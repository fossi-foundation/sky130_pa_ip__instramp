magic
tech sky130A
timestamp 1730992408
<< pwell >>
rect -164 -379 164 379
<< mvnmos >>
rect -50 -250 50 250
<< mvndiff >>
rect -79 244 -50 250
rect -79 -244 -73 244
rect -56 -244 -50 244
rect -79 -250 -50 -244
rect 50 244 79 250
rect 50 -244 56 244
rect 73 -244 79 244
rect 50 -250 79 -244
<< mvndiffc >>
rect -73 -244 -56 244
rect 56 -244 73 244
<< mvpsubdiff >>
rect -146 355 146 361
rect -146 338 -92 355
rect 92 338 146 355
rect -146 332 146 338
rect -146 307 -117 332
rect -146 -307 -140 307
rect -123 -307 -117 307
rect 117 307 146 332
rect -146 -332 -117 -307
rect 117 -307 123 307
rect 140 -307 146 307
rect 117 -332 146 -307
rect -146 -338 146 -332
rect -146 -355 -92 -338
rect 92 -355 146 -338
rect -146 -361 146 -355
<< mvpsubdiffcont >>
rect -92 338 92 355
rect -140 -307 -123 307
rect 123 -307 140 307
rect -92 -355 92 -338
<< poly >>
rect -50 286 50 294
rect -50 269 -42 286
rect 42 269 50 286
rect -50 250 50 269
rect -50 -269 50 -250
rect -50 -286 -42 -269
rect 42 -286 50 -269
rect -50 -294 50 -286
<< polycont >>
rect -42 269 42 286
rect -42 -286 42 -269
<< locali >>
rect -140 338 -92 355
rect 92 338 140 355
rect -140 307 -123 338
rect 123 307 140 338
rect -50 269 -42 286
rect 42 269 50 286
rect -73 244 -56 252
rect -73 -252 -56 -244
rect 56 244 73 252
rect 56 -252 73 -244
rect -50 -286 -42 -269
rect 42 -286 50 -269
rect -140 -338 -123 -307
rect 123 -338 140 -307
rect -140 -355 -92 -338
rect 92 -355 140 -338
<< viali >>
rect -42 269 42 286
rect -73 -244 -56 244
rect 56 -244 73 244
rect -42 -286 42 -269
<< metal1 >>
rect -48 286 48 289
rect -48 269 -42 286
rect 42 269 48 286
rect -48 266 48 269
rect -76 244 -53 250
rect -76 -244 -73 244
rect -56 -244 -53 244
rect -76 -250 -53 -244
rect 53 244 76 250
rect 53 -244 56 244
rect 73 -244 76 244
rect 53 -250 76 -244
rect -48 -269 48 -266
rect -48 -286 -42 -269
rect 42 -286 48 -269
rect -48 -289 48 -286
<< properties >>
string FIXED_BBOX -131 -346 131 346
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 ad {int((nf+1)/2) * W/nf * 0.29} as {int((nf+2)/2) * W/nf * 0.29} pd {2*int((nf+1)/2) * (W/nf + 0.29)} ps {2*int((nf+2)/2) * (W/nf + 0.29)} nrd {0.29 / W} nrs {0.29 / W} sa 0 sb 0 sd 0 mult 1
<< end >>
