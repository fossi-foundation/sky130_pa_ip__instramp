magic
tech sky130A
magscale 1 2
timestamp 1748312405
<< dnwell >>
rect 84 80 29486 37640
<< nwell >>
rect 4 37432 29566 37720
rect 4 33252 290 37432
rect 29280 33252 29566 37432
rect 4 24578 348 33252
rect 29218 24578 29566 33252
rect 4 23504 290 24578
rect 29280 23532 29566 24578
rect 4 14830 356 23504
rect 29220 14858 29566 23532
rect 4 13784 290 14830
rect 29278 14434 29566 14858
rect 29280 13784 29566 14434
rect 4 5110 356 13784
rect 29222 5110 29566 13784
rect 4 308 290 5110
rect 29278 4686 29566 5110
rect 29280 308 29566 4686
rect 4 0 29566 308
<< nsubdiff >>
rect 136 37580 29446 37592
rect 136 37526 268 37580
rect 29322 37526 29446 37580
rect 136 37514 29446 37526
rect 136 37472 214 37514
rect 136 262 146 37472
rect 202 262 214 37472
rect 136 181 214 262
rect 29367 37488 29446 37514
rect 29367 278 29378 37488
rect 29434 278 29446 37488
rect 29367 181 29446 278
rect 136 170 29446 181
rect 136 116 290 170
rect 29344 116 29446 170
rect 136 102 29446 116
<< nsubdiffcont >>
rect 268 37526 29322 37580
rect 146 262 202 37472
rect 29378 278 29434 37488
rect 290 116 29344 170
<< locali >>
rect 136 37562 268 37580
rect 136 120 144 37562
rect 204 37526 268 37562
rect 29322 37560 29446 37580
rect 29322 37526 29374 37560
rect 204 37468 346 37526
rect 2816 37468 29374 37526
rect 204 37442 29374 37468
rect 204 181 214 37442
rect 14464 26920 16102 27532
rect 13472 17176 16096 17816
rect 13466 7458 16104 8062
rect 29367 181 29374 37442
rect 204 174 29374 181
rect 204 120 290 174
rect 29316 170 29374 174
rect 136 110 290 120
rect 29344 116 29374 170
rect 29316 114 29374 116
rect 29436 114 29446 37560
rect 29316 110 29446 114
rect 136 102 29446 110
<< viali >>
rect 144 37472 204 37562
rect 346 37526 2816 37536
rect 144 262 146 37472
rect 146 262 202 37472
rect 202 262 204 37472
rect 346 37468 2816 37526
rect 29374 37488 29436 37560
rect 144 120 204 262
rect 29374 278 29378 37488
rect 29378 278 29434 37488
rect 29434 278 29436 37488
rect 290 170 29316 174
rect 290 116 29316 170
rect 290 110 29316 116
rect 29374 114 29436 278
<< metal1 >>
rect 1636 39187 1836 39814
rect 2824 39614 3049 39814
rect 436 39112 936 39134
rect 1636 39130 3211 39187
rect 5271 39130 5563 39187
rect 436 38846 454 39112
rect 916 39102 936 39112
rect 916 38852 2908 39102
rect 916 38846 936 38852
rect 436 38828 936 38846
rect 1986 37854 2668 37870
rect 1986 37652 2022 37854
rect 2654 37782 2668 37854
rect 2654 37652 5122 37782
rect 1986 37638 5122 37652
rect 136 37572 214 37580
rect 136 37562 2872 37572
rect 136 25116 144 37562
rect 204 37536 2872 37562
rect 204 37468 346 37536
rect 2816 37468 2872 37536
rect 204 37442 2872 37468
rect 29366 37560 29446 37580
rect 136 24158 142 25116
rect 136 15364 144 24158
rect 204 19616 214 37442
rect 1278 33645 1344 34079
rect 1278 33579 2876 33645
rect 2810 32735 2876 33579
rect 29366 29368 29374 37560
rect 29436 29368 29446 37560
rect 29366 28528 29372 29368
rect 29438 28528 29446 29368
rect 206 18782 214 19616
rect 204 15364 214 18782
rect 2812 15594 3166 15608
rect 2812 15502 2830 15594
rect 3148 15502 3166 15594
rect 2812 15490 3166 15502
rect 136 14414 142 15364
rect 206 14414 214 15364
rect 136 120 144 14414
rect 204 5644 214 14414
rect 29366 15390 29374 28528
rect 29436 19646 29446 28528
rect 29440 18812 29446 19646
rect 29436 15390 29446 18812
rect 29366 14446 29372 15390
rect 29438 14446 29446 15390
rect 26370 14280 26762 14290
rect 26370 14188 26390 14280
rect 26748 14188 26762 14280
rect 26370 14174 26762 14188
rect 13460 7456 14596 8028
rect 14954 7456 16106 8066
rect 206 4696 214 5644
rect 204 182 214 4696
rect 14281 4594 14754 4672
rect 13904 4578 14360 4594
rect 13904 4484 13918 4578
rect 14342 4484 14360 4578
rect 13904 4472 14360 4484
rect 29366 182 29374 14446
rect 29436 9896 29446 14446
rect 29438 9064 29446 9896
rect 204 174 29374 182
rect 204 120 290 174
rect 136 110 290 120
rect 29316 114 29374 174
rect 29436 114 29446 9064
rect 29316 110 29446 114
rect 136 102 29446 110
<< via1 >>
rect 454 38846 916 39112
rect 2022 37652 2654 37854
rect 146 28530 204 29362
rect 142 24158 144 25116
rect 144 24158 204 25116
rect 1144 35326 1344 35462
rect 29372 28528 29374 29368
rect 29374 28528 29436 29368
rect 29436 28528 29438 29368
rect 15256 23346 19932 23398
rect 146 18782 204 19616
rect 204 18782 206 19616
rect 2830 15502 3148 15594
rect 142 14414 144 15364
rect 144 14414 204 15364
rect 204 14414 206 15364
rect 146 9058 204 9898
rect 29380 24168 29436 25108
rect 29374 18812 29436 19646
rect 29436 18812 29440 19646
rect 29372 14446 29374 15390
rect 29374 14446 29436 15390
rect 29436 14446 29438 15390
rect 26390 14188 26748 14280
rect 144 4696 204 5644
rect 204 4696 206 5644
rect 144 2482 202 3624
rect 13918 4484 14342 4578
rect 29374 9064 29436 9896
rect 29436 9064 29438 9896
rect 29380 4696 29432 5640
rect 29376 2482 29434 3622
<< metal2 >>
rect 4718 39842 4918 40042
rect 7118 39842 7318 40042
rect 9518 39842 9718 40042
rect 11918 39842 12118 40042
rect 14318 39842 14518 40042
rect 16718 39842 16918 40042
rect 19118 39842 19318 40042
rect 21518 39842 21718 40042
rect 23918 39842 24118 40042
rect 26318 39842 26518 40042
rect 436 39112 936 39134
rect 436 38846 454 39112
rect 916 38846 936 39112
rect 436 38828 936 38846
rect 1986 37854 2668 37870
rect 1986 37652 2022 37854
rect 2654 37652 2668 37854
rect 1986 37638 2668 37652
rect 0 35462 200 35490
rect 0 35326 1144 35462
rect 1344 35326 1362 35462
rect 0 35290 200 35326
rect 2278 34482 2682 34498
rect 2278 33710 2408 34482
rect 2656 33710 2682 34482
rect 2278 33696 2682 33710
rect 132 29362 444 29376
rect 132 28530 146 29362
rect 204 28530 444 29362
rect 132 28520 444 28530
rect 29122 29368 29448 29376
rect 29122 28528 29372 29368
rect 29438 28528 29448 29368
rect 29122 28520 29448 28528
rect 134 25116 442 25122
rect 134 24158 142 25116
rect 204 24158 442 25116
rect 134 24152 442 24158
rect 29118 25108 29446 25122
rect 29118 24168 29380 25108
rect 29436 24168 29446 25108
rect 29118 24152 29446 24168
rect 2 23842 316 24042
rect 29122 19646 29450 19656
rect 122 19616 450 19628
rect 122 18782 146 19616
rect 206 18782 450 19616
rect 29122 18812 29374 19646
rect 29440 18812 29450 19646
rect 29122 18800 29450 18812
rect 122 18772 450 18782
rect 2812 15594 3166 15608
rect 2812 15502 2830 15594
rect 3148 15502 3166 15594
rect 2812 15490 3166 15502
rect 29116 15390 29458 15402
rect 126 15364 450 15374
rect 126 14414 142 15364
rect 206 14414 450 15364
rect 29116 14446 29372 15390
rect 29438 14446 29458 15390
rect 29116 14432 29458 14446
rect 126 14404 450 14414
rect 4 14118 312 14318
rect 26370 14280 26762 14290
rect 26370 14188 26390 14280
rect 26748 14188 26762 14280
rect 26370 14174 26762 14188
rect 128 9898 450 9908
rect 128 9058 146 9898
rect 204 9058 450 9898
rect 128 9052 450 9058
rect 29122 9896 29450 9908
rect 29122 9064 29374 9896
rect 29438 9064 29450 9896
rect 29122 9052 29450 9064
rect 130 5644 450 5654
rect 130 4696 144 5644
rect 206 4696 450 5644
rect 130 4684 450 4696
rect 29128 5640 29452 5654
rect 29128 4696 29380 5640
rect 29432 4696 29452 5640
rect 29128 4684 29452 4696
rect 2 4424 402 4624
rect 7386 4578 14356 4592
rect 7386 4484 13918 4578
rect 14342 4484 14356 4578
rect 7386 4464 14356 4484
rect 20 3624 29530 3636
rect 20 2482 144 3624
rect 202 3622 29530 3624
rect 202 3598 29376 3622
rect 202 2496 476 3598
rect 906 3596 29376 3598
rect 906 2496 28678 3596
rect 202 2494 28678 2496
rect 29108 2494 29376 3596
rect 202 2482 29376 2494
rect 29434 2482 29530 3622
rect 20 2472 29530 2482
rect 22 2210 29532 2238
rect 22 2204 26926 2210
rect 22 1096 2428 2204
rect 2646 1102 26926 2204
rect 27144 1102 29532 2210
rect 2646 1096 29532 1102
rect 22 1074 29532 1096
<< via2 >>
rect 454 38846 916 39112
rect 2022 37652 2654 37854
rect 2408 33710 2656 34482
rect 2830 15502 3148 15594
rect 26390 14188 26748 14280
rect 476 2496 906 3598
rect 28678 2494 29108 3596
rect 2428 1096 2646 2204
rect 26926 1102 27144 2210
<< metal3 >>
rect 436 39112 936 39822
rect 436 38846 454 39112
rect 916 38846 936 39112
rect 436 33508 936 38846
rect 2010 38012 2668 39822
rect 2010 37854 27166 38012
rect 2010 37652 2022 37854
rect 2654 37652 27166 37854
rect 2010 37643 27166 37652
rect 2010 34482 2668 37643
rect 2010 33710 2408 34482
rect 2656 33710 2668 34482
rect 2010 33522 2668 33710
rect 2010 33174 2400 33522
rect 2812 15594 3166 15608
rect 2812 15502 2830 15594
rect 3148 15502 3166 15594
rect 2812 15490 3166 15502
rect 2822 14280 2922 15490
rect 26370 14280 26762 14290
rect 2816 14188 26390 14280
rect 26748 14188 26762 14280
rect 2816 14180 26762 14188
rect 26370 14174 26762 14180
rect 444 3598 944 4694
rect 444 2496 476 3598
rect 906 2496 944 3598
rect 444 304 944 2496
rect 2406 2204 2676 5914
rect 2406 1096 2428 2204
rect 2646 1096 2676 2204
rect 2406 320 2676 1096
rect 14840 0 15052 200
use Parallel_10B_Block2  x1
timestamp 1748312405
transform -1 0 29706 0 1 11584
box 364 -11384 29514 28258
use Input_Stage_v1  x2
timestamp 1748312405
transform -1 0 29402 0 1 41468
box 14048 -37044 29188 -7862
use vbias_gen_pga  x3
timestamp 1730992408
transform 1 0 1455 0 1 34561
box -311 -865 845 909
<< labels >>
flabel metal2 0 35290 200 35490 0 FreeSans 256 0 0 0 IBIAS
port 11 nsew
flabel metal2 2 23842 202 24042 0 FreeSans 256 0 0 0 VCM
port 10 nsew
flabel metal3 14848 0 15048 200 0 FreeSans 256 0 0 0 VOUT
port 15 nsew
flabel metal3 564 39612 764 39812 0 FreeSans 256 0 0 0 AVDD
port 12 nsew
flabel metal3 2256 39614 2456 39814 0 FreeSans 256 0 0 0 AVSS
port 16 nsew
flabel metal2 26318 39842 26518 40042 0 FreeSans 256 90 0 0 V[0]
port 9 nsew
flabel metal2 23918 39842 24118 40042 0 FreeSans 256 90 0 0 V[1]
port 8 nsew
flabel metal2 21518 39842 21718 40042 0 FreeSans 256 90 0 0 V[2]
port 7 nsew
flabel metal2 19118 39842 19318 40042 0 FreeSans 256 90 0 0 V[3]
port 6 nsew
flabel metal2 16718 39842 16918 40042 0 FreeSans 256 90 0 0 V[4]
port 5 nsew
flabel metal2 14318 39842 14518 40042 0 FreeSans 256 90 0 0 V[5]
port 4 nsew
flabel metal2 11918 39842 12118 40042 0 FreeSans 256 90 0 0 V[6]
port 3 nsew
flabel metal2 9518 39842 9718 40042 0 FreeSans 256 90 0 0 V[7]
port 2 nsew
flabel metal2 7118 39842 7318 40042 0 FreeSans 256 90 0 0 V[8]
port 1 nsew
flabel metal2 4718 39842 4918 40042 0 FreeSans 256 90 0 0 V[9]
port 0 nsew
flabel metal1 2824 39614 3024 39814 0 FreeSans 256 0 0 0 DVSS
port 17 nsew
flabel metal1 1636 39614 1836 39814 0 FreeSans 256 0 0 0 DVDD
port 14 nsew
flabel metal2 4 14118 204 14318 0 FreeSans 256 0 0 0 VINP
port 13 nsew
flabel metal2 2 4424 202 4624 0 FreeSans 480 0 0 0 VINN
port 18 nsew
<< properties >>
string MASKHINTS_HVI 2806 39814 26901 39875
<< end >>
