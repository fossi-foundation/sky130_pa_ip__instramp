magic
tech sky130A
magscale 1 2
timestamp 1730739923
<< metal3 >>
rect -3798 5652 -1426 5680
rect -3798 3628 -1510 5652
rect -1446 3628 -1426 5652
rect -3798 3600 -1426 3628
rect -1186 5652 1186 5680
rect -1186 3628 1102 5652
rect 1166 3628 1186 5652
rect -1186 3600 1186 3628
rect 1426 5652 3798 5680
rect 1426 3628 3714 5652
rect 3778 3628 3798 5652
rect 1426 3600 3798 3628
rect -3798 3332 -1426 3360
rect -3798 1308 -1510 3332
rect -1446 1308 -1426 3332
rect -3798 1280 -1426 1308
rect -1186 3332 1186 3360
rect -1186 1308 1102 3332
rect 1166 1308 1186 3332
rect -1186 1280 1186 1308
rect 1426 3332 3798 3360
rect 1426 1308 3714 3332
rect 3778 1308 3798 3332
rect 1426 1280 3798 1308
rect -3798 1012 -1426 1040
rect -3798 -1012 -1510 1012
rect -1446 -1012 -1426 1012
rect -3798 -1040 -1426 -1012
rect -1186 1012 1186 1040
rect -1186 -1012 1102 1012
rect 1166 -1012 1186 1012
rect -1186 -1040 1186 -1012
rect 1426 1012 3798 1040
rect 1426 -1012 3714 1012
rect 3778 -1012 3798 1012
rect 1426 -1040 3798 -1012
rect -3798 -1308 -1426 -1280
rect -3798 -3332 -1510 -1308
rect -1446 -3332 -1426 -1308
rect -3798 -3360 -1426 -3332
rect -1186 -1308 1186 -1280
rect -1186 -3332 1102 -1308
rect 1166 -3332 1186 -1308
rect -1186 -3360 1186 -3332
rect 1426 -1308 3798 -1280
rect 1426 -3332 3714 -1308
rect 3778 -3332 3798 -1308
rect 1426 -3360 3798 -3332
rect -3798 -3628 -1426 -3600
rect -3798 -5652 -1510 -3628
rect -1446 -5652 -1426 -3628
rect -3798 -5680 -1426 -5652
rect -1186 -3628 1186 -3600
rect -1186 -5652 1102 -3628
rect 1166 -5652 1186 -3628
rect -1186 -5680 1186 -5652
rect 1426 -3628 3798 -3600
rect 1426 -5652 3714 -3628
rect 3778 -5652 3798 -3628
rect 1426 -5680 3798 -5652
<< via3 >>
rect -1510 3628 -1446 5652
rect 1102 3628 1166 5652
rect 3714 3628 3778 5652
rect -1510 1308 -1446 3332
rect 1102 1308 1166 3332
rect 3714 1308 3778 3332
rect -1510 -1012 -1446 1012
rect 1102 -1012 1166 1012
rect 3714 -1012 3778 1012
rect -1510 -3332 -1446 -1308
rect 1102 -3332 1166 -1308
rect 3714 -3332 3778 -1308
rect -1510 -5652 -1446 -3628
rect 1102 -5652 1166 -3628
rect 3714 -5652 3778 -3628
<< mimcap >>
rect -3758 5600 -1758 5640
rect -3758 3680 -3718 5600
rect -1798 3680 -1758 5600
rect -3758 3640 -1758 3680
rect -1146 5600 854 5640
rect -1146 3680 -1106 5600
rect 814 3680 854 5600
rect -1146 3640 854 3680
rect 1466 5600 3466 5640
rect 1466 3680 1506 5600
rect 3426 3680 3466 5600
rect 1466 3640 3466 3680
rect -3758 3280 -1758 3320
rect -3758 1360 -3718 3280
rect -1798 1360 -1758 3280
rect -3758 1320 -1758 1360
rect -1146 3280 854 3320
rect -1146 1360 -1106 3280
rect 814 1360 854 3280
rect -1146 1320 854 1360
rect 1466 3280 3466 3320
rect 1466 1360 1506 3280
rect 3426 1360 3466 3280
rect 1466 1320 3466 1360
rect -3758 960 -1758 1000
rect -3758 -960 -3718 960
rect -1798 -960 -1758 960
rect -3758 -1000 -1758 -960
rect -1146 960 854 1000
rect -1146 -960 -1106 960
rect 814 -960 854 960
rect -1146 -1000 854 -960
rect 1466 960 3466 1000
rect 1466 -960 1506 960
rect 3426 -960 3466 960
rect 1466 -1000 3466 -960
rect -3758 -1360 -1758 -1320
rect -3758 -3280 -3718 -1360
rect -1798 -3280 -1758 -1360
rect -3758 -3320 -1758 -3280
rect -1146 -1360 854 -1320
rect -1146 -3280 -1106 -1360
rect 814 -3280 854 -1360
rect -1146 -3320 854 -3280
rect 1466 -1360 3466 -1320
rect 1466 -3280 1506 -1360
rect 3426 -3280 3466 -1360
rect 1466 -3320 3466 -3280
rect -3758 -3680 -1758 -3640
rect -3758 -5600 -3718 -3680
rect -1798 -5600 -1758 -3680
rect -3758 -5640 -1758 -5600
rect -1146 -3680 854 -3640
rect -1146 -5600 -1106 -3680
rect 814 -5600 854 -3680
rect -1146 -5640 854 -5600
rect 1466 -3680 3466 -3640
rect 1466 -5600 1506 -3680
rect 3426 -5600 3466 -3680
rect 1466 -5640 3466 -5600
<< mimcapcontact >>
rect -3718 3680 -1798 5600
rect -1106 3680 814 5600
rect 1506 3680 3426 5600
rect -3718 1360 -1798 3280
rect -1106 1360 814 3280
rect 1506 1360 3426 3280
rect -3718 -960 -1798 960
rect -1106 -960 814 960
rect 1506 -960 3426 960
rect -3718 -3280 -1798 -1360
rect -1106 -3280 814 -1360
rect 1506 -3280 3426 -1360
rect -3718 -5600 -1798 -3680
rect -1106 -5600 814 -3680
rect 1506 -5600 3426 -3680
<< metal4 >>
rect -2810 5601 -2706 5800
rect -1530 5652 -1426 5800
rect -3719 5600 -1797 5601
rect -3719 3680 -3718 5600
rect -1798 3680 -1797 5600
rect -3719 3679 -1797 3680
rect -2810 3281 -2706 3679
rect -1530 3628 -1510 5652
rect -1446 3628 -1426 5652
rect -198 5601 -94 5800
rect 1082 5652 1186 5800
rect -1107 5600 815 5601
rect -1107 3680 -1106 5600
rect 814 3680 815 5600
rect -1107 3679 815 3680
rect -1530 3332 -1426 3628
rect -3719 3280 -1797 3281
rect -3719 1360 -3718 3280
rect -1798 1360 -1797 3280
rect -3719 1359 -1797 1360
rect -2810 961 -2706 1359
rect -1530 1308 -1510 3332
rect -1446 1308 -1426 3332
rect -198 3281 -94 3679
rect 1082 3628 1102 5652
rect 1166 3628 1186 5652
rect 2414 5601 2518 5800
rect 3694 5652 3798 5800
rect 1505 5600 3427 5601
rect 1505 3680 1506 5600
rect 3426 3680 3427 5600
rect 1505 3679 3427 3680
rect 1082 3332 1186 3628
rect -1107 3280 815 3281
rect -1107 1360 -1106 3280
rect 814 1360 815 3280
rect -1107 1359 815 1360
rect -1530 1012 -1426 1308
rect -3719 960 -1797 961
rect -3719 -960 -3718 960
rect -1798 -960 -1797 960
rect -3719 -961 -1797 -960
rect -2810 -1359 -2706 -961
rect -1530 -1012 -1510 1012
rect -1446 -1012 -1426 1012
rect -198 961 -94 1359
rect 1082 1308 1102 3332
rect 1166 1308 1186 3332
rect 2414 3281 2518 3679
rect 3694 3628 3714 5652
rect 3778 3628 3798 5652
rect 3694 3332 3798 3628
rect 1505 3280 3427 3281
rect 1505 1360 1506 3280
rect 3426 1360 3427 3280
rect 1505 1359 3427 1360
rect 1082 1012 1186 1308
rect -1107 960 815 961
rect -1107 -960 -1106 960
rect 814 -960 815 960
rect -1107 -961 815 -960
rect -1530 -1308 -1426 -1012
rect -3719 -1360 -1797 -1359
rect -3719 -3280 -3718 -1360
rect -1798 -3280 -1797 -1360
rect -3719 -3281 -1797 -3280
rect -2810 -3679 -2706 -3281
rect -1530 -3332 -1510 -1308
rect -1446 -3332 -1426 -1308
rect -198 -1359 -94 -961
rect 1082 -1012 1102 1012
rect 1166 -1012 1186 1012
rect 2414 961 2518 1359
rect 3694 1308 3714 3332
rect 3778 1308 3798 3332
rect 3694 1012 3798 1308
rect 1505 960 3427 961
rect 1505 -960 1506 960
rect 3426 -960 3427 960
rect 1505 -961 3427 -960
rect 1082 -1308 1186 -1012
rect -1107 -1360 815 -1359
rect -1107 -3280 -1106 -1360
rect 814 -3280 815 -1360
rect -1107 -3281 815 -3280
rect -1530 -3628 -1426 -3332
rect -3719 -3680 -1797 -3679
rect -3719 -5600 -3718 -3680
rect -1798 -5600 -1797 -3680
rect -3719 -5601 -1797 -5600
rect -2810 -5800 -2706 -5601
rect -1530 -5652 -1510 -3628
rect -1446 -5652 -1426 -3628
rect -198 -3679 -94 -3281
rect 1082 -3332 1102 -1308
rect 1166 -3332 1186 -1308
rect 2414 -1359 2518 -961
rect 3694 -1012 3714 1012
rect 3778 -1012 3798 1012
rect 3694 -1308 3798 -1012
rect 1505 -1360 3427 -1359
rect 1505 -3280 1506 -1360
rect 3426 -3280 3427 -1360
rect 1505 -3281 3427 -3280
rect 1082 -3628 1186 -3332
rect -1107 -3680 815 -3679
rect -1107 -5600 -1106 -3680
rect 814 -5600 815 -3680
rect -1107 -5601 815 -5600
rect -1530 -5800 -1426 -5652
rect -198 -5800 -94 -5601
rect 1082 -5652 1102 -3628
rect 1166 -5652 1186 -3628
rect 2414 -3679 2518 -3281
rect 3694 -3332 3714 -1308
rect 3778 -3332 3798 -1308
rect 3694 -3628 3798 -3332
rect 1505 -3680 3427 -3679
rect 1505 -5600 1506 -3680
rect 3426 -5600 3427 -3680
rect 1505 -5601 3427 -5600
rect 1082 -5800 1186 -5652
rect 2414 -5800 2518 -5601
rect 3694 -5652 3714 -3628
rect 3778 -5652 3798 -3628
rect 3694 -5800 3798 -5652
<< properties >>
string FIXED_BBOX 1426 3600 3506 5680
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10.0 l 10.0 val 207.6 carea 2.00 cperi 0.19 class capacitor nx 3 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
