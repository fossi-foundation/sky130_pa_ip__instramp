magic
tech sky130A
magscale 1 2
timestamp 1729620069
<< pwell >>
rect -30070 -8050 30070 8050
<< psubdiff >>
rect -30034 7980 -29938 8014
rect 29938 7980 30034 8014
rect -30034 7918 -30000 7980
rect 30000 7918 30034 7980
rect -30034 -7980 -30000 -7918
rect 30000 -7980 30034 -7918
rect -30034 -8014 -29938 -7980
rect 29938 -8014 30034 -7980
<< psubdiffcont >>
rect -29938 7980 29938 8014
rect -30034 -7918 -30000 7918
rect 30000 -7918 30034 7918
rect -29938 -8014 29938 -7980
<< xpolycontact >>
rect -29904 7452 -29766 7884
rect -29904 52 -29766 484
rect -29670 7452 -29532 7884
rect -29670 52 -29532 484
rect -29436 7452 -29298 7884
rect -29436 52 -29298 484
rect -29202 7452 -29064 7884
rect -29202 52 -29064 484
rect -28968 7452 -28830 7884
rect -28968 52 -28830 484
rect -28734 7452 -28596 7884
rect -28734 52 -28596 484
rect -28500 7452 -28362 7884
rect -28500 52 -28362 484
rect -28266 7452 -28128 7884
rect -28266 52 -28128 484
rect -28032 7452 -27894 7884
rect -28032 52 -27894 484
rect -27798 7452 -27660 7884
rect -27798 52 -27660 484
rect -27564 7452 -27426 7884
rect -27564 52 -27426 484
rect -27330 7452 -27192 7884
rect -27330 52 -27192 484
rect -27096 7452 -26958 7884
rect -27096 52 -26958 484
rect -26862 7452 -26724 7884
rect -26862 52 -26724 484
rect -26628 7452 -26490 7884
rect -26628 52 -26490 484
rect -26394 7452 -26256 7884
rect -26394 52 -26256 484
rect -26160 7452 -26022 7884
rect -26160 52 -26022 484
rect -25926 7452 -25788 7884
rect -25926 52 -25788 484
rect -25692 7452 -25554 7884
rect -25692 52 -25554 484
rect -25458 7452 -25320 7884
rect -25458 52 -25320 484
rect -25224 7452 -25086 7884
rect -25224 52 -25086 484
rect -24990 7452 -24852 7884
rect -24990 52 -24852 484
rect -24756 7452 -24618 7884
rect -24756 52 -24618 484
rect -24522 7452 -24384 7884
rect -24522 52 -24384 484
rect -24288 7452 -24150 7884
rect -24288 52 -24150 484
rect -24054 7452 -23916 7884
rect -24054 52 -23916 484
rect -23820 7452 -23682 7884
rect -23820 52 -23682 484
rect -23586 7452 -23448 7884
rect -23586 52 -23448 484
rect -23352 7452 -23214 7884
rect -23352 52 -23214 484
rect -23118 7452 -22980 7884
rect -23118 52 -22980 484
rect -22884 7452 -22746 7884
rect -22884 52 -22746 484
rect -22650 7452 -22512 7884
rect -22650 52 -22512 484
rect -22416 7452 -22278 7884
rect -22416 52 -22278 484
rect -22182 7452 -22044 7884
rect -22182 52 -22044 484
rect -21948 7452 -21810 7884
rect -21948 52 -21810 484
rect -21714 7452 -21576 7884
rect -21714 52 -21576 484
rect -21480 7452 -21342 7884
rect -21480 52 -21342 484
rect -21246 7452 -21108 7884
rect -21246 52 -21108 484
rect -21012 7452 -20874 7884
rect -21012 52 -20874 484
rect -20778 7452 -20640 7884
rect -20778 52 -20640 484
rect -20544 7452 -20406 7884
rect -20544 52 -20406 484
rect -20310 7452 -20172 7884
rect -20310 52 -20172 484
rect -20076 7452 -19938 7884
rect -20076 52 -19938 484
rect -19842 7452 -19704 7884
rect -19842 52 -19704 484
rect -19608 7452 -19470 7884
rect -19608 52 -19470 484
rect -19374 7452 -19236 7884
rect -19374 52 -19236 484
rect -19140 7452 -19002 7884
rect -19140 52 -19002 484
rect -18906 7452 -18768 7884
rect -18906 52 -18768 484
rect -18672 7452 -18534 7884
rect -18672 52 -18534 484
rect -18438 7452 -18300 7884
rect -18438 52 -18300 484
rect -18204 7452 -18066 7884
rect -18204 52 -18066 484
rect -17970 7452 -17832 7884
rect -17970 52 -17832 484
rect -17736 7452 -17598 7884
rect -17736 52 -17598 484
rect -17502 7452 -17364 7884
rect -17502 52 -17364 484
rect -17268 7452 -17130 7884
rect -17268 52 -17130 484
rect -17034 7452 -16896 7884
rect -17034 52 -16896 484
rect -16800 7452 -16662 7884
rect -16800 52 -16662 484
rect -16566 7452 -16428 7884
rect -16566 52 -16428 484
rect -16332 7452 -16194 7884
rect -16332 52 -16194 484
rect -16098 7452 -15960 7884
rect -16098 52 -15960 484
rect -15864 7452 -15726 7884
rect -15864 52 -15726 484
rect -15630 7452 -15492 7884
rect -15630 52 -15492 484
rect -15396 7452 -15258 7884
rect -15396 52 -15258 484
rect -15162 7452 -15024 7884
rect -15162 52 -15024 484
rect -14928 7452 -14790 7884
rect -14928 52 -14790 484
rect -14694 7452 -14556 7884
rect -14694 52 -14556 484
rect -14460 7452 -14322 7884
rect -14460 52 -14322 484
rect -14226 7452 -14088 7884
rect -14226 52 -14088 484
rect -13992 7452 -13854 7884
rect -13992 52 -13854 484
rect -13758 7452 -13620 7884
rect -13758 52 -13620 484
rect -13524 7452 -13386 7884
rect -13524 52 -13386 484
rect -13290 7452 -13152 7884
rect -13290 52 -13152 484
rect -13056 7452 -12918 7884
rect -13056 52 -12918 484
rect -12822 7452 -12684 7884
rect -12822 52 -12684 484
rect -12588 7452 -12450 7884
rect -12588 52 -12450 484
rect -12354 7452 -12216 7884
rect -12354 52 -12216 484
rect -12120 7452 -11982 7884
rect -12120 52 -11982 484
rect -11886 7452 -11748 7884
rect -11886 52 -11748 484
rect -11652 7452 -11514 7884
rect -11652 52 -11514 484
rect -11418 7452 -11280 7884
rect -11418 52 -11280 484
rect -11184 7452 -11046 7884
rect -11184 52 -11046 484
rect -10950 7452 -10812 7884
rect -10950 52 -10812 484
rect -10716 7452 -10578 7884
rect -10716 52 -10578 484
rect -10482 7452 -10344 7884
rect -10482 52 -10344 484
rect -10248 7452 -10110 7884
rect -10248 52 -10110 484
rect -10014 7452 -9876 7884
rect -10014 52 -9876 484
rect -9780 7452 -9642 7884
rect -9780 52 -9642 484
rect -9546 7452 -9408 7884
rect -9546 52 -9408 484
rect -9312 7452 -9174 7884
rect -9312 52 -9174 484
rect -9078 7452 -8940 7884
rect -9078 52 -8940 484
rect -8844 7452 -8706 7884
rect -8844 52 -8706 484
rect -8610 7452 -8472 7884
rect -8610 52 -8472 484
rect -8376 7452 -8238 7884
rect -8376 52 -8238 484
rect -8142 7452 -8004 7884
rect -8142 52 -8004 484
rect -7908 7452 -7770 7884
rect -7908 52 -7770 484
rect -7674 7452 -7536 7884
rect -7674 52 -7536 484
rect -7440 7452 -7302 7884
rect -7440 52 -7302 484
rect -7206 7452 -7068 7884
rect -7206 52 -7068 484
rect -6972 7452 -6834 7884
rect -6972 52 -6834 484
rect -6738 7452 -6600 7884
rect -6738 52 -6600 484
rect -6504 7452 -6366 7884
rect -6504 52 -6366 484
rect -6270 7452 -6132 7884
rect -6270 52 -6132 484
rect -6036 7452 -5898 7884
rect -6036 52 -5898 484
rect -5802 7452 -5664 7884
rect -5802 52 -5664 484
rect -5568 7452 -5430 7884
rect -5568 52 -5430 484
rect -5334 7452 -5196 7884
rect -5334 52 -5196 484
rect -5100 7452 -4962 7884
rect -5100 52 -4962 484
rect -4866 7452 -4728 7884
rect -4866 52 -4728 484
rect -4632 7452 -4494 7884
rect -4632 52 -4494 484
rect -4398 7452 -4260 7884
rect -4398 52 -4260 484
rect -4164 7452 -4026 7884
rect -4164 52 -4026 484
rect -3930 7452 -3792 7884
rect -3930 52 -3792 484
rect -3696 7452 -3558 7884
rect -3696 52 -3558 484
rect -3462 7452 -3324 7884
rect -3462 52 -3324 484
rect -3228 7452 -3090 7884
rect -3228 52 -3090 484
rect -2994 7452 -2856 7884
rect -2994 52 -2856 484
rect -2760 7452 -2622 7884
rect -2760 52 -2622 484
rect -2526 7452 -2388 7884
rect -2526 52 -2388 484
rect -2292 7452 -2154 7884
rect -2292 52 -2154 484
rect -2058 7452 -1920 7884
rect -2058 52 -1920 484
rect -1824 7452 -1686 7884
rect -1824 52 -1686 484
rect -1590 7452 -1452 7884
rect -1590 52 -1452 484
rect -1356 7452 -1218 7884
rect -1356 52 -1218 484
rect -1122 7452 -984 7884
rect -1122 52 -984 484
rect -888 7452 -750 7884
rect -888 52 -750 484
rect -654 7452 -516 7884
rect -654 52 -516 484
rect -420 7452 -282 7884
rect -420 52 -282 484
rect -186 7452 -48 7884
rect -186 52 -48 484
rect 48 7452 186 7884
rect 48 52 186 484
rect 282 7452 420 7884
rect 282 52 420 484
rect 516 7452 654 7884
rect 516 52 654 484
rect 750 7452 888 7884
rect 750 52 888 484
rect 984 7452 1122 7884
rect 984 52 1122 484
rect 1218 7452 1356 7884
rect 1218 52 1356 484
rect 1452 7452 1590 7884
rect 1452 52 1590 484
rect 1686 7452 1824 7884
rect 1686 52 1824 484
rect 1920 7452 2058 7884
rect 1920 52 2058 484
rect 2154 7452 2292 7884
rect 2154 52 2292 484
rect 2388 7452 2526 7884
rect 2388 52 2526 484
rect 2622 7452 2760 7884
rect 2622 52 2760 484
rect 2856 7452 2994 7884
rect 2856 52 2994 484
rect 3090 7452 3228 7884
rect 3090 52 3228 484
rect 3324 7452 3462 7884
rect 3324 52 3462 484
rect 3558 7452 3696 7884
rect 3558 52 3696 484
rect 3792 7452 3930 7884
rect 3792 52 3930 484
rect 4026 7452 4164 7884
rect 4026 52 4164 484
rect 4260 7452 4398 7884
rect 4260 52 4398 484
rect 4494 7452 4632 7884
rect 4494 52 4632 484
rect 4728 7452 4866 7884
rect 4728 52 4866 484
rect 4962 7452 5100 7884
rect 4962 52 5100 484
rect 5196 7452 5334 7884
rect 5196 52 5334 484
rect 5430 7452 5568 7884
rect 5430 52 5568 484
rect 5664 7452 5802 7884
rect 5664 52 5802 484
rect 5898 7452 6036 7884
rect 5898 52 6036 484
rect 6132 7452 6270 7884
rect 6132 52 6270 484
rect 6366 7452 6504 7884
rect 6366 52 6504 484
rect 6600 7452 6738 7884
rect 6600 52 6738 484
rect 6834 7452 6972 7884
rect 6834 52 6972 484
rect 7068 7452 7206 7884
rect 7068 52 7206 484
rect 7302 7452 7440 7884
rect 7302 52 7440 484
rect 7536 7452 7674 7884
rect 7536 52 7674 484
rect 7770 7452 7908 7884
rect 7770 52 7908 484
rect 8004 7452 8142 7884
rect 8004 52 8142 484
rect 8238 7452 8376 7884
rect 8238 52 8376 484
rect 8472 7452 8610 7884
rect 8472 52 8610 484
rect 8706 7452 8844 7884
rect 8706 52 8844 484
rect 8940 7452 9078 7884
rect 8940 52 9078 484
rect 9174 7452 9312 7884
rect 9174 52 9312 484
rect 9408 7452 9546 7884
rect 9408 52 9546 484
rect 9642 7452 9780 7884
rect 9642 52 9780 484
rect 9876 7452 10014 7884
rect 9876 52 10014 484
rect 10110 7452 10248 7884
rect 10110 52 10248 484
rect 10344 7452 10482 7884
rect 10344 52 10482 484
rect 10578 7452 10716 7884
rect 10578 52 10716 484
rect 10812 7452 10950 7884
rect 10812 52 10950 484
rect 11046 7452 11184 7884
rect 11046 52 11184 484
rect 11280 7452 11418 7884
rect 11280 52 11418 484
rect 11514 7452 11652 7884
rect 11514 52 11652 484
rect 11748 7452 11886 7884
rect 11748 52 11886 484
rect 11982 7452 12120 7884
rect 11982 52 12120 484
rect 12216 7452 12354 7884
rect 12216 52 12354 484
rect 12450 7452 12588 7884
rect 12450 52 12588 484
rect 12684 7452 12822 7884
rect 12684 52 12822 484
rect 12918 7452 13056 7884
rect 12918 52 13056 484
rect 13152 7452 13290 7884
rect 13152 52 13290 484
rect 13386 7452 13524 7884
rect 13386 52 13524 484
rect 13620 7452 13758 7884
rect 13620 52 13758 484
rect 13854 7452 13992 7884
rect 13854 52 13992 484
rect 14088 7452 14226 7884
rect 14088 52 14226 484
rect 14322 7452 14460 7884
rect 14322 52 14460 484
rect 14556 7452 14694 7884
rect 14556 52 14694 484
rect 14790 7452 14928 7884
rect 14790 52 14928 484
rect 15024 7452 15162 7884
rect 15024 52 15162 484
rect 15258 7452 15396 7884
rect 15258 52 15396 484
rect 15492 7452 15630 7884
rect 15492 52 15630 484
rect 15726 7452 15864 7884
rect 15726 52 15864 484
rect 15960 7452 16098 7884
rect 15960 52 16098 484
rect 16194 7452 16332 7884
rect 16194 52 16332 484
rect 16428 7452 16566 7884
rect 16428 52 16566 484
rect 16662 7452 16800 7884
rect 16662 52 16800 484
rect 16896 7452 17034 7884
rect 16896 52 17034 484
rect 17130 7452 17268 7884
rect 17130 52 17268 484
rect 17364 7452 17502 7884
rect 17364 52 17502 484
rect 17598 7452 17736 7884
rect 17598 52 17736 484
rect 17832 7452 17970 7884
rect 17832 52 17970 484
rect 18066 7452 18204 7884
rect 18066 52 18204 484
rect 18300 7452 18438 7884
rect 18300 52 18438 484
rect 18534 7452 18672 7884
rect 18534 52 18672 484
rect 18768 7452 18906 7884
rect 18768 52 18906 484
rect 19002 7452 19140 7884
rect 19002 52 19140 484
rect 19236 7452 19374 7884
rect 19236 52 19374 484
rect 19470 7452 19608 7884
rect 19470 52 19608 484
rect 19704 7452 19842 7884
rect 19704 52 19842 484
rect 19938 7452 20076 7884
rect 19938 52 20076 484
rect 20172 7452 20310 7884
rect 20172 52 20310 484
rect 20406 7452 20544 7884
rect 20406 52 20544 484
rect 20640 7452 20778 7884
rect 20640 52 20778 484
rect 20874 7452 21012 7884
rect 20874 52 21012 484
rect 21108 7452 21246 7884
rect 21108 52 21246 484
rect 21342 7452 21480 7884
rect 21342 52 21480 484
rect 21576 7452 21714 7884
rect 21576 52 21714 484
rect 21810 7452 21948 7884
rect 21810 52 21948 484
rect 22044 7452 22182 7884
rect 22044 52 22182 484
rect 22278 7452 22416 7884
rect 22278 52 22416 484
rect 22512 7452 22650 7884
rect 22512 52 22650 484
rect 22746 7452 22884 7884
rect 22746 52 22884 484
rect 22980 7452 23118 7884
rect 22980 52 23118 484
rect 23214 7452 23352 7884
rect 23214 52 23352 484
rect 23448 7452 23586 7884
rect 23448 52 23586 484
rect 23682 7452 23820 7884
rect 23682 52 23820 484
rect 23916 7452 24054 7884
rect 23916 52 24054 484
rect 24150 7452 24288 7884
rect 24150 52 24288 484
rect 24384 7452 24522 7884
rect 24384 52 24522 484
rect 24618 7452 24756 7884
rect 24618 52 24756 484
rect 24852 7452 24990 7884
rect 24852 52 24990 484
rect 25086 7452 25224 7884
rect 25086 52 25224 484
rect 25320 7452 25458 7884
rect 25320 52 25458 484
rect 25554 7452 25692 7884
rect 25554 52 25692 484
rect 25788 7452 25926 7884
rect 25788 52 25926 484
rect 26022 7452 26160 7884
rect 26022 52 26160 484
rect 26256 7452 26394 7884
rect 26256 52 26394 484
rect 26490 7452 26628 7884
rect 26490 52 26628 484
rect 26724 7452 26862 7884
rect 26724 52 26862 484
rect 26958 7452 27096 7884
rect 26958 52 27096 484
rect 27192 7452 27330 7884
rect 27192 52 27330 484
rect 27426 7452 27564 7884
rect 27426 52 27564 484
rect 27660 7452 27798 7884
rect 27660 52 27798 484
rect 27894 7452 28032 7884
rect 27894 52 28032 484
rect 28128 7452 28266 7884
rect 28128 52 28266 484
rect 28362 7452 28500 7884
rect 28362 52 28500 484
rect 28596 7452 28734 7884
rect 28596 52 28734 484
rect 28830 7452 28968 7884
rect 28830 52 28968 484
rect 29064 7452 29202 7884
rect 29064 52 29202 484
rect 29298 7452 29436 7884
rect 29298 52 29436 484
rect 29532 7452 29670 7884
rect 29532 52 29670 484
rect 29766 7452 29904 7884
rect 29766 52 29904 484
rect -29904 -484 -29766 -52
rect -29904 -7884 -29766 -7452
rect -29670 -484 -29532 -52
rect -29670 -7884 -29532 -7452
rect -29436 -484 -29298 -52
rect -29436 -7884 -29298 -7452
rect -29202 -484 -29064 -52
rect -29202 -7884 -29064 -7452
rect -28968 -484 -28830 -52
rect -28968 -7884 -28830 -7452
rect -28734 -484 -28596 -52
rect -28734 -7884 -28596 -7452
rect -28500 -484 -28362 -52
rect -28500 -7884 -28362 -7452
rect -28266 -484 -28128 -52
rect -28266 -7884 -28128 -7452
rect -28032 -484 -27894 -52
rect -28032 -7884 -27894 -7452
rect -27798 -484 -27660 -52
rect -27798 -7884 -27660 -7452
rect -27564 -484 -27426 -52
rect -27564 -7884 -27426 -7452
rect -27330 -484 -27192 -52
rect -27330 -7884 -27192 -7452
rect -27096 -484 -26958 -52
rect -27096 -7884 -26958 -7452
rect -26862 -484 -26724 -52
rect -26862 -7884 -26724 -7452
rect -26628 -484 -26490 -52
rect -26628 -7884 -26490 -7452
rect -26394 -484 -26256 -52
rect -26394 -7884 -26256 -7452
rect -26160 -484 -26022 -52
rect -26160 -7884 -26022 -7452
rect -25926 -484 -25788 -52
rect -25926 -7884 -25788 -7452
rect -25692 -484 -25554 -52
rect -25692 -7884 -25554 -7452
rect -25458 -484 -25320 -52
rect -25458 -7884 -25320 -7452
rect -25224 -484 -25086 -52
rect -25224 -7884 -25086 -7452
rect -24990 -484 -24852 -52
rect -24990 -7884 -24852 -7452
rect -24756 -484 -24618 -52
rect -24756 -7884 -24618 -7452
rect -24522 -484 -24384 -52
rect -24522 -7884 -24384 -7452
rect -24288 -484 -24150 -52
rect -24288 -7884 -24150 -7452
rect -24054 -484 -23916 -52
rect -24054 -7884 -23916 -7452
rect -23820 -484 -23682 -52
rect -23820 -7884 -23682 -7452
rect -23586 -484 -23448 -52
rect -23586 -7884 -23448 -7452
rect -23352 -484 -23214 -52
rect -23352 -7884 -23214 -7452
rect -23118 -484 -22980 -52
rect -23118 -7884 -22980 -7452
rect -22884 -484 -22746 -52
rect -22884 -7884 -22746 -7452
rect -22650 -484 -22512 -52
rect -22650 -7884 -22512 -7452
rect -22416 -484 -22278 -52
rect -22416 -7884 -22278 -7452
rect -22182 -484 -22044 -52
rect -22182 -7884 -22044 -7452
rect -21948 -484 -21810 -52
rect -21948 -7884 -21810 -7452
rect -21714 -484 -21576 -52
rect -21714 -7884 -21576 -7452
rect -21480 -484 -21342 -52
rect -21480 -7884 -21342 -7452
rect -21246 -484 -21108 -52
rect -21246 -7884 -21108 -7452
rect -21012 -484 -20874 -52
rect -21012 -7884 -20874 -7452
rect -20778 -484 -20640 -52
rect -20778 -7884 -20640 -7452
rect -20544 -484 -20406 -52
rect -20544 -7884 -20406 -7452
rect -20310 -484 -20172 -52
rect -20310 -7884 -20172 -7452
rect -20076 -484 -19938 -52
rect -20076 -7884 -19938 -7452
rect -19842 -484 -19704 -52
rect -19842 -7884 -19704 -7452
rect -19608 -484 -19470 -52
rect -19608 -7884 -19470 -7452
rect -19374 -484 -19236 -52
rect -19374 -7884 -19236 -7452
rect -19140 -484 -19002 -52
rect -19140 -7884 -19002 -7452
rect -18906 -484 -18768 -52
rect -18906 -7884 -18768 -7452
rect -18672 -484 -18534 -52
rect -18672 -7884 -18534 -7452
rect -18438 -484 -18300 -52
rect -18438 -7884 -18300 -7452
rect -18204 -484 -18066 -52
rect -18204 -7884 -18066 -7452
rect -17970 -484 -17832 -52
rect -17970 -7884 -17832 -7452
rect -17736 -484 -17598 -52
rect -17736 -7884 -17598 -7452
rect -17502 -484 -17364 -52
rect -17502 -7884 -17364 -7452
rect -17268 -484 -17130 -52
rect -17268 -7884 -17130 -7452
rect -17034 -484 -16896 -52
rect -17034 -7884 -16896 -7452
rect -16800 -484 -16662 -52
rect -16800 -7884 -16662 -7452
rect -16566 -484 -16428 -52
rect -16566 -7884 -16428 -7452
rect -16332 -484 -16194 -52
rect -16332 -7884 -16194 -7452
rect -16098 -484 -15960 -52
rect -16098 -7884 -15960 -7452
rect -15864 -484 -15726 -52
rect -15864 -7884 -15726 -7452
rect -15630 -484 -15492 -52
rect -15630 -7884 -15492 -7452
rect -15396 -484 -15258 -52
rect -15396 -7884 -15258 -7452
rect -15162 -484 -15024 -52
rect -15162 -7884 -15024 -7452
rect -14928 -484 -14790 -52
rect -14928 -7884 -14790 -7452
rect -14694 -484 -14556 -52
rect -14694 -7884 -14556 -7452
rect -14460 -484 -14322 -52
rect -14460 -7884 -14322 -7452
rect -14226 -484 -14088 -52
rect -14226 -7884 -14088 -7452
rect -13992 -484 -13854 -52
rect -13992 -7884 -13854 -7452
rect -13758 -484 -13620 -52
rect -13758 -7884 -13620 -7452
rect -13524 -484 -13386 -52
rect -13524 -7884 -13386 -7452
rect -13290 -484 -13152 -52
rect -13290 -7884 -13152 -7452
rect -13056 -484 -12918 -52
rect -13056 -7884 -12918 -7452
rect -12822 -484 -12684 -52
rect -12822 -7884 -12684 -7452
rect -12588 -484 -12450 -52
rect -12588 -7884 -12450 -7452
rect -12354 -484 -12216 -52
rect -12354 -7884 -12216 -7452
rect -12120 -484 -11982 -52
rect -12120 -7884 -11982 -7452
rect -11886 -484 -11748 -52
rect -11886 -7884 -11748 -7452
rect -11652 -484 -11514 -52
rect -11652 -7884 -11514 -7452
rect -11418 -484 -11280 -52
rect -11418 -7884 -11280 -7452
rect -11184 -484 -11046 -52
rect -11184 -7884 -11046 -7452
rect -10950 -484 -10812 -52
rect -10950 -7884 -10812 -7452
rect -10716 -484 -10578 -52
rect -10716 -7884 -10578 -7452
rect -10482 -484 -10344 -52
rect -10482 -7884 -10344 -7452
rect -10248 -484 -10110 -52
rect -10248 -7884 -10110 -7452
rect -10014 -484 -9876 -52
rect -10014 -7884 -9876 -7452
rect -9780 -484 -9642 -52
rect -9780 -7884 -9642 -7452
rect -9546 -484 -9408 -52
rect -9546 -7884 -9408 -7452
rect -9312 -484 -9174 -52
rect -9312 -7884 -9174 -7452
rect -9078 -484 -8940 -52
rect -9078 -7884 -8940 -7452
rect -8844 -484 -8706 -52
rect -8844 -7884 -8706 -7452
rect -8610 -484 -8472 -52
rect -8610 -7884 -8472 -7452
rect -8376 -484 -8238 -52
rect -8376 -7884 -8238 -7452
rect -8142 -484 -8004 -52
rect -8142 -7884 -8004 -7452
rect -7908 -484 -7770 -52
rect -7908 -7884 -7770 -7452
rect -7674 -484 -7536 -52
rect -7674 -7884 -7536 -7452
rect -7440 -484 -7302 -52
rect -7440 -7884 -7302 -7452
rect -7206 -484 -7068 -52
rect -7206 -7884 -7068 -7452
rect -6972 -484 -6834 -52
rect -6972 -7884 -6834 -7452
rect -6738 -484 -6600 -52
rect -6738 -7884 -6600 -7452
rect -6504 -484 -6366 -52
rect -6504 -7884 -6366 -7452
rect -6270 -484 -6132 -52
rect -6270 -7884 -6132 -7452
rect -6036 -484 -5898 -52
rect -6036 -7884 -5898 -7452
rect -5802 -484 -5664 -52
rect -5802 -7884 -5664 -7452
rect -5568 -484 -5430 -52
rect -5568 -7884 -5430 -7452
rect -5334 -484 -5196 -52
rect -5334 -7884 -5196 -7452
rect -5100 -484 -4962 -52
rect -5100 -7884 -4962 -7452
rect -4866 -484 -4728 -52
rect -4866 -7884 -4728 -7452
rect -4632 -484 -4494 -52
rect -4632 -7884 -4494 -7452
rect -4398 -484 -4260 -52
rect -4398 -7884 -4260 -7452
rect -4164 -484 -4026 -52
rect -4164 -7884 -4026 -7452
rect -3930 -484 -3792 -52
rect -3930 -7884 -3792 -7452
rect -3696 -484 -3558 -52
rect -3696 -7884 -3558 -7452
rect -3462 -484 -3324 -52
rect -3462 -7884 -3324 -7452
rect -3228 -484 -3090 -52
rect -3228 -7884 -3090 -7452
rect -2994 -484 -2856 -52
rect -2994 -7884 -2856 -7452
rect -2760 -484 -2622 -52
rect -2760 -7884 -2622 -7452
rect -2526 -484 -2388 -52
rect -2526 -7884 -2388 -7452
rect -2292 -484 -2154 -52
rect -2292 -7884 -2154 -7452
rect -2058 -484 -1920 -52
rect -2058 -7884 -1920 -7452
rect -1824 -484 -1686 -52
rect -1824 -7884 -1686 -7452
rect -1590 -484 -1452 -52
rect -1590 -7884 -1452 -7452
rect -1356 -484 -1218 -52
rect -1356 -7884 -1218 -7452
rect -1122 -484 -984 -52
rect -1122 -7884 -984 -7452
rect -888 -484 -750 -52
rect -888 -7884 -750 -7452
rect -654 -484 -516 -52
rect -654 -7884 -516 -7452
rect -420 -484 -282 -52
rect -420 -7884 -282 -7452
rect -186 -484 -48 -52
rect -186 -7884 -48 -7452
rect 48 -484 186 -52
rect 48 -7884 186 -7452
rect 282 -484 420 -52
rect 282 -7884 420 -7452
rect 516 -484 654 -52
rect 516 -7884 654 -7452
rect 750 -484 888 -52
rect 750 -7884 888 -7452
rect 984 -484 1122 -52
rect 984 -7884 1122 -7452
rect 1218 -484 1356 -52
rect 1218 -7884 1356 -7452
rect 1452 -484 1590 -52
rect 1452 -7884 1590 -7452
rect 1686 -484 1824 -52
rect 1686 -7884 1824 -7452
rect 1920 -484 2058 -52
rect 1920 -7884 2058 -7452
rect 2154 -484 2292 -52
rect 2154 -7884 2292 -7452
rect 2388 -484 2526 -52
rect 2388 -7884 2526 -7452
rect 2622 -484 2760 -52
rect 2622 -7884 2760 -7452
rect 2856 -484 2994 -52
rect 2856 -7884 2994 -7452
rect 3090 -484 3228 -52
rect 3090 -7884 3228 -7452
rect 3324 -484 3462 -52
rect 3324 -7884 3462 -7452
rect 3558 -484 3696 -52
rect 3558 -7884 3696 -7452
rect 3792 -484 3930 -52
rect 3792 -7884 3930 -7452
rect 4026 -484 4164 -52
rect 4026 -7884 4164 -7452
rect 4260 -484 4398 -52
rect 4260 -7884 4398 -7452
rect 4494 -484 4632 -52
rect 4494 -7884 4632 -7452
rect 4728 -484 4866 -52
rect 4728 -7884 4866 -7452
rect 4962 -484 5100 -52
rect 4962 -7884 5100 -7452
rect 5196 -484 5334 -52
rect 5196 -7884 5334 -7452
rect 5430 -484 5568 -52
rect 5430 -7884 5568 -7452
rect 5664 -484 5802 -52
rect 5664 -7884 5802 -7452
rect 5898 -484 6036 -52
rect 5898 -7884 6036 -7452
rect 6132 -484 6270 -52
rect 6132 -7884 6270 -7452
rect 6366 -484 6504 -52
rect 6366 -7884 6504 -7452
rect 6600 -484 6738 -52
rect 6600 -7884 6738 -7452
rect 6834 -484 6972 -52
rect 6834 -7884 6972 -7452
rect 7068 -484 7206 -52
rect 7068 -7884 7206 -7452
rect 7302 -484 7440 -52
rect 7302 -7884 7440 -7452
rect 7536 -484 7674 -52
rect 7536 -7884 7674 -7452
rect 7770 -484 7908 -52
rect 7770 -7884 7908 -7452
rect 8004 -484 8142 -52
rect 8004 -7884 8142 -7452
rect 8238 -484 8376 -52
rect 8238 -7884 8376 -7452
rect 8472 -484 8610 -52
rect 8472 -7884 8610 -7452
rect 8706 -484 8844 -52
rect 8706 -7884 8844 -7452
rect 8940 -484 9078 -52
rect 8940 -7884 9078 -7452
rect 9174 -484 9312 -52
rect 9174 -7884 9312 -7452
rect 9408 -484 9546 -52
rect 9408 -7884 9546 -7452
rect 9642 -484 9780 -52
rect 9642 -7884 9780 -7452
rect 9876 -484 10014 -52
rect 9876 -7884 10014 -7452
rect 10110 -484 10248 -52
rect 10110 -7884 10248 -7452
rect 10344 -484 10482 -52
rect 10344 -7884 10482 -7452
rect 10578 -484 10716 -52
rect 10578 -7884 10716 -7452
rect 10812 -484 10950 -52
rect 10812 -7884 10950 -7452
rect 11046 -484 11184 -52
rect 11046 -7884 11184 -7452
rect 11280 -484 11418 -52
rect 11280 -7884 11418 -7452
rect 11514 -484 11652 -52
rect 11514 -7884 11652 -7452
rect 11748 -484 11886 -52
rect 11748 -7884 11886 -7452
rect 11982 -484 12120 -52
rect 11982 -7884 12120 -7452
rect 12216 -484 12354 -52
rect 12216 -7884 12354 -7452
rect 12450 -484 12588 -52
rect 12450 -7884 12588 -7452
rect 12684 -484 12822 -52
rect 12684 -7884 12822 -7452
rect 12918 -484 13056 -52
rect 12918 -7884 13056 -7452
rect 13152 -484 13290 -52
rect 13152 -7884 13290 -7452
rect 13386 -484 13524 -52
rect 13386 -7884 13524 -7452
rect 13620 -484 13758 -52
rect 13620 -7884 13758 -7452
rect 13854 -484 13992 -52
rect 13854 -7884 13992 -7452
rect 14088 -484 14226 -52
rect 14088 -7884 14226 -7452
rect 14322 -484 14460 -52
rect 14322 -7884 14460 -7452
rect 14556 -484 14694 -52
rect 14556 -7884 14694 -7452
rect 14790 -484 14928 -52
rect 14790 -7884 14928 -7452
rect 15024 -484 15162 -52
rect 15024 -7884 15162 -7452
rect 15258 -484 15396 -52
rect 15258 -7884 15396 -7452
rect 15492 -484 15630 -52
rect 15492 -7884 15630 -7452
rect 15726 -484 15864 -52
rect 15726 -7884 15864 -7452
rect 15960 -484 16098 -52
rect 15960 -7884 16098 -7452
rect 16194 -484 16332 -52
rect 16194 -7884 16332 -7452
rect 16428 -484 16566 -52
rect 16428 -7884 16566 -7452
rect 16662 -484 16800 -52
rect 16662 -7884 16800 -7452
rect 16896 -484 17034 -52
rect 16896 -7884 17034 -7452
rect 17130 -484 17268 -52
rect 17130 -7884 17268 -7452
rect 17364 -484 17502 -52
rect 17364 -7884 17502 -7452
rect 17598 -484 17736 -52
rect 17598 -7884 17736 -7452
rect 17832 -484 17970 -52
rect 17832 -7884 17970 -7452
rect 18066 -484 18204 -52
rect 18066 -7884 18204 -7452
rect 18300 -484 18438 -52
rect 18300 -7884 18438 -7452
rect 18534 -484 18672 -52
rect 18534 -7884 18672 -7452
rect 18768 -484 18906 -52
rect 18768 -7884 18906 -7452
rect 19002 -484 19140 -52
rect 19002 -7884 19140 -7452
rect 19236 -484 19374 -52
rect 19236 -7884 19374 -7452
rect 19470 -484 19608 -52
rect 19470 -7884 19608 -7452
rect 19704 -484 19842 -52
rect 19704 -7884 19842 -7452
rect 19938 -484 20076 -52
rect 19938 -7884 20076 -7452
rect 20172 -484 20310 -52
rect 20172 -7884 20310 -7452
rect 20406 -484 20544 -52
rect 20406 -7884 20544 -7452
rect 20640 -484 20778 -52
rect 20640 -7884 20778 -7452
rect 20874 -484 21012 -52
rect 20874 -7884 21012 -7452
rect 21108 -484 21246 -52
rect 21108 -7884 21246 -7452
rect 21342 -484 21480 -52
rect 21342 -7884 21480 -7452
rect 21576 -484 21714 -52
rect 21576 -7884 21714 -7452
rect 21810 -484 21948 -52
rect 21810 -7884 21948 -7452
rect 22044 -484 22182 -52
rect 22044 -7884 22182 -7452
rect 22278 -484 22416 -52
rect 22278 -7884 22416 -7452
rect 22512 -484 22650 -52
rect 22512 -7884 22650 -7452
rect 22746 -484 22884 -52
rect 22746 -7884 22884 -7452
rect 22980 -484 23118 -52
rect 22980 -7884 23118 -7452
rect 23214 -484 23352 -52
rect 23214 -7884 23352 -7452
rect 23448 -484 23586 -52
rect 23448 -7884 23586 -7452
rect 23682 -484 23820 -52
rect 23682 -7884 23820 -7452
rect 23916 -484 24054 -52
rect 23916 -7884 24054 -7452
rect 24150 -484 24288 -52
rect 24150 -7884 24288 -7452
rect 24384 -484 24522 -52
rect 24384 -7884 24522 -7452
rect 24618 -484 24756 -52
rect 24618 -7884 24756 -7452
rect 24852 -484 24990 -52
rect 24852 -7884 24990 -7452
rect 25086 -484 25224 -52
rect 25086 -7884 25224 -7452
rect 25320 -484 25458 -52
rect 25320 -7884 25458 -7452
rect 25554 -484 25692 -52
rect 25554 -7884 25692 -7452
rect 25788 -484 25926 -52
rect 25788 -7884 25926 -7452
rect 26022 -484 26160 -52
rect 26022 -7884 26160 -7452
rect 26256 -484 26394 -52
rect 26256 -7884 26394 -7452
rect 26490 -484 26628 -52
rect 26490 -7884 26628 -7452
rect 26724 -484 26862 -52
rect 26724 -7884 26862 -7452
rect 26958 -484 27096 -52
rect 26958 -7884 27096 -7452
rect 27192 -484 27330 -52
rect 27192 -7884 27330 -7452
rect 27426 -484 27564 -52
rect 27426 -7884 27564 -7452
rect 27660 -484 27798 -52
rect 27660 -7884 27798 -7452
rect 27894 -484 28032 -52
rect 27894 -7884 28032 -7452
rect 28128 -484 28266 -52
rect 28128 -7884 28266 -7452
rect 28362 -484 28500 -52
rect 28362 -7884 28500 -7452
rect 28596 -484 28734 -52
rect 28596 -7884 28734 -7452
rect 28830 -484 28968 -52
rect 28830 -7884 28968 -7452
rect 29064 -484 29202 -52
rect 29064 -7884 29202 -7452
rect 29298 -484 29436 -52
rect 29298 -7884 29436 -7452
rect 29532 -484 29670 -52
rect 29532 -7884 29670 -7452
rect 29766 -484 29904 -52
rect 29766 -7884 29904 -7452
<< ppolyres >>
rect -29904 484 -29766 7452
rect -29670 484 -29532 7452
rect -29436 484 -29298 7452
rect -29202 484 -29064 7452
rect -28968 484 -28830 7452
rect -28734 484 -28596 7452
rect -28500 484 -28362 7452
rect -28266 484 -28128 7452
rect -28032 484 -27894 7452
rect -27798 484 -27660 7452
rect -27564 484 -27426 7452
rect -27330 484 -27192 7452
rect -27096 484 -26958 7452
rect -26862 484 -26724 7452
rect -26628 484 -26490 7452
rect -26394 484 -26256 7452
rect -26160 484 -26022 7452
rect -25926 484 -25788 7452
rect -25692 484 -25554 7452
rect -25458 484 -25320 7452
rect -25224 484 -25086 7452
rect -24990 484 -24852 7452
rect -24756 484 -24618 7452
rect -24522 484 -24384 7452
rect -24288 484 -24150 7452
rect -24054 484 -23916 7452
rect -23820 484 -23682 7452
rect -23586 484 -23448 7452
rect -23352 484 -23214 7452
rect -23118 484 -22980 7452
rect -22884 484 -22746 7452
rect -22650 484 -22512 7452
rect -22416 484 -22278 7452
rect -22182 484 -22044 7452
rect -21948 484 -21810 7452
rect -21714 484 -21576 7452
rect -21480 484 -21342 7452
rect -21246 484 -21108 7452
rect -21012 484 -20874 7452
rect -20778 484 -20640 7452
rect -20544 484 -20406 7452
rect -20310 484 -20172 7452
rect -20076 484 -19938 7452
rect -19842 484 -19704 7452
rect -19608 484 -19470 7452
rect -19374 484 -19236 7452
rect -19140 484 -19002 7452
rect -18906 484 -18768 7452
rect -18672 484 -18534 7452
rect -18438 484 -18300 7452
rect -18204 484 -18066 7452
rect -17970 484 -17832 7452
rect -17736 484 -17598 7452
rect -17502 484 -17364 7452
rect -17268 484 -17130 7452
rect -17034 484 -16896 7452
rect -16800 484 -16662 7452
rect -16566 484 -16428 7452
rect -16332 484 -16194 7452
rect -16098 484 -15960 7452
rect -15864 484 -15726 7452
rect -15630 484 -15492 7452
rect -15396 484 -15258 7452
rect -15162 484 -15024 7452
rect -14928 484 -14790 7452
rect -14694 484 -14556 7452
rect -14460 484 -14322 7452
rect -14226 484 -14088 7452
rect -13992 484 -13854 7452
rect -13758 484 -13620 7452
rect -13524 484 -13386 7452
rect -13290 484 -13152 7452
rect -13056 484 -12918 7452
rect -12822 484 -12684 7452
rect -12588 484 -12450 7452
rect -12354 484 -12216 7452
rect -12120 484 -11982 7452
rect -11886 484 -11748 7452
rect -11652 484 -11514 7452
rect -11418 484 -11280 7452
rect -11184 484 -11046 7452
rect -10950 484 -10812 7452
rect -10716 484 -10578 7452
rect -10482 484 -10344 7452
rect -10248 484 -10110 7452
rect -10014 484 -9876 7452
rect -9780 484 -9642 7452
rect -9546 484 -9408 7452
rect -9312 484 -9174 7452
rect -9078 484 -8940 7452
rect -8844 484 -8706 7452
rect -8610 484 -8472 7452
rect -8376 484 -8238 7452
rect -8142 484 -8004 7452
rect -7908 484 -7770 7452
rect -7674 484 -7536 7452
rect -7440 484 -7302 7452
rect -7206 484 -7068 7452
rect -6972 484 -6834 7452
rect -6738 484 -6600 7452
rect -6504 484 -6366 7452
rect -6270 484 -6132 7452
rect -6036 484 -5898 7452
rect -5802 484 -5664 7452
rect -5568 484 -5430 7452
rect -5334 484 -5196 7452
rect -5100 484 -4962 7452
rect -4866 484 -4728 7452
rect -4632 484 -4494 7452
rect -4398 484 -4260 7452
rect -4164 484 -4026 7452
rect -3930 484 -3792 7452
rect -3696 484 -3558 7452
rect -3462 484 -3324 7452
rect -3228 484 -3090 7452
rect -2994 484 -2856 7452
rect -2760 484 -2622 7452
rect -2526 484 -2388 7452
rect -2292 484 -2154 7452
rect -2058 484 -1920 7452
rect -1824 484 -1686 7452
rect -1590 484 -1452 7452
rect -1356 484 -1218 7452
rect -1122 484 -984 7452
rect -888 484 -750 7452
rect -654 484 -516 7452
rect -420 484 -282 7452
rect -186 484 -48 7452
rect 48 484 186 7452
rect 282 484 420 7452
rect 516 484 654 7452
rect 750 484 888 7452
rect 984 484 1122 7452
rect 1218 484 1356 7452
rect 1452 484 1590 7452
rect 1686 484 1824 7452
rect 1920 484 2058 7452
rect 2154 484 2292 7452
rect 2388 484 2526 7452
rect 2622 484 2760 7452
rect 2856 484 2994 7452
rect 3090 484 3228 7452
rect 3324 484 3462 7452
rect 3558 484 3696 7452
rect 3792 484 3930 7452
rect 4026 484 4164 7452
rect 4260 484 4398 7452
rect 4494 484 4632 7452
rect 4728 484 4866 7452
rect 4962 484 5100 7452
rect 5196 484 5334 7452
rect 5430 484 5568 7452
rect 5664 484 5802 7452
rect 5898 484 6036 7452
rect 6132 484 6270 7452
rect 6366 484 6504 7452
rect 6600 484 6738 7452
rect 6834 484 6972 7452
rect 7068 484 7206 7452
rect 7302 484 7440 7452
rect 7536 484 7674 7452
rect 7770 484 7908 7452
rect 8004 484 8142 7452
rect 8238 484 8376 7452
rect 8472 484 8610 7452
rect 8706 484 8844 7452
rect 8940 484 9078 7452
rect 9174 484 9312 7452
rect 9408 484 9546 7452
rect 9642 484 9780 7452
rect 9876 484 10014 7452
rect 10110 484 10248 7452
rect 10344 484 10482 7452
rect 10578 484 10716 7452
rect 10812 484 10950 7452
rect 11046 484 11184 7452
rect 11280 484 11418 7452
rect 11514 484 11652 7452
rect 11748 484 11886 7452
rect 11982 484 12120 7452
rect 12216 484 12354 7452
rect 12450 484 12588 7452
rect 12684 484 12822 7452
rect 12918 484 13056 7452
rect 13152 484 13290 7452
rect 13386 484 13524 7452
rect 13620 484 13758 7452
rect 13854 484 13992 7452
rect 14088 484 14226 7452
rect 14322 484 14460 7452
rect 14556 484 14694 7452
rect 14790 484 14928 7452
rect 15024 484 15162 7452
rect 15258 484 15396 7452
rect 15492 484 15630 7452
rect 15726 484 15864 7452
rect 15960 484 16098 7452
rect 16194 484 16332 7452
rect 16428 484 16566 7452
rect 16662 484 16800 7452
rect 16896 484 17034 7452
rect 17130 484 17268 7452
rect 17364 484 17502 7452
rect 17598 484 17736 7452
rect 17832 484 17970 7452
rect 18066 484 18204 7452
rect 18300 484 18438 7452
rect 18534 484 18672 7452
rect 18768 484 18906 7452
rect 19002 484 19140 7452
rect 19236 484 19374 7452
rect 19470 484 19608 7452
rect 19704 484 19842 7452
rect 19938 484 20076 7452
rect 20172 484 20310 7452
rect 20406 484 20544 7452
rect 20640 484 20778 7452
rect 20874 484 21012 7452
rect 21108 484 21246 7452
rect 21342 484 21480 7452
rect 21576 484 21714 7452
rect 21810 484 21948 7452
rect 22044 484 22182 7452
rect 22278 484 22416 7452
rect 22512 484 22650 7452
rect 22746 484 22884 7452
rect 22980 484 23118 7452
rect 23214 484 23352 7452
rect 23448 484 23586 7452
rect 23682 484 23820 7452
rect 23916 484 24054 7452
rect 24150 484 24288 7452
rect 24384 484 24522 7452
rect 24618 484 24756 7452
rect 24852 484 24990 7452
rect 25086 484 25224 7452
rect 25320 484 25458 7452
rect 25554 484 25692 7452
rect 25788 484 25926 7452
rect 26022 484 26160 7452
rect 26256 484 26394 7452
rect 26490 484 26628 7452
rect 26724 484 26862 7452
rect 26958 484 27096 7452
rect 27192 484 27330 7452
rect 27426 484 27564 7452
rect 27660 484 27798 7452
rect 27894 484 28032 7452
rect 28128 484 28266 7452
rect 28362 484 28500 7452
rect 28596 484 28734 7452
rect 28830 484 28968 7452
rect 29064 484 29202 7452
rect 29298 484 29436 7452
rect 29532 484 29670 7452
rect 29766 484 29904 7452
rect -29904 -7452 -29766 -484
rect -29670 -7452 -29532 -484
rect -29436 -7452 -29298 -484
rect -29202 -7452 -29064 -484
rect -28968 -7452 -28830 -484
rect -28734 -7452 -28596 -484
rect -28500 -7452 -28362 -484
rect -28266 -7452 -28128 -484
rect -28032 -7452 -27894 -484
rect -27798 -7452 -27660 -484
rect -27564 -7452 -27426 -484
rect -27330 -7452 -27192 -484
rect -27096 -7452 -26958 -484
rect -26862 -7452 -26724 -484
rect -26628 -7452 -26490 -484
rect -26394 -7452 -26256 -484
rect -26160 -7452 -26022 -484
rect -25926 -7452 -25788 -484
rect -25692 -7452 -25554 -484
rect -25458 -7452 -25320 -484
rect -25224 -7452 -25086 -484
rect -24990 -7452 -24852 -484
rect -24756 -7452 -24618 -484
rect -24522 -7452 -24384 -484
rect -24288 -7452 -24150 -484
rect -24054 -7452 -23916 -484
rect -23820 -7452 -23682 -484
rect -23586 -7452 -23448 -484
rect -23352 -7452 -23214 -484
rect -23118 -7452 -22980 -484
rect -22884 -7452 -22746 -484
rect -22650 -7452 -22512 -484
rect -22416 -7452 -22278 -484
rect -22182 -7452 -22044 -484
rect -21948 -7452 -21810 -484
rect -21714 -7452 -21576 -484
rect -21480 -7452 -21342 -484
rect -21246 -7452 -21108 -484
rect -21012 -7452 -20874 -484
rect -20778 -7452 -20640 -484
rect -20544 -7452 -20406 -484
rect -20310 -7452 -20172 -484
rect -20076 -7452 -19938 -484
rect -19842 -7452 -19704 -484
rect -19608 -7452 -19470 -484
rect -19374 -7452 -19236 -484
rect -19140 -7452 -19002 -484
rect -18906 -7452 -18768 -484
rect -18672 -7452 -18534 -484
rect -18438 -7452 -18300 -484
rect -18204 -7452 -18066 -484
rect -17970 -7452 -17832 -484
rect -17736 -7452 -17598 -484
rect -17502 -7452 -17364 -484
rect -17268 -7452 -17130 -484
rect -17034 -7452 -16896 -484
rect -16800 -7452 -16662 -484
rect -16566 -7452 -16428 -484
rect -16332 -7452 -16194 -484
rect -16098 -7452 -15960 -484
rect -15864 -7452 -15726 -484
rect -15630 -7452 -15492 -484
rect -15396 -7452 -15258 -484
rect -15162 -7452 -15024 -484
rect -14928 -7452 -14790 -484
rect -14694 -7452 -14556 -484
rect -14460 -7452 -14322 -484
rect -14226 -7452 -14088 -484
rect -13992 -7452 -13854 -484
rect -13758 -7452 -13620 -484
rect -13524 -7452 -13386 -484
rect -13290 -7452 -13152 -484
rect -13056 -7452 -12918 -484
rect -12822 -7452 -12684 -484
rect -12588 -7452 -12450 -484
rect -12354 -7452 -12216 -484
rect -12120 -7452 -11982 -484
rect -11886 -7452 -11748 -484
rect -11652 -7452 -11514 -484
rect -11418 -7452 -11280 -484
rect -11184 -7452 -11046 -484
rect -10950 -7452 -10812 -484
rect -10716 -7452 -10578 -484
rect -10482 -7452 -10344 -484
rect -10248 -7452 -10110 -484
rect -10014 -7452 -9876 -484
rect -9780 -7452 -9642 -484
rect -9546 -7452 -9408 -484
rect -9312 -7452 -9174 -484
rect -9078 -7452 -8940 -484
rect -8844 -7452 -8706 -484
rect -8610 -7452 -8472 -484
rect -8376 -7452 -8238 -484
rect -8142 -7452 -8004 -484
rect -7908 -7452 -7770 -484
rect -7674 -7452 -7536 -484
rect -7440 -7452 -7302 -484
rect -7206 -7452 -7068 -484
rect -6972 -7452 -6834 -484
rect -6738 -7452 -6600 -484
rect -6504 -7452 -6366 -484
rect -6270 -7452 -6132 -484
rect -6036 -7452 -5898 -484
rect -5802 -7452 -5664 -484
rect -5568 -7452 -5430 -484
rect -5334 -7452 -5196 -484
rect -5100 -7452 -4962 -484
rect -4866 -7452 -4728 -484
rect -4632 -7452 -4494 -484
rect -4398 -7452 -4260 -484
rect -4164 -7452 -4026 -484
rect -3930 -7452 -3792 -484
rect -3696 -7452 -3558 -484
rect -3462 -7452 -3324 -484
rect -3228 -7452 -3090 -484
rect -2994 -7452 -2856 -484
rect -2760 -7452 -2622 -484
rect -2526 -7452 -2388 -484
rect -2292 -7452 -2154 -484
rect -2058 -7452 -1920 -484
rect -1824 -7452 -1686 -484
rect -1590 -7452 -1452 -484
rect -1356 -7452 -1218 -484
rect -1122 -7452 -984 -484
rect -888 -7452 -750 -484
rect -654 -7452 -516 -484
rect -420 -7452 -282 -484
rect -186 -7452 -48 -484
rect 48 -7452 186 -484
rect 282 -7452 420 -484
rect 516 -7452 654 -484
rect 750 -7452 888 -484
rect 984 -7452 1122 -484
rect 1218 -7452 1356 -484
rect 1452 -7452 1590 -484
rect 1686 -7452 1824 -484
rect 1920 -7452 2058 -484
rect 2154 -7452 2292 -484
rect 2388 -7452 2526 -484
rect 2622 -7452 2760 -484
rect 2856 -7452 2994 -484
rect 3090 -7452 3228 -484
rect 3324 -7452 3462 -484
rect 3558 -7452 3696 -484
rect 3792 -7452 3930 -484
rect 4026 -7452 4164 -484
rect 4260 -7452 4398 -484
rect 4494 -7452 4632 -484
rect 4728 -7452 4866 -484
rect 4962 -7452 5100 -484
rect 5196 -7452 5334 -484
rect 5430 -7452 5568 -484
rect 5664 -7452 5802 -484
rect 5898 -7452 6036 -484
rect 6132 -7452 6270 -484
rect 6366 -7452 6504 -484
rect 6600 -7452 6738 -484
rect 6834 -7452 6972 -484
rect 7068 -7452 7206 -484
rect 7302 -7452 7440 -484
rect 7536 -7452 7674 -484
rect 7770 -7452 7908 -484
rect 8004 -7452 8142 -484
rect 8238 -7452 8376 -484
rect 8472 -7452 8610 -484
rect 8706 -7452 8844 -484
rect 8940 -7452 9078 -484
rect 9174 -7452 9312 -484
rect 9408 -7452 9546 -484
rect 9642 -7452 9780 -484
rect 9876 -7452 10014 -484
rect 10110 -7452 10248 -484
rect 10344 -7452 10482 -484
rect 10578 -7452 10716 -484
rect 10812 -7452 10950 -484
rect 11046 -7452 11184 -484
rect 11280 -7452 11418 -484
rect 11514 -7452 11652 -484
rect 11748 -7452 11886 -484
rect 11982 -7452 12120 -484
rect 12216 -7452 12354 -484
rect 12450 -7452 12588 -484
rect 12684 -7452 12822 -484
rect 12918 -7452 13056 -484
rect 13152 -7452 13290 -484
rect 13386 -7452 13524 -484
rect 13620 -7452 13758 -484
rect 13854 -7452 13992 -484
rect 14088 -7452 14226 -484
rect 14322 -7452 14460 -484
rect 14556 -7452 14694 -484
rect 14790 -7452 14928 -484
rect 15024 -7452 15162 -484
rect 15258 -7452 15396 -484
rect 15492 -7452 15630 -484
rect 15726 -7452 15864 -484
rect 15960 -7452 16098 -484
rect 16194 -7452 16332 -484
rect 16428 -7452 16566 -484
rect 16662 -7452 16800 -484
rect 16896 -7452 17034 -484
rect 17130 -7452 17268 -484
rect 17364 -7452 17502 -484
rect 17598 -7452 17736 -484
rect 17832 -7452 17970 -484
rect 18066 -7452 18204 -484
rect 18300 -7452 18438 -484
rect 18534 -7452 18672 -484
rect 18768 -7452 18906 -484
rect 19002 -7452 19140 -484
rect 19236 -7452 19374 -484
rect 19470 -7452 19608 -484
rect 19704 -7452 19842 -484
rect 19938 -7452 20076 -484
rect 20172 -7452 20310 -484
rect 20406 -7452 20544 -484
rect 20640 -7452 20778 -484
rect 20874 -7452 21012 -484
rect 21108 -7452 21246 -484
rect 21342 -7452 21480 -484
rect 21576 -7452 21714 -484
rect 21810 -7452 21948 -484
rect 22044 -7452 22182 -484
rect 22278 -7452 22416 -484
rect 22512 -7452 22650 -484
rect 22746 -7452 22884 -484
rect 22980 -7452 23118 -484
rect 23214 -7452 23352 -484
rect 23448 -7452 23586 -484
rect 23682 -7452 23820 -484
rect 23916 -7452 24054 -484
rect 24150 -7452 24288 -484
rect 24384 -7452 24522 -484
rect 24618 -7452 24756 -484
rect 24852 -7452 24990 -484
rect 25086 -7452 25224 -484
rect 25320 -7452 25458 -484
rect 25554 -7452 25692 -484
rect 25788 -7452 25926 -484
rect 26022 -7452 26160 -484
rect 26256 -7452 26394 -484
rect 26490 -7452 26628 -484
rect 26724 -7452 26862 -484
rect 26958 -7452 27096 -484
rect 27192 -7452 27330 -484
rect 27426 -7452 27564 -484
rect 27660 -7452 27798 -484
rect 27894 -7452 28032 -484
rect 28128 -7452 28266 -484
rect 28362 -7452 28500 -484
rect 28596 -7452 28734 -484
rect 28830 -7452 28968 -484
rect 29064 -7452 29202 -484
rect 29298 -7452 29436 -484
rect 29532 -7452 29670 -484
rect 29766 -7452 29904 -484
<< locali >>
rect -30034 7980 -29938 8014
rect 29938 7980 30034 8014
rect -30034 7918 -30000 7980
rect 30000 7918 30034 7980
rect -30034 -7980 -30000 -7918
rect 30000 -7980 30034 -7918
rect -30034 -8014 -29938 -7980
rect 29938 -8014 30034 -7980
<< viali >>
rect -29888 7469 -29782 7866
rect -29654 7469 -29548 7866
rect -29420 7469 -29314 7866
rect -29186 7469 -29080 7866
rect -28952 7469 -28846 7866
rect -28718 7469 -28612 7866
rect -28484 7469 -28378 7866
rect -28250 7469 -28144 7866
rect -28016 7469 -27910 7866
rect -27782 7469 -27676 7866
rect -27548 7469 -27442 7866
rect -27314 7469 -27208 7866
rect -27080 7469 -26974 7866
rect -26846 7469 -26740 7866
rect -26612 7469 -26506 7866
rect -26378 7469 -26272 7866
rect -26144 7469 -26038 7866
rect -25910 7469 -25804 7866
rect -25676 7469 -25570 7866
rect -25442 7469 -25336 7866
rect -25208 7469 -25102 7866
rect -24974 7469 -24868 7866
rect -24740 7469 -24634 7866
rect -24506 7469 -24400 7866
rect -24272 7469 -24166 7866
rect -24038 7469 -23932 7866
rect -23804 7469 -23698 7866
rect -23570 7469 -23464 7866
rect -23336 7469 -23230 7866
rect -23102 7469 -22996 7866
rect -22868 7469 -22762 7866
rect -22634 7469 -22528 7866
rect -22400 7469 -22294 7866
rect -22166 7469 -22060 7866
rect -21932 7469 -21826 7866
rect -21698 7469 -21592 7866
rect -21464 7469 -21358 7866
rect -21230 7469 -21124 7866
rect -20996 7469 -20890 7866
rect -20762 7469 -20656 7866
rect -20528 7469 -20422 7866
rect -20294 7469 -20188 7866
rect -20060 7469 -19954 7866
rect -19826 7469 -19720 7866
rect -19592 7469 -19486 7866
rect -19358 7469 -19252 7866
rect -19124 7469 -19018 7866
rect -18890 7469 -18784 7866
rect -18656 7469 -18550 7866
rect -18422 7469 -18316 7866
rect -18188 7469 -18082 7866
rect -17954 7469 -17848 7866
rect -17720 7469 -17614 7866
rect -17486 7469 -17380 7866
rect -17252 7469 -17146 7866
rect -17018 7469 -16912 7866
rect -16784 7469 -16678 7866
rect -16550 7469 -16444 7866
rect -16316 7469 -16210 7866
rect -16082 7469 -15976 7866
rect -15848 7469 -15742 7866
rect -15614 7469 -15508 7866
rect -15380 7469 -15274 7866
rect -15146 7469 -15040 7866
rect -14912 7469 -14806 7866
rect -14678 7469 -14572 7866
rect -14444 7469 -14338 7866
rect -14210 7469 -14104 7866
rect -13976 7469 -13870 7866
rect -13742 7469 -13636 7866
rect -13508 7469 -13402 7866
rect -13274 7469 -13168 7866
rect -13040 7469 -12934 7866
rect -12806 7469 -12700 7866
rect -12572 7469 -12466 7866
rect -12338 7469 -12232 7866
rect -12104 7469 -11998 7866
rect -11870 7469 -11764 7866
rect -11636 7469 -11530 7866
rect -11402 7469 -11296 7866
rect -11168 7469 -11062 7866
rect -10934 7469 -10828 7866
rect -10700 7469 -10594 7866
rect -10466 7469 -10360 7866
rect -10232 7469 -10126 7866
rect -9998 7469 -9892 7866
rect -9764 7469 -9658 7866
rect -9530 7469 -9424 7866
rect -9296 7469 -9190 7866
rect -9062 7469 -8956 7866
rect -8828 7469 -8722 7866
rect -8594 7469 -8488 7866
rect -8360 7469 -8254 7866
rect -8126 7469 -8020 7866
rect -7892 7469 -7786 7866
rect -7658 7469 -7552 7866
rect -7424 7469 -7318 7866
rect -7190 7469 -7084 7866
rect -6956 7469 -6850 7866
rect -6722 7469 -6616 7866
rect -6488 7469 -6382 7866
rect -6254 7469 -6148 7866
rect -6020 7469 -5914 7866
rect -5786 7469 -5680 7866
rect -5552 7469 -5446 7866
rect -5318 7469 -5212 7866
rect -5084 7469 -4978 7866
rect -4850 7469 -4744 7866
rect -4616 7469 -4510 7866
rect -4382 7469 -4276 7866
rect -4148 7469 -4042 7866
rect -3914 7469 -3808 7866
rect -3680 7469 -3574 7866
rect -3446 7469 -3340 7866
rect -3212 7469 -3106 7866
rect -2978 7469 -2872 7866
rect -2744 7469 -2638 7866
rect -2510 7469 -2404 7866
rect -2276 7469 -2170 7866
rect -2042 7469 -1936 7866
rect -1808 7469 -1702 7866
rect -1574 7469 -1468 7866
rect -1340 7469 -1234 7866
rect -1106 7469 -1000 7866
rect -872 7469 -766 7866
rect -638 7469 -532 7866
rect -404 7469 -298 7866
rect -170 7469 -64 7866
rect 64 7469 170 7866
rect 298 7469 404 7866
rect 532 7469 638 7866
rect 766 7469 872 7866
rect 1000 7469 1106 7866
rect 1234 7469 1340 7866
rect 1468 7469 1574 7866
rect 1702 7469 1808 7866
rect 1936 7469 2042 7866
rect 2170 7469 2276 7866
rect 2404 7469 2510 7866
rect 2638 7469 2744 7866
rect 2872 7469 2978 7866
rect 3106 7469 3212 7866
rect 3340 7469 3446 7866
rect 3574 7469 3680 7866
rect 3808 7469 3914 7866
rect 4042 7469 4148 7866
rect 4276 7469 4382 7866
rect 4510 7469 4616 7866
rect 4744 7469 4850 7866
rect 4978 7469 5084 7866
rect 5212 7469 5318 7866
rect 5446 7469 5552 7866
rect 5680 7469 5786 7866
rect 5914 7469 6020 7866
rect 6148 7469 6254 7866
rect 6382 7469 6488 7866
rect 6616 7469 6722 7866
rect 6850 7469 6956 7866
rect 7084 7469 7190 7866
rect 7318 7469 7424 7866
rect 7552 7469 7658 7866
rect 7786 7469 7892 7866
rect 8020 7469 8126 7866
rect 8254 7469 8360 7866
rect 8488 7469 8594 7866
rect 8722 7469 8828 7866
rect 8956 7469 9062 7866
rect 9190 7469 9296 7866
rect 9424 7469 9530 7866
rect 9658 7469 9764 7866
rect 9892 7469 9998 7866
rect 10126 7469 10232 7866
rect 10360 7469 10466 7866
rect 10594 7469 10700 7866
rect 10828 7469 10934 7866
rect 11062 7469 11168 7866
rect 11296 7469 11402 7866
rect 11530 7469 11636 7866
rect 11764 7469 11870 7866
rect 11998 7469 12104 7866
rect 12232 7469 12338 7866
rect 12466 7469 12572 7866
rect 12700 7469 12806 7866
rect 12934 7469 13040 7866
rect 13168 7469 13274 7866
rect 13402 7469 13508 7866
rect 13636 7469 13742 7866
rect 13870 7469 13976 7866
rect 14104 7469 14210 7866
rect 14338 7469 14444 7866
rect 14572 7469 14678 7866
rect 14806 7469 14912 7866
rect 15040 7469 15146 7866
rect 15274 7469 15380 7866
rect 15508 7469 15614 7866
rect 15742 7469 15848 7866
rect 15976 7469 16082 7866
rect 16210 7469 16316 7866
rect 16444 7469 16550 7866
rect 16678 7469 16784 7866
rect 16912 7469 17018 7866
rect 17146 7469 17252 7866
rect 17380 7469 17486 7866
rect 17614 7469 17720 7866
rect 17848 7469 17954 7866
rect 18082 7469 18188 7866
rect 18316 7469 18422 7866
rect 18550 7469 18656 7866
rect 18784 7469 18890 7866
rect 19018 7469 19124 7866
rect 19252 7469 19358 7866
rect 19486 7469 19592 7866
rect 19720 7469 19826 7866
rect 19954 7469 20060 7866
rect 20188 7469 20294 7866
rect 20422 7469 20528 7866
rect 20656 7469 20762 7866
rect 20890 7469 20996 7866
rect 21124 7469 21230 7866
rect 21358 7469 21464 7866
rect 21592 7469 21698 7866
rect 21826 7469 21932 7866
rect 22060 7469 22166 7866
rect 22294 7469 22400 7866
rect 22528 7469 22634 7866
rect 22762 7469 22868 7866
rect 22996 7469 23102 7866
rect 23230 7469 23336 7866
rect 23464 7469 23570 7866
rect 23698 7469 23804 7866
rect 23932 7469 24038 7866
rect 24166 7469 24272 7866
rect 24400 7469 24506 7866
rect 24634 7469 24740 7866
rect 24868 7469 24974 7866
rect 25102 7469 25208 7866
rect 25336 7469 25442 7866
rect 25570 7469 25676 7866
rect 25804 7469 25910 7866
rect 26038 7469 26144 7866
rect 26272 7469 26378 7866
rect 26506 7469 26612 7866
rect 26740 7469 26846 7866
rect 26974 7469 27080 7866
rect 27208 7469 27314 7866
rect 27442 7469 27548 7866
rect 27676 7469 27782 7866
rect 27910 7469 28016 7866
rect 28144 7469 28250 7866
rect 28378 7469 28484 7866
rect 28612 7469 28718 7866
rect 28846 7469 28952 7866
rect 29080 7469 29186 7866
rect 29314 7469 29420 7866
rect 29548 7469 29654 7866
rect 29782 7469 29888 7866
rect -29888 70 -29782 467
rect -29654 70 -29548 467
rect -29420 70 -29314 467
rect -29186 70 -29080 467
rect -28952 70 -28846 467
rect -28718 70 -28612 467
rect -28484 70 -28378 467
rect -28250 70 -28144 467
rect -28016 70 -27910 467
rect -27782 70 -27676 467
rect -27548 70 -27442 467
rect -27314 70 -27208 467
rect -27080 70 -26974 467
rect -26846 70 -26740 467
rect -26612 70 -26506 467
rect -26378 70 -26272 467
rect -26144 70 -26038 467
rect -25910 70 -25804 467
rect -25676 70 -25570 467
rect -25442 70 -25336 467
rect -25208 70 -25102 467
rect -24974 70 -24868 467
rect -24740 70 -24634 467
rect -24506 70 -24400 467
rect -24272 70 -24166 467
rect -24038 70 -23932 467
rect -23804 70 -23698 467
rect -23570 70 -23464 467
rect -23336 70 -23230 467
rect -23102 70 -22996 467
rect -22868 70 -22762 467
rect -22634 70 -22528 467
rect -22400 70 -22294 467
rect -22166 70 -22060 467
rect -21932 70 -21826 467
rect -21698 70 -21592 467
rect -21464 70 -21358 467
rect -21230 70 -21124 467
rect -20996 70 -20890 467
rect -20762 70 -20656 467
rect -20528 70 -20422 467
rect -20294 70 -20188 467
rect -20060 70 -19954 467
rect -19826 70 -19720 467
rect -19592 70 -19486 467
rect -19358 70 -19252 467
rect -19124 70 -19018 467
rect -18890 70 -18784 467
rect -18656 70 -18550 467
rect -18422 70 -18316 467
rect -18188 70 -18082 467
rect -17954 70 -17848 467
rect -17720 70 -17614 467
rect -17486 70 -17380 467
rect -17252 70 -17146 467
rect -17018 70 -16912 467
rect -16784 70 -16678 467
rect -16550 70 -16444 467
rect -16316 70 -16210 467
rect -16082 70 -15976 467
rect -15848 70 -15742 467
rect -15614 70 -15508 467
rect -15380 70 -15274 467
rect -15146 70 -15040 467
rect -14912 70 -14806 467
rect -14678 70 -14572 467
rect -14444 70 -14338 467
rect -14210 70 -14104 467
rect -13976 70 -13870 467
rect -13742 70 -13636 467
rect -13508 70 -13402 467
rect -13274 70 -13168 467
rect -13040 70 -12934 467
rect -12806 70 -12700 467
rect -12572 70 -12466 467
rect -12338 70 -12232 467
rect -12104 70 -11998 467
rect -11870 70 -11764 467
rect -11636 70 -11530 467
rect -11402 70 -11296 467
rect -11168 70 -11062 467
rect -10934 70 -10828 467
rect -10700 70 -10594 467
rect -10466 70 -10360 467
rect -10232 70 -10126 467
rect -9998 70 -9892 467
rect -9764 70 -9658 467
rect -9530 70 -9424 467
rect -9296 70 -9190 467
rect -9062 70 -8956 467
rect -8828 70 -8722 467
rect -8594 70 -8488 467
rect -8360 70 -8254 467
rect -8126 70 -8020 467
rect -7892 70 -7786 467
rect -7658 70 -7552 467
rect -7424 70 -7318 467
rect -7190 70 -7084 467
rect -6956 70 -6850 467
rect -6722 70 -6616 467
rect -6488 70 -6382 467
rect -6254 70 -6148 467
rect -6020 70 -5914 467
rect -5786 70 -5680 467
rect -5552 70 -5446 467
rect -5318 70 -5212 467
rect -5084 70 -4978 467
rect -4850 70 -4744 467
rect -4616 70 -4510 467
rect -4382 70 -4276 467
rect -4148 70 -4042 467
rect -3914 70 -3808 467
rect -3680 70 -3574 467
rect -3446 70 -3340 467
rect -3212 70 -3106 467
rect -2978 70 -2872 467
rect -2744 70 -2638 467
rect -2510 70 -2404 467
rect -2276 70 -2170 467
rect -2042 70 -1936 467
rect -1808 70 -1702 467
rect -1574 70 -1468 467
rect -1340 70 -1234 467
rect -1106 70 -1000 467
rect -872 70 -766 467
rect -638 70 -532 467
rect -404 70 -298 467
rect -170 70 -64 467
rect 64 70 170 467
rect 298 70 404 467
rect 532 70 638 467
rect 766 70 872 467
rect 1000 70 1106 467
rect 1234 70 1340 467
rect 1468 70 1574 467
rect 1702 70 1808 467
rect 1936 70 2042 467
rect 2170 70 2276 467
rect 2404 70 2510 467
rect 2638 70 2744 467
rect 2872 70 2978 467
rect 3106 70 3212 467
rect 3340 70 3446 467
rect 3574 70 3680 467
rect 3808 70 3914 467
rect 4042 70 4148 467
rect 4276 70 4382 467
rect 4510 70 4616 467
rect 4744 70 4850 467
rect 4978 70 5084 467
rect 5212 70 5318 467
rect 5446 70 5552 467
rect 5680 70 5786 467
rect 5914 70 6020 467
rect 6148 70 6254 467
rect 6382 70 6488 467
rect 6616 70 6722 467
rect 6850 70 6956 467
rect 7084 70 7190 467
rect 7318 70 7424 467
rect 7552 70 7658 467
rect 7786 70 7892 467
rect 8020 70 8126 467
rect 8254 70 8360 467
rect 8488 70 8594 467
rect 8722 70 8828 467
rect 8956 70 9062 467
rect 9190 70 9296 467
rect 9424 70 9530 467
rect 9658 70 9764 467
rect 9892 70 9998 467
rect 10126 70 10232 467
rect 10360 70 10466 467
rect 10594 70 10700 467
rect 10828 70 10934 467
rect 11062 70 11168 467
rect 11296 70 11402 467
rect 11530 70 11636 467
rect 11764 70 11870 467
rect 11998 70 12104 467
rect 12232 70 12338 467
rect 12466 70 12572 467
rect 12700 70 12806 467
rect 12934 70 13040 467
rect 13168 70 13274 467
rect 13402 70 13508 467
rect 13636 70 13742 467
rect 13870 70 13976 467
rect 14104 70 14210 467
rect 14338 70 14444 467
rect 14572 70 14678 467
rect 14806 70 14912 467
rect 15040 70 15146 467
rect 15274 70 15380 467
rect 15508 70 15614 467
rect 15742 70 15848 467
rect 15976 70 16082 467
rect 16210 70 16316 467
rect 16444 70 16550 467
rect 16678 70 16784 467
rect 16912 70 17018 467
rect 17146 70 17252 467
rect 17380 70 17486 467
rect 17614 70 17720 467
rect 17848 70 17954 467
rect 18082 70 18188 467
rect 18316 70 18422 467
rect 18550 70 18656 467
rect 18784 70 18890 467
rect 19018 70 19124 467
rect 19252 70 19358 467
rect 19486 70 19592 467
rect 19720 70 19826 467
rect 19954 70 20060 467
rect 20188 70 20294 467
rect 20422 70 20528 467
rect 20656 70 20762 467
rect 20890 70 20996 467
rect 21124 70 21230 467
rect 21358 70 21464 467
rect 21592 70 21698 467
rect 21826 70 21932 467
rect 22060 70 22166 467
rect 22294 70 22400 467
rect 22528 70 22634 467
rect 22762 70 22868 467
rect 22996 70 23102 467
rect 23230 70 23336 467
rect 23464 70 23570 467
rect 23698 70 23804 467
rect 23932 70 24038 467
rect 24166 70 24272 467
rect 24400 70 24506 467
rect 24634 70 24740 467
rect 24868 70 24974 467
rect 25102 70 25208 467
rect 25336 70 25442 467
rect 25570 70 25676 467
rect 25804 70 25910 467
rect 26038 70 26144 467
rect 26272 70 26378 467
rect 26506 70 26612 467
rect 26740 70 26846 467
rect 26974 70 27080 467
rect 27208 70 27314 467
rect 27442 70 27548 467
rect 27676 70 27782 467
rect 27910 70 28016 467
rect 28144 70 28250 467
rect 28378 70 28484 467
rect 28612 70 28718 467
rect 28846 70 28952 467
rect 29080 70 29186 467
rect 29314 70 29420 467
rect 29548 70 29654 467
rect 29782 70 29888 467
rect -29888 -467 -29782 -70
rect -29654 -467 -29548 -70
rect -29420 -467 -29314 -70
rect -29186 -467 -29080 -70
rect -28952 -467 -28846 -70
rect -28718 -467 -28612 -70
rect -28484 -467 -28378 -70
rect -28250 -467 -28144 -70
rect -28016 -467 -27910 -70
rect -27782 -467 -27676 -70
rect -27548 -467 -27442 -70
rect -27314 -467 -27208 -70
rect -27080 -467 -26974 -70
rect -26846 -467 -26740 -70
rect -26612 -467 -26506 -70
rect -26378 -467 -26272 -70
rect -26144 -467 -26038 -70
rect -25910 -467 -25804 -70
rect -25676 -467 -25570 -70
rect -25442 -467 -25336 -70
rect -25208 -467 -25102 -70
rect -24974 -467 -24868 -70
rect -24740 -467 -24634 -70
rect -24506 -467 -24400 -70
rect -24272 -467 -24166 -70
rect -24038 -467 -23932 -70
rect -23804 -467 -23698 -70
rect -23570 -467 -23464 -70
rect -23336 -467 -23230 -70
rect -23102 -467 -22996 -70
rect -22868 -467 -22762 -70
rect -22634 -467 -22528 -70
rect -22400 -467 -22294 -70
rect -22166 -467 -22060 -70
rect -21932 -467 -21826 -70
rect -21698 -467 -21592 -70
rect -21464 -467 -21358 -70
rect -21230 -467 -21124 -70
rect -20996 -467 -20890 -70
rect -20762 -467 -20656 -70
rect -20528 -467 -20422 -70
rect -20294 -467 -20188 -70
rect -20060 -467 -19954 -70
rect -19826 -467 -19720 -70
rect -19592 -467 -19486 -70
rect -19358 -467 -19252 -70
rect -19124 -467 -19018 -70
rect -18890 -467 -18784 -70
rect -18656 -467 -18550 -70
rect -18422 -467 -18316 -70
rect -18188 -467 -18082 -70
rect -17954 -467 -17848 -70
rect -17720 -467 -17614 -70
rect -17486 -467 -17380 -70
rect -17252 -467 -17146 -70
rect -17018 -467 -16912 -70
rect -16784 -467 -16678 -70
rect -16550 -467 -16444 -70
rect -16316 -467 -16210 -70
rect -16082 -467 -15976 -70
rect -15848 -467 -15742 -70
rect -15614 -467 -15508 -70
rect -15380 -467 -15274 -70
rect -15146 -467 -15040 -70
rect -14912 -467 -14806 -70
rect -14678 -467 -14572 -70
rect -14444 -467 -14338 -70
rect -14210 -467 -14104 -70
rect -13976 -467 -13870 -70
rect -13742 -467 -13636 -70
rect -13508 -467 -13402 -70
rect -13274 -467 -13168 -70
rect -13040 -467 -12934 -70
rect -12806 -467 -12700 -70
rect -12572 -467 -12466 -70
rect -12338 -467 -12232 -70
rect -12104 -467 -11998 -70
rect -11870 -467 -11764 -70
rect -11636 -467 -11530 -70
rect -11402 -467 -11296 -70
rect -11168 -467 -11062 -70
rect -10934 -467 -10828 -70
rect -10700 -467 -10594 -70
rect -10466 -467 -10360 -70
rect -10232 -467 -10126 -70
rect -9998 -467 -9892 -70
rect -9764 -467 -9658 -70
rect -9530 -467 -9424 -70
rect -9296 -467 -9190 -70
rect -9062 -467 -8956 -70
rect -8828 -467 -8722 -70
rect -8594 -467 -8488 -70
rect -8360 -467 -8254 -70
rect -8126 -467 -8020 -70
rect -7892 -467 -7786 -70
rect -7658 -467 -7552 -70
rect -7424 -467 -7318 -70
rect -7190 -467 -7084 -70
rect -6956 -467 -6850 -70
rect -6722 -467 -6616 -70
rect -6488 -467 -6382 -70
rect -6254 -467 -6148 -70
rect -6020 -467 -5914 -70
rect -5786 -467 -5680 -70
rect -5552 -467 -5446 -70
rect -5318 -467 -5212 -70
rect -5084 -467 -4978 -70
rect -4850 -467 -4744 -70
rect -4616 -467 -4510 -70
rect -4382 -467 -4276 -70
rect -4148 -467 -4042 -70
rect -3914 -467 -3808 -70
rect -3680 -467 -3574 -70
rect -3446 -467 -3340 -70
rect -3212 -467 -3106 -70
rect -2978 -467 -2872 -70
rect -2744 -467 -2638 -70
rect -2510 -467 -2404 -70
rect -2276 -467 -2170 -70
rect -2042 -467 -1936 -70
rect -1808 -467 -1702 -70
rect -1574 -467 -1468 -70
rect -1340 -467 -1234 -70
rect -1106 -467 -1000 -70
rect -872 -467 -766 -70
rect -638 -467 -532 -70
rect -404 -467 -298 -70
rect -170 -467 -64 -70
rect 64 -467 170 -70
rect 298 -467 404 -70
rect 532 -467 638 -70
rect 766 -467 872 -70
rect 1000 -467 1106 -70
rect 1234 -467 1340 -70
rect 1468 -467 1574 -70
rect 1702 -467 1808 -70
rect 1936 -467 2042 -70
rect 2170 -467 2276 -70
rect 2404 -467 2510 -70
rect 2638 -467 2744 -70
rect 2872 -467 2978 -70
rect 3106 -467 3212 -70
rect 3340 -467 3446 -70
rect 3574 -467 3680 -70
rect 3808 -467 3914 -70
rect 4042 -467 4148 -70
rect 4276 -467 4382 -70
rect 4510 -467 4616 -70
rect 4744 -467 4850 -70
rect 4978 -467 5084 -70
rect 5212 -467 5318 -70
rect 5446 -467 5552 -70
rect 5680 -467 5786 -70
rect 5914 -467 6020 -70
rect 6148 -467 6254 -70
rect 6382 -467 6488 -70
rect 6616 -467 6722 -70
rect 6850 -467 6956 -70
rect 7084 -467 7190 -70
rect 7318 -467 7424 -70
rect 7552 -467 7658 -70
rect 7786 -467 7892 -70
rect 8020 -467 8126 -70
rect 8254 -467 8360 -70
rect 8488 -467 8594 -70
rect 8722 -467 8828 -70
rect 8956 -467 9062 -70
rect 9190 -467 9296 -70
rect 9424 -467 9530 -70
rect 9658 -467 9764 -70
rect 9892 -467 9998 -70
rect 10126 -467 10232 -70
rect 10360 -467 10466 -70
rect 10594 -467 10700 -70
rect 10828 -467 10934 -70
rect 11062 -467 11168 -70
rect 11296 -467 11402 -70
rect 11530 -467 11636 -70
rect 11764 -467 11870 -70
rect 11998 -467 12104 -70
rect 12232 -467 12338 -70
rect 12466 -467 12572 -70
rect 12700 -467 12806 -70
rect 12934 -467 13040 -70
rect 13168 -467 13274 -70
rect 13402 -467 13508 -70
rect 13636 -467 13742 -70
rect 13870 -467 13976 -70
rect 14104 -467 14210 -70
rect 14338 -467 14444 -70
rect 14572 -467 14678 -70
rect 14806 -467 14912 -70
rect 15040 -467 15146 -70
rect 15274 -467 15380 -70
rect 15508 -467 15614 -70
rect 15742 -467 15848 -70
rect 15976 -467 16082 -70
rect 16210 -467 16316 -70
rect 16444 -467 16550 -70
rect 16678 -467 16784 -70
rect 16912 -467 17018 -70
rect 17146 -467 17252 -70
rect 17380 -467 17486 -70
rect 17614 -467 17720 -70
rect 17848 -467 17954 -70
rect 18082 -467 18188 -70
rect 18316 -467 18422 -70
rect 18550 -467 18656 -70
rect 18784 -467 18890 -70
rect 19018 -467 19124 -70
rect 19252 -467 19358 -70
rect 19486 -467 19592 -70
rect 19720 -467 19826 -70
rect 19954 -467 20060 -70
rect 20188 -467 20294 -70
rect 20422 -467 20528 -70
rect 20656 -467 20762 -70
rect 20890 -467 20996 -70
rect 21124 -467 21230 -70
rect 21358 -467 21464 -70
rect 21592 -467 21698 -70
rect 21826 -467 21932 -70
rect 22060 -467 22166 -70
rect 22294 -467 22400 -70
rect 22528 -467 22634 -70
rect 22762 -467 22868 -70
rect 22996 -467 23102 -70
rect 23230 -467 23336 -70
rect 23464 -467 23570 -70
rect 23698 -467 23804 -70
rect 23932 -467 24038 -70
rect 24166 -467 24272 -70
rect 24400 -467 24506 -70
rect 24634 -467 24740 -70
rect 24868 -467 24974 -70
rect 25102 -467 25208 -70
rect 25336 -467 25442 -70
rect 25570 -467 25676 -70
rect 25804 -467 25910 -70
rect 26038 -467 26144 -70
rect 26272 -467 26378 -70
rect 26506 -467 26612 -70
rect 26740 -467 26846 -70
rect 26974 -467 27080 -70
rect 27208 -467 27314 -70
rect 27442 -467 27548 -70
rect 27676 -467 27782 -70
rect 27910 -467 28016 -70
rect 28144 -467 28250 -70
rect 28378 -467 28484 -70
rect 28612 -467 28718 -70
rect 28846 -467 28952 -70
rect 29080 -467 29186 -70
rect 29314 -467 29420 -70
rect 29548 -467 29654 -70
rect 29782 -467 29888 -70
rect -29888 -7866 -29782 -7469
rect -29654 -7866 -29548 -7469
rect -29420 -7866 -29314 -7469
rect -29186 -7866 -29080 -7469
rect -28952 -7866 -28846 -7469
rect -28718 -7866 -28612 -7469
rect -28484 -7866 -28378 -7469
rect -28250 -7866 -28144 -7469
rect -28016 -7866 -27910 -7469
rect -27782 -7866 -27676 -7469
rect -27548 -7866 -27442 -7469
rect -27314 -7866 -27208 -7469
rect -27080 -7866 -26974 -7469
rect -26846 -7866 -26740 -7469
rect -26612 -7866 -26506 -7469
rect -26378 -7866 -26272 -7469
rect -26144 -7866 -26038 -7469
rect -25910 -7866 -25804 -7469
rect -25676 -7866 -25570 -7469
rect -25442 -7866 -25336 -7469
rect -25208 -7866 -25102 -7469
rect -24974 -7866 -24868 -7469
rect -24740 -7866 -24634 -7469
rect -24506 -7866 -24400 -7469
rect -24272 -7866 -24166 -7469
rect -24038 -7866 -23932 -7469
rect -23804 -7866 -23698 -7469
rect -23570 -7866 -23464 -7469
rect -23336 -7866 -23230 -7469
rect -23102 -7866 -22996 -7469
rect -22868 -7866 -22762 -7469
rect -22634 -7866 -22528 -7469
rect -22400 -7866 -22294 -7469
rect -22166 -7866 -22060 -7469
rect -21932 -7866 -21826 -7469
rect -21698 -7866 -21592 -7469
rect -21464 -7866 -21358 -7469
rect -21230 -7866 -21124 -7469
rect -20996 -7866 -20890 -7469
rect -20762 -7866 -20656 -7469
rect -20528 -7866 -20422 -7469
rect -20294 -7866 -20188 -7469
rect -20060 -7866 -19954 -7469
rect -19826 -7866 -19720 -7469
rect -19592 -7866 -19486 -7469
rect -19358 -7866 -19252 -7469
rect -19124 -7866 -19018 -7469
rect -18890 -7866 -18784 -7469
rect -18656 -7866 -18550 -7469
rect -18422 -7866 -18316 -7469
rect -18188 -7866 -18082 -7469
rect -17954 -7866 -17848 -7469
rect -17720 -7866 -17614 -7469
rect -17486 -7866 -17380 -7469
rect -17252 -7866 -17146 -7469
rect -17018 -7866 -16912 -7469
rect -16784 -7866 -16678 -7469
rect -16550 -7866 -16444 -7469
rect -16316 -7866 -16210 -7469
rect -16082 -7866 -15976 -7469
rect -15848 -7866 -15742 -7469
rect -15614 -7866 -15508 -7469
rect -15380 -7866 -15274 -7469
rect -15146 -7866 -15040 -7469
rect -14912 -7866 -14806 -7469
rect -14678 -7866 -14572 -7469
rect -14444 -7866 -14338 -7469
rect -14210 -7866 -14104 -7469
rect -13976 -7866 -13870 -7469
rect -13742 -7866 -13636 -7469
rect -13508 -7866 -13402 -7469
rect -13274 -7866 -13168 -7469
rect -13040 -7866 -12934 -7469
rect -12806 -7866 -12700 -7469
rect -12572 -7866 -12466 -7469
rect -12338 -7866 -12232 -7469
rect -12104 -7866 -11998 -7469
rect -11870 -7866 -11764 -7469
rect -11636 -7866 -11530 -7469
rect -11402 -7866 -11296 -7469
rect -11168 -7866 -11062 -7469
rect -10934 -7866 -10828 -7469
rect -10700 -7866 -10594 -7469
rect -10466 -7866 -10360 -7469
rect -10232 -7866 -10126 -7469
rect -9998 -7866 -9892 -7469
rect -9764 -7866 -9658 -7469
rect -9530 -7866 -9424 -7469
rect -9296 -7866 -9190 -7469
rect -9062 -7866 -8956 -7469
rect -8828 -7866 -8722 -7469
rect -8594 -7866 -8488 -7469
rect -8360 -7866 -8254 -7469
rect -8126 -7866 -8020 -7469
rect -7892 -7866 -7786 -7469
rect -7658 -7866 -7552 -7469
rect -7424 -7866 -7318 -7469
rect -7190 -7866 -7084 -7469
rect -6956 -7866 -6850 -7469
rect -6722 -7866 -6616 -7469
rect -6488 -7866 -6382 -7469
rect -6254 -7866 -6148 -7469
rect -6020 -7866 -5914 -7469
rect -5786 -7866 -5680 -7469
rect -5552 -7866 -5446 -7469
rect -5318 -7866 -5212 -7469
rect -5084 -7866 -4978 -7469
rect -4850 -7866 -4744 -7469
rect -4616 -7866 -4510 -7469
rect -4382 -7866 -4276 -7469
rect -4148 -7866 -4042 -7469
rect -3914 -7866 -3808 -7469
rect -3680 -7866 -3574 -7469
rect -3446 -7866 -3340 -7469
rect -3212 -7866 -3106 -7469
rect -2978 -7866 -2872 -7469
rect -2744 -7866 -2638 -7469
rect -2510 -7866 -2404 -7469
rect -2276 -7866 -2170 -7469
rect -2042 -7866 -1936 -7469
rect -1808 -7866 -1702 -7469
rect -1574 -7866 -1468 -7469
rect -1340 -7866 -1234 -7469
rect -1106 -7866 -1000 -7469
rect -872 -7866 -766 -7469
rect -638 -7866 -532 -7469
rect -404 -7866 -298 -7469
rect -170 -7866 -64 -7469
rect 64 -7866 170 -7469
rect 298 -7866 404 -7469
rect 532 -7866 638 -7469
rect 766 -7866 872 -7469
rect 1000 -7866 1106 -7469
rect 1234 -7866 1340 -7469
rect 1468 -7866 1574 -7469
rect 1702 -7866 1808 -7469
rect 1936 -7866 2042 -7469
rect 2170 -7866 2276 -7469
rect 2404 -7866 2510 -7469
rect 2638 -7866 2744 -7469
rect 2872 -7866 2978 -7469
rect 3106 -7866 3212 -7469
rect 3340 -7866 3446 -7469
rect 3574 -7866 3680 -7469
rect 3808 -7866 3914 -7469
rect 4042 -7866 4148 -7469
rect 4276 -7866 4382 -7469
rect 4510 -7866 4616 -7469
rect 4744 -7866 4850 -7469
rect 4978 -7866 5084 -7469
rect 5212 -7866 5318 -7469
rect 5446 -7866 5552 -7469
rect 5680 -7866 5786 -7469
rect 5914 -7866 6020 -7469
rect 6148 -7866 6254 -7469
rect 6382 -7866 6488 -7469
rect 6616 -7866 6722 -7469
rect 6850 -7866 6956 -7469
rect 7084 -7866 7190 -7469
rect 7318 -7866 7424 -7469
rect 7552 -7866 7658 -7469
rect 7786 -7866 7892 -7469
rect 8020 -7866 8126 -7469
rect 8254 -7866 8360 -7469
rect 8488 -7866 8594 -7469
rect 8722 -7866 8828 -7469
rect 8956 -7866 9062 -7469
rect 9190 -7866 9296 -7469
rect 9424 -7866 9530 -7469
rect 9658 -7866 9764 -7469
rect 9892 -7866 9998 -7469
rect 10126 -7866 10232 -7469
rect 10360 -7866 10466 -7469
rect 10594 -7866 10700 -7469
rect 10828 -7866 10934 -7469
rect 11062 -7866 11168 -7469
rect 11296 -7866 11402 -7469
rect 11530 -7866 11636 -7469
rect 11764 -7866 11870 -7469
rect 11998 -7866 12104 -7469
rect 12232 -7866 12338 -7469
rect 12466 -7866 12572 -7469
rect 12700 -7866 12806 -7469
rect 12934 -7866 13040 -7469
rect 13168 -7866 13274 -7469
rect 13402 -7866 13508 -7469
rect 13636 -7866 13742 -7469
rect 13870 -7866 13976 -7469
rect 14104 -7866 14210 -7469
rect 14338 -7866 14444 -7469
rect 14572 -7866 14678 -7469
rect 14806 -7866 14912 -7469
rect 15040 -7866 15146 -7469
rect 15274 -7866 15380 -7469
rect 15508 -7866 15614 -7469
rect 15742 -7866 15848 -7469
rect 15976 -7866 16082 -7469
rect 16210 -7866 16316 -7469
rect 16444 -7866 16550 -7469
rect 16678 -7866 16784 -7469
rect 16912 -7866 17018 -7469
rect 17146 -7866 17252 -7469
rect 17380 -7866 17486 -7469
rect 17614 -7866 17720 -7469
rect 17848 -7866 17954 -7469
rect 18082 -7866 18188 -7469
rect 18316 -7866 18422 -7469
rect 18550 -7866 18656 -7469
rect 18784 -7866 18890 -7469
rect 19018 -7866 19124 -7469
rect 19252 -7866 19358 -7469
rect 19486 -7866 19592 -7469
rect 19720 -7866 19826 -7469
rect 19954 -7866 20060 -7469
rect 20188 -7866 20294 -7469
rect 20422 -7866 20528 -7469
rect 20656 -7866 20762 -7469
rect 20890 -7866 20996 -7469
rect 21124 -7866 21230 -7469
rect 21358 -7866 21464 -7469
rect 21592 -7866 21698 -7469
rect 21826 -7866 21932 -7469
rect 22060 -7866 22166 -7469
rect 22294 -7866 22400 -7469
rect 22528 -7866 22634 -7469
rect 22762 -7866 22868 -7469
rect 22996 -7866 23102 -7469
rect 23230 -7866 23336 -7469
rect 23464 -7866 23570 -7469
rect 23698 -7866 23804 -7469
rect 23932 -7866 24038 -7469
rect 24166 -7866 24272 -7469
rect 24400 -7866 24506 -7469
rect 24634 -7866 24740 -7469
rect 24868 -7866 24974 -7469
rect 25102 -7866 25208 -7469
rect 25336 -7866 25442 -7469
rect 25570 -7866 25676 -7469
rect 25804 -7866 25910 -7469
rect 26038 -7866 26144 -7469
rect 26272 -7866 26378 -7469
rect 26506 -7866 26612 -7469
rect 26740 -7866 26846 -7469
rect 26974 -7866 27080 -7469
rect 27208 -7866 27314 -7469
rect 27442 -7866 27548 -7469
rect 27676 -7866 27782 -7469
rect 27910 -7866 28016 -7469
rect 28144 -7866 28250 -7469
rect 28378 -7866 28484 -7469
rect 28612 -7866 28718 -7469
rect 28846 -7866 28952 -7469
rect 29080 -7866 29186 -7469
rect 29314 -7866 29420 -7469
rect 29548 -7866 29654 -7469
rect 29782 -7866 29888 -7469
<< metal1 >>
rect -29894 7866 -29776 7878
rect -29894 7469 -29888 7866
rect -29782 7469 -29776 7866
rect -29894 7457 -29776 7469
rect -29660 7866 -29542 7878
rect -29660 7469 -29654 7866
rect -29548 7469 -29542 7866
rect -29660 7457 -29542 7469
rect -29426 7866 -29308 7878
rect -29426 7469 -29420 7866
rect -29314 7469 -29308 7866
rect -29426 7457 -29308 7469
rect -29192 7866 -29074 7878
rect -29192 7469 -29186 7866
rect -29080 7469 -29074 7866
rect -29192 7457 -29074 7469
rect -28958 7866 -28840 7878
rect -28958 7469 -28952 7866
rect -28846 7469 -28840 7866
rect -28958 7457 -28840 7469
rect -28724 7866 -28606 7878
rect -28724 7469 -28718 7866
rect -28612 7469 -28606 7866
rect -28724 7457 -28606 7469
rect -28490 7866 -28372 7878
rect -28490 7469 -28484 7866
rect -28378 7469 -28372 7866
rect -28490 7457 -28372 7469
rect -28256 7866 -28138 7878
rect -28256 7469 -28250 7866
rect -28144 7469 -28138 7866
rect -28256 7457 -28138 7469
rect -28022 7866 -27904 7878
rect -28022 7469 -28016 7866
rect -27910 7469 -27904 7866
rect -28022 7457 -27904 7469
rect -27788 7866 -27670 7878
rect -27788 7469 -27782 7866
rect -27676 7469 -27670 7866
rect -27788 7457 -27670 7469
rect -27554 7866 -27436 7878
rect -27554 7469 -27548 7866
rect -27442 7469 -27436 7866
rect -27554 7457 -27436 7469
rect -27320 7866 -27202 7878
rect -27320 7469 -27314 7866
rect -27208 7469 -27202 7866
rect -27320 7457 -27202 7469
rect -27086 7866 -26968 7878
rect -27086 7469 -27080 7866
rect -26974 7469 -26968 7866
rect -27086 7457 -26968 7469
rect -26852 7866 -26734 7878
rect -26852 7469 -26846 7866
rect -26740 7469 -26734 7866
rect -26852 7457 -26734 7469
rect -26618 7866 -26500 7878
rect -26618 7469 -26612 7866
rect -26506 7469 -26500 7866
rect -26618 7457 -26500 7469
rect -26384 7866 -26266 7878
rect -26384 7469 -26378 7866
rect -26272 7469 -26266 7866
rect -26384 7457 -26266 7469
rect -26150 7866 -26032 7878
rect -26150 7469 -26144 7866
rect -26038 7469 -26032 7866
rect -26150 7457 -26032 7469
rect -25916 7866 -25798 7878
rect -25916 7469 -25910 7866
rect -25804 7469 -25798 7866
rect -25916 7457 -25798 7469
rect -25682 7866 -25564 7878
rect -25682 7469 -25676 7866
rect -25570 7469 -25564 7866
rect -25682 7457 -25564 7469
rect -25448 7866 -25330 7878
rect -25448 7469 -25442 7866
rect -25336 7469 -25330 7866
rect -25448 7457 -25330 7469
rect -25214 7866 -25096 7878
rect -25214 7469 -25208 7866
rect -25102 7469 -25096 7866
rect -25214 7457 -25096 7469
rect -24980 7866 -24862 7878
rect -24980 7469 -24974 7866
rect -24868 7469 -24862 7866
rect -24980 7457 -24862 7469
rect -24746 7866 -24628 7878
rect -24746 7469 -24740 7866
rect -24634 7469 -24628 7866
rect -24746 7457 -24628 7469
rect -24512 7866 -24394 7878
rect -24512 7469 -24506 7866
rect -24400 7469 -24394 7866
rect -24512 7457 -24394 7469
rect -24278 7866 -24160 7878
rect -24278 7469 -24272 7866
rect -24166 7469 -24160 7866
rect -24278 7457 -24160 7469
rect -24044 7866 -23926 7878
rect -24044 7469 -24038 7866
rect -23932 7469 -23926 7866
rect -24044 7457 -23926 7469
rect -23810 7866 -23692 7878
rect -23810 7469 -23804 7866
rect -23698 7469 -23692 7866
rect -23810 7457 -23692 7469
rect -23576 7866 -23458 7878
rect -23576 7469 -23570 7866
rect -23464 7469 -23458 7866
rect -23576 7457 -23458 7469
rect -23342 7866 -23224 7878
rect -23342 7469 -23336 7866
rect -23230 7469 -23224 7866
rect -23342 7457 -23224 7469
rect -23108 7866 -22990 7878
rect -23108 7469 -23102 7866
rect -22996 7469 -22990 7866
rect -23108 7457 -22990 7469
rect -22874 7866 -22756 7878
rect -22874 7469 -22868 7866
rect -22762 7469 -22756 7866
rect -22874 7457 -22756 7469
rect -22640 7866 -22522 7878
rect -22640 7469 -22634 7866
rect -22528 7469 -22522 7866
rect -22640 7457 -22522 7469
rect -22406 7866 -22288 7878
rect -22406 7469 -22400 7866
rect -22294 7469 -22288 7866
rect -22406 7457 -22288 7469
rect -22172 7866 -22054 7878
rect -22172 7469 -22166 7866
rect -22060 7469 -22054 7866
rect -22172 7457 -22054 7469
rect -21938 7866 -21820 7878
rect -21938 7469 -21932 7866
rect -21826 7469 -21820 7866
rect -21938 7457 -21820 7469
rect -21704 7866 -21586 7878
rect -21704 7469 -21698 7866
rect -21592 7469 -21586 7866
rect -21704 7457 -21586 7469
rect -21470 7866 -21352 7878
rect -21470 7469 -21464 7866
rect -21358 7469 -21352 7866
rect -21470 7457 -21352 7469
rect -21236 7866 -21118 7878
rect -21236 7469 -21230 7866
rect -21124 7469 -21118 7866
rect -21236 7457 -21118 7469
rect -21002 7866 -20884 7878
rect -21002 7469 -20996 7866
rect -20890 7469 -20884 7866
rect -21002 7457 -20884 7469
rect -20768 7866 -20650 7878
rect -20768 7469 -20762 7866
rect -20656 7469 -20650 7866
rect -20768 7457 -20650 7469
rect -20534 7866 -20416 7878
rect -20534 7469 -20528 7866
rect -20422 7469 -20416 7866
rect -20534 7457 -20416 7469
rect -20300 7866 -20182 7878
rect -20300 7469 -20294 7866
rect -20188 7469 -20182 7866
rect -20300 7457 -20182 7469
rect -20066 7866 -19948 7878
rect -20066 7469 -20060 7866
rect -19954 7469 -19948 7866
rect -20066 7457 -19948 7469
rect -19832 7866 -19714 7878
rect -19832 7469 -19826 7866
rect -19720 7469 -19714 7866
rect -19832 7457 -19714 7469
rect -19598 7866 -19480 7878
rect -19598 7469 -19592 7866
rect -19486 7469 -19480 7866
rect -19598 7457 -19480 7469
rect -19364 7866 -19246 7878
rect -19364 7469 -19358 7866
rect -19252 7469 -19246 7866
rect -19364 7457 -19246 7469
rect -19130 7866 -19012 7878
rect -19130 7469 -19124 7866
rect -19018 7469 -19012 7866
rect -19130 7457 -19012 7469
rect -18896 7866 -18778 7878
rect -18896 7469 -18890 7866
rect -18784 7469 -18778 7866
rect -18896 7457 -18778 7469
rect -18662 7866 -18544 7878
rect -18662 7469 -18656 7866
rect -18550 7469 -18544 7866
rect -18662 7457 -18544 7469
rect -18428 7866 -18310 7878
rect -18428 7469 -18422 7866
rect -18316 7469 -18310 7866
rect -18428 7457 -18310 7469
rect -18194 7866 -18076 7878
rect -18194 7469 -18188 7866
rect -18082 7469 -18076 7866
rect -18194 7457 -18076 7469
rect -17960 7866 -17842 7878
rect -17960 7469 -17954 7866
rect -17848 7469 -17842 7866
rect -17960 7457 -17842 7469
rect -17726 7866 -17608 7878
rect -17726 7469 -17720 7866
rect -17614 7469 -17608 7866
rect -17726 7457 -17608 7469
rect -17492 7866 -17374 7878
rect -17492 7469 -17486 7866
rect -17380 7469 -17374 7866
rect -17492 7457 -17374 7469
rect -17258 7866 -17140 7878
rect -17258 7469 -17252 7866
rect -17146 7469 -17140 7866
rect -17258 7457 -17140 7469
rect -17024 7866 -16906 7878
rect -17024 7469 -17018 7866
rect -16912 7469 -16906 7866
rect -17024 7457 -16906 7469
rect -16790 7866 -16672 7878
rect -16790 7469 -16784 7866
rect -16678 7469 -16672 7866
rect -16790 7457 -16672 7469
rect -16556 7866 -16438 7878
rect -16556 7469 -16550 7866
rect -16444 7469 -16438 7866
rect -16556 7457 -16438 7469
rect -16322 7866 -16204 7878
rect -16322 7469 -16316 7866
rect -16210 7469 -16204 7866
rect -16322 7457 -16204 7469
rect -16088 7866 -15970 7878
rect -16088 7469 -16082 7866
rect -15976 7469 -15970 7866
rect -16088 7457 -15970 7469
rect -15854 7866 -15736 7878
rect -15854 7469 -15848 7866
rect -15742 7469 -15736 7866
rect -15854 7457 -15736 7469
rect -15620 7866 -15502 7878
rect -15620 7469 -15614 7866
rect -15508 7469 -15502 7866
rect -15620 7457 -15502 7469
rect -15386 7866 -15268 7878
rect -15386 7469 -15380 7866
rect -15274 7469 -15268 7866
rect -15386 7457 -15268 7469
rect -15152 7866 -15034 7878
rect -15152 7469 -15146 7866
rect -15040 7469 -15034 7866
rect -15152 7457 -15034 7469
rect -14918 7866 -14800 7878
rect -14918 7469 -14912 7866
rect -14806 7469 -14800 7866
rect -14918 7457 -14800 7469
rect -14684 7866 -14566 7878
rect -14684 7469 -14678 7866
rect -14572 7469 -14566 7866
rect -14684 7457 -14566 7469
rect -14450 7866 -14332 7878
rect -14450 7469 -14444 7866
rect -14338 7469 -14332 7866
rect -14450 7457 -14332 7469
rect -14216 7866 -14098 7878
rect -14216 7469 -14210 7866
rect -14104 7469 -14098 7866
rect -14216 7457 -14098 7469
rect -13982 7866 -13864 7878
rect -13982 7469 -13976 7866
rect -13870 7469 -13864 7866
rect -13982 7457 -13864 7469
rect -13748 7866 -13630 7878
rect -13748 7469 -13742 7866
rect -13636 7469 -13630 7866
rect -13748 7457 -13630 7469
rect -13514 7866 -13396 7878
rect -13514 7469 -13508 7866
rect -13402 7469 -13396 7866
rect -13514 7457 -13396 7469
rect -13280 7866 -13162 7878
rect -13280 7469 -13274 7866
rect -13168 7469 -13162 7866
rect -13280 7457 -13162 7469
rect -13046 7866 -12928 7878
rect -13046 7469 -13040 7866
rect -12934 7469 -12928 7866
rect -13046 7457 -12928 7469
rect -12812 7866 -12694 7878
rect -12812 7469 -12806 7866
rect -12700 7469 -12694 7866
rect -12812 7457 -12694 7469
rect -12578 7866 -12460 7878
rect -12578 7469 -12572 7866
rect -12466 7469 -12460 7866
rect -12578 7457 -12460 7469
rect -12344 7866 -12226 7878
rect -12344 7469 -12338 7866
rect -12232 7469 -12226 7866
rect -12344 7457 -12226 7469
rect -12110 7866 -11992 7878
rect -12110 7469 -12104 7866
rect -11998 7469 -11992 7866
rect -12110 7457 -11992 7469
rect -11876 7866 -11758 7878
rect -11876 7469 -11870 7866
rect -11764 7469 -11758 7866
rect -11876 7457 -11758 7469
rect -11642 7866 -11524 7878
rect -11642 7469 -11636 7866
rect -11530 7469 -11524 7866
rect -11642 7457 -11524 7469
rect -11408 7866 -11290 7878
rect -11408 7469 -11402 7866
rect -11296 7469 -11290 7866
rect -11408 7457 -11290 7469
rect -11174 7866 -11056 7878
rect -11174 7469 -11168 7866
rect -11062 7469 -11056 7866
rect -11174 7457 -11056 7469
rect -10940 7866 -10822 7878
rect -10940 7469 -10934 7866
rect -10828 7469 -10822 7866
rect -10940 7457 -10822 7469
rect -10706 7866 -10588 7878
rect -10706 7469 -10700 7866
rect -10594 7469 -10588 7866
rect -10706 7457 -10588 7469
rect -10472 7866 -10354 7878
rect -10472 7469 -10466 7866
rect -10360 7469 -10354 7866
rect -10472 7457 -10354 7469
rect -10238 7866 -10120 7878
rect -10238 7469 -10232 7866
rect -10126 7469 -10120 7866
rect -10238 7457 -10120 7469
rect -10004 7866 -9886 7878
rect -10004 7469 -9998 7866
rect -9892 7469 -9886 7866
rect -10004 7457 -9886 7469
rect -9770 7866 -9652 7878
rect -9770 7469 -9764 7866
rect -9658 7469 -9652 7866
rect -9770 7457 -9652 7469
rect -9536 7866 -9418 7878
rect -9536 7469 -9530 7866
rect -9424 7469 -9418 7866
rect -9536 7457 -9418 7469
rect -9302 7866 -9184 7878
rect -9302 7469 -9296 7866
rect -9190 7469 -9184 7866
rect -9302 7457 -9184 7469
rect -9068 7866 -8950 7878
rect -9068 7469 -9062 7866
rect -8956 7469 -8950 7866
rect -9068 7457 -8950 7469
rect -8834 7866 -8716 7878
rect -8834 7469 -8828 7866
rect -8722 7469 -8716 7866
rect -8834 7457 -8716 7469
rect -8600 7866 -8482 7878
rect -8600 7469 -8594 7866
rect -8488 7469 -8482 7866
rect -8600 7457 -8482 7469
rect -8366 7866 -8248 7878
rect -8366 7469 -8360 7866
rect -8254 7469 -8248 7866
rect -8366 7457 -8248 7469
rect -8132 7866 -8014 7878
rect -8132 7469 -8126 7866
rect -8020 7469 -8014 7866
rect -8132 7457 -8014 7469
rect -7898 7866 -7780 7878
rect -7898 7469 -7892 7866
rect -7786 7469 -7780 7866
rect -7898 7457 -7780 7469
rect -7664 7866 -7546 7878
rect -7664 7469 -7658 7866
rect -7552 7469 -7546 7866
rect -7664 7457 -7546 7469
rect -7430 7866 -7312 7878
rect -7430 7469 -7424 7866
rect -7318 7469 -7312 7866
rect -7430 7457 -7312 7469
rect -7196 7866 -7078 7878
rect -7196 7469 -7190 7866
rect -7084 7469 -7078 7866
rect -7196 7457 -7078 7469
rect -6962 7866 -6844 7878
rect -6962 7469 -6956 7866
rect -6850 7469 -6844 7866
rect -6962 7457 -6844 7469
rect -6728 7866 -6610 7878
rect -6728 7469 -6722 7866
rect -6616 7469 -6610 7866
rect -6728 7457 -6610 7469
rect -6494 7866 -6376 7878
rect -6494 7469 -6488 7866
rect -6382 7469 -6376 7866
rect -6494 7457 -6376 7469
rect -6260 7866 -6142 7878
rect -6260 7469 -6254 7866
rect -6148 7469 -6142 7866
rect -6260 7457 -6142 7469
rect -6026 7866 -5908 7878
rect -6026 7469 -6020 7866
rect -5914 7469 -5908 7866
rect -6026 7457 -5908 7469
rect -5792 7866 -5674 7878
rect -5792 7469 -5786 7866
rect -5680 7469 -5674 7866
rect -5792 7457 -5674 7469
rect -5558 7866 -5440 7878
rect -5558 7469 -5552 7866
rect -5446 7469 -5440 7866
rect -5558 7457 -5440 7469
rect -5324 7866 -5206 7878
rect -5324 7469 -5318 7866
rect -5212 7469 -5206 7866
rect -5324 7457 -5206 7469
rect -5090 7866 -4972 7878
rect -5090 7469 -5084 7866
rect -4978 7469 -4972 7866
rect -5090 7457 -4972 7469
rect -4856 7866 -4738 7878
rect -4856 7469 -4850 7866
rect -4744 7469 -4738 7866
rect -4856 7457 -4738 7469
rect -4622 7866 -4504 7878
rect -4622 7469 -4616 7866
rect -4510 7469 -4504 7866
rect -4622 7457 -4504 7469
rect -4388 7866 -4270 7878
rect -4388 7469 -4382 7866
rect -4276 7469 -4270 7866
rect -4388 7457 -4270 7469
rect -4154 7866 -4036 7878
rect -4154 7469 -4148 7866
rect -4042 7469 -4036 7866
rect -4154 7457 -4036 7469
rect -3920 7866 -3802 7878
rect -3920 7469 -3914 7866
rect -3808 7469 -3802 7866
rect -3920 7457 -3802 7469
rect -3686 7866 -3568 7878
rect -3686 7469 -3680 7866
rect -3574 7469 -3568 7866
rect -3686 7457 -3568 7469
rect -3452 7866 -3334 7878
rect -3452 7469 -3446 7866
rect -3340 7469 -3334 7866
rect -3452 7457 -3334 7469
rect -3218 7866 -3100 7878
rect -3218 7469 -3212 7866
rect -3106 7469 -3100 7866
rect -3218 7457 -3100 7469
rect -2984 7866 -2866 7878
rect -2984 7469 -2978 7866
rect -2872 7469 -2866 7866
rect -2984 7457 -2866 7469
rect -2750 7866 -2632 7878
rect -2750 7469 -2744 7866
rect -2638 7469 -2632 7866
rect -2750 7457 -2632 7469
rect -2516 7866 -2398 7878
rect -2516 7469 -2510 7866
rect -2404 7469 -2398 7866
rect -2516 7457 -2398 7469
rect -2282 7866 -2164 7878
rect -2282 7469 -2276 7866
rect -2170 7469 -2164 7866
rect -2282 7457 -2164 7469
rect -2048 7866 -1930 7878
rect -2048 7469 -2042 7866
rect -1936 7469 -1930 7866
rect -2048 7457 -1930 7469
rect -1814 7866 -1696 7878
rect -1814 7469 -1808 7866
rect -1702 7469 -1696 7866
rect -1814 7457 -1696 7469
rect -1580 7866 -1462 7878
rect -1580 7469 -1574 7866
rect -1468 7469 -1462 7866
rect -1580 7457 -1462 7469
rect -1346 7866 -1228 7878
rect -1346 7469 -1340 7866
rect -1234 7469 -1228 7866
rect -1346 7457 -1228 7469
rect -1112 7866 -994 7878
rect -1112 7469 -1106 7866
rect -1000 7469 -994 7866
rect -1112 7457 -994 7469
rect -878 7866 -760 7878
rect -878 7469 -872 7866
rect -766 7469 -760 7866
rect -878 7457 -760 7469
rect -644 7866 -526 7878
rect -644 7469 -638 7866
rect -532 7469 -526 7866
rect -644 7457 -526 7469
rect -410 7866 -292 7878
rect -410 7469 -404 7866
rect -298 7469 -292 7866
rect -410 7457 -292 7469
rect -176 7866 -58 7878
rect -176 7469 -170 7866
rect -64 7469 -58 7866
rect -176 7457 -58 7469
rect 58 7866 176 7878
rect 58 7469 64 7866
rect 170 7469 176 7866
rect 58 7457 176 7469
rect 292 7866 410 7878
rect 292 7469 298 7866
rect 404 7469 410 7866
rect 292 7457 410 7469
rect 526 7866 644 7878
rect 526 7469 532 7866
rect 638 7469 644 7866
rect 526 7457 644 7469
rect 760 7866 878 7878
rect 760 7469 766 7866
rect 872 7469 878 7866
rect 760 7457 878 7469
rect 994 7866 1112 7878
rect 994 7469 1000 7866
rect 1106 7469 1112 7866
rect 994 7457 1112 7469
rect 1228 7866 1346 7878
rect 1228 7469 1234 7866
rect 1340 7469 1346 7866
rect 1228 7457 1346 7469
rect 1462 7866 1580 7878
rect 1462 7469 1468 7866
rect 1574 7469 1580 7866
rect 1462 7457 1580 7469
rect 1696 7866 1814 7878
rect 1696 7469 1702 7866
rect 1808 7469 1814 7866
rect 1696 7457 1814 7469
rect 1930 7866 2048 7878
rect 1930 7469 1936 7866
rect 2042 7469 2048 7866
rect 1930 7457 2048 7469
rect 2164 7866 2282 7878
rect 2164 7469 2170 7866
rect 2276 7469 2282 7866
rect 2164 7457 2282 7469
rect 2398 7866 2516 7878
rect 2398 7469 2404 7866
rect 2510 7469 2516 7866
rect 2398 7457 2516 7469
rect 2632 7866 2750 7878
rect 2632 7469 2638 7866
rect 2744 7469 2750 7866
rect 2632 7457 2750 7469
rect 2866 7866 2984 7878
rect 2866 7469 2872 7866
rect 2978 7469 2984 7866
rect 2866 7457 2984 7469
rect 3100 7866 3218 7878
rect 3100 7469 3106 7866
rect 3212 7469 3218 7866
rect 3100 7457 3218 7469
rect 3334 7866 3452 7878
rect 3334 7469 3340 7866
rect 3446 7469 3452 7866
rect 3334 7457 3452 7469
rect 3568 7866 3686 7878
rect 3568 7469 3574 7866
rect 3680 7469 3686 7866
rect 3568 7457 3686 7469
rect 3802 7866 3920 7878
rect 3802 7469 3808 7866
rect 3914 7469 3920 7866
rect 3802 7457 3920 7469
rect 4036 7866 4154 7878
rect 4036 7469 4042 7866
rect 4148 7469 4154 7866
rect 4036 7457 4154 7469
rect 4270 7866 4388 7878
rect 4270 7469 4276 7866
rect 4382 7469 4388 7866
rect 4270 7457 4388 7469
rect 4504 7866 4622 7878
rect 4504 7469 4510 7866
rect 4616 7469 4622 7866
rect 4504 7457 4622 7469
rect 4738 7866 4856 7878
rect 4738 7469 4744 7866
rect 4850 7469 4856 7866
rect 4738 7457 4856 7469
rect 4972 7866 5090 7878
rect 4972 7469 4978 7866
rect 5084 7469 5090 7866
rect 4972 7457 5090 7469
rect 5206 7866 5324 7878
rect 5206 7469 5212 7866
rect 5318 7469 5324 7866
rect 5206 7457 5324 7469
rect 5440 7866 5558 7878
rect 5440 7469 5446 7866
rect 5552 7469 5558 7866
rect 5440 7457 5558 7469
rect 5674 7866 5792 7878
rect 5674 7469 5680 7866
rect 5786 7469 5792 7866
rect 5674 7457 5792 7469
rect 5908 7866 6026 7878
rect 5908 7469 5914 7866
rect 6020 7469 6026 7866
rect 5908 7457 6026 7469
rect 6142 7866 6260 7878
rect 6142 7469 6148 7866
rect 6254 7469 6260 7866
rect 6142 7457 6260 7469
rect 6376 7866 6494 7878
rect 6376 7469 6382 7866
rect 6488 7469 6494 7866
rect 6376 7457 6494 7469
rect 6610 7866 6728 7878
rect 6610 7469 6616 7866
rect 6722 7469 6728 7866
rect 6610 7457 6728 7469
rect 6844 7866 6962 7878
rect 6844 7469 6850 7866
rect 6956 7469 6962 7866
rect 6844 7457 6962 7469
rect 7078 7866 7196 7878
rect 7078 7469 7084 7866
rect 7190 7469 7196 7866
rect 7078 7457 7196 7469
rect 7312 7866 7430 7878
rect 7312 7469 7318 7866
rect 7424 7469 7430 7866
rect 7312 7457 7430 7469
rect 7546 7866 7664 7878
rect 7546 7469 7552 7866
rect 7658 7469 7664 7866
rect 7546 7457 7664 7469
rect 7780 7866 7898 7878
rect 7780 7469 7786 7866
rect 7892 7469 7898 7866
rect 7780 7457 7898 7469
rect 8014 7866 8132 7878
rect 8014 7469 8020 7866
rect 8126 7469 8132 7866
rect 8014 7457 8132 7469
rect 8248 7866 8366 7878
rect 8248 7469 8254 7866
rect 8360 7469 8366 7866
rect 8248 7457 8366 7469
rect 8482 7866 8600 7878
rect 8482 7469 8488 7866
rect 8594 7469 8600 7866
rect 8482 7457 8600 7469
rect 8716 7866 8834 7878
rect 8716 7469 8722 7866
rect 8828 7469 8834 7866
rect 8716 7457 8834 7469
rect 8950 7866 9068 7878
rect 8950 7469 8956 7866
rect 9062 7469 9068 7866
rect 8950 7457 9068 7469
rect 9184 7866 9302 7878
rect 9184 7469 9190 7866
rect 9296 7469 9302 7866
rect 9184 7457 9302 7469
rect 9418 7866 9536 7878
rect 9418 7469 9424 7866
rect 9530 7469 9536 7866
rect 9418 7457 9536 7469
rect 9652 7866 9770 7878
rect 9652 7469 9658 7866
rect 9764 7469 9770 7866
rect 9652 7457 9770 7469
rect 9886 7866 10004 7878
rect 9886 7469 9892 7866
rect 9998 7469 10004 7866
rect 9886 7457 10004 7469
rect 10120 7866 10238 7878
rect 10120 7469 10126 7866
rect 10232 7469 10238 7866
rect 10120 7457 10238 7469
rect 10354 7866 10472 7878
rect 10354 7469 10360 7866
rect 10466 7469 10472 7866
rect 10354 7457 10472 7469
rect 10588 7866 10706 7878
rect 10588 7469 10594 7866
rect 10700 7469 10706 7866
rect 10588 7457 10706 7469
rect 10822 7866 10940 7878
rect 10822 7469 10828 7866
rect 10934 7469 10940 7866
rect 10822 7457 10940 7469
rect 11056 7866 11174 7878
rect 11056 7469 11062 7866
rect 11168 7469 11174 7866
rect 11056 7457 11174 7469
rect 11290 7866 11408 7878
rect 11290 7469 11296 7866
rect 11402 7469 11408 7866
rect 11290 7457 11408 7469
rect 11524 7866 11642 7878
rect 11524 7469 11530 7866
rect 11636 7469 11642 7866
rect 11524 7457 11642 7469
rect 11758 7866 11876 7878
rect 11758 7469 11764 7866
rect 11870 7469 11876 7866
rect 11758 7457 11876 7469
rect 11992 7866 12110 7878
rect 11992 7469 11998 7866
rect 12104 7469 12110 7866
rect 11992 7457 12110 7469
rect 12226 7866 12344 7878
rect 12226 7469 12232 7866
rect 12338 7469 12344 7866
rect 12226 7457 12344 7469
rect 12460 7866 12578 7878
rect 12460 7469 12466 7866
rect 12572 7469 12578 7866
rect 12460 7457 12578 7469
rect 12694 7866 12812 7878
rect 12694 7469 12700 7866
rect 12806 7469 12812 7866
rect 12694 7457 12812 7469
rect 12928 7866 13046 7878
rect 12928 7469 12934 7866
rect 13040 7469 13046 7866
rect 12928 7457 13046 7469
rect 13162 7866 13280 7878
rect 13162 7469 13168 7866
rect 13274 7469 13280 7866
rect 13162 7457 13280 7469
rect 13396 7866 13514 7878
rect 13396 7469 13402 7866
rect 13508 7469 13514 7866
rect 13396 7457 13514 7469
rect 13630 7866 13748 7878
rect 13630 7469 13636 7866
rect 13742 7469 13748 7866
rect 13630 7457 13748 7469
rect 13864 7866 13982 7878
rect 13864 7469 13870 7866
rect 13976 7469 13982 7866
rect 13864 7457 13982 7469
rect 14098 7866 14216 7878
rect 14098 7469 14104 7866
rect 14210 7469 14216 7866
rect 14098 7457 14216 7469
rect 14332 7866 14450 7878
rect 14332 7469 14338 7866
rect 14444 7469 14450 7866
rect 14332 7457 14450 7469
rect 14566 7866 14684 7878
rect 14566 7469 14572 7866
rect 14678 7469 14684 7866
rect 14566 7457 14684 7469
rect 14800 7866 14918 7878
rect 14800 7469 14806 7866
rect 14912 7469 14918 7866
rect 14800 7457 14918 7469
rect 15034 7866 15152 7878
rect 15034 7469 15040 7866
rect 15146 7469 15152 7866
rect 15034 7457 15152 7469
rect 15268 7866 15386 7878
rect 15268 7469 15274 7866
rect 15380 7469 15386 7866
rect 15268 7457 15386 7469
rect 15502 7866 15620 7878
rect 15502 7469 15508 7866
rect 15614 7469 15620 7866
rect 15502 7457 15620 7469
rect 15736 7866 15854 7878
rect 15736 7469 15742 7866
rect 15848 7469 15854 7866
rect 15736 7457 15854 7469
rect 15970 7866 16088 7878
rect 15970 7469 15976 7866
rect 16082 7469 16088 7866
rect 15970 7457 16088 7469
rect 16204 7866 16322 7878
rect 16204 7469 16210 7866
rect 16316 7469 16322 7866
rect 16204 7457 16322 7469
rect 16438 7866 16556 7878
rect 16438 7469 16444 7866
rect 16550 7469 16556 7866
rect 16438 7457 16556 7469
rect 16672 7866 16790 7878
rect 16672 7469 16678 7866
rect 16784 7469 16790 7866
rect 16672 7457 16790 7469
rect 16906 7866 17024 7878
rect 16906 7469 16912 7866
rect 17018 7469 17024 7866
rect 16906 7457 17024 7469
rect 17140 7866 17258 7878
rect 17140 7469 17146 7866
rect 17252 7469 17258 7866
rect 17140 7457 17258 7469
rect 17374 7866 17492 7878
rect 17374 7469 17380 7866
rect 17486 7469 17492 7866
rect 17374 7457 17492 7469
rect 17608 7866 17726 7878
rect 17608 7469 17614 7866
rect 17720 7469 17726 7866
rect 17608 7457 17726 7469
rect 17842 7866 17960 7878
rect 17842 7469 17848 7866
rect 17954 7469 17960 7866
rect 17842 7457 17960 7469
rect 18076 7866 18194 7878
rect 18076 7469 18082 7866
rect 18188 7469 18194 7866
rect 18076 7457 18194 7469
rect 18310 7866 18428 7878
rect 18310 7469 18316 7866
rect 18422 7469 18428 7866
rect 18310 7457 18428 7469
rect 18544 7866 18662 7878
rect 18544 7469 18550 7866
rect 18656 7469 18662 7866
rect 18544 7457 18662 7469
rect 18778 7866 18896 7878
rect 18778 7469 18784 7866
rect 18890 7469 18896 7866
rect 18778 7457 18896 7469
rect 19012 7866 19130 7878
rect 19012 7469 19018 7866
rect 19124 7469 19130 7866
rect 19012 7457 19130 7469
rect 19246 7866 19364 7878
rect 19246 7469 19252 7866
rect 19358 7469 19364 7866
rect 19246 7457 19364 7469
rect 19480 7866 19598 7878
rect 19480 7469 19486 7866
rect 19592 7469 19598 7866
rect 19480 7457 19598 7469
rect 19714 7866 19832 7878
rect 19714 7469 19720 7866
rect 19826 7469 19832 7866
rect 19714 7457 19832 7469
rect 19948 7866 20066 7878
rect 19948 7469 19954 7866
rect 20060 7469 20066 7866
rect 19948 7457 20066 7469
rect 20182 7866 20300 7878
rect 20182 7469 20188 7866
rect 20294 7469 20300 7866
rect 20182 7457 20300 7469
rect 20416 7866 20534 7878
rect 20416 7469 20422 7866
rect 20528 7469 20534 7866
rect 20416 7457 20534 7469
rect 20650 7866 20768 7878
rect 20650 7469 20656 7866
rect 20762 7469 20768 7866
rect 20650 7457 20768 7469
rect 20884 7866 21002 7878
rect 20884 7469 20890 7866
rect 20996 7469 21002 7866
rect 20884 7457 21002 7469
rect 21118 7866 21236 7878
rect 21118 7469 21124 7866
rect 21230 7469 21236 7866
rect 21118 7457 21236 7469
rect 21352 7866 21470 7878
rect 21352 7469 21358 7866
rect 21464 7469 21470 7866
rect 21352 7457 21470 7469
rect 21586 7866 21704 7878
rect 21586 7469 21592 7866
rect 21698 7469 21704 7866
rect 21586 7457 21704 7469
rect 21820 7866 21938 7878
rect 21820 7469 21826 7866
rect 21932 7469 21938 7866
rect 21820 7457 21938 7469
rect 22054 7866 22172 7878
rect 22054 7469 22060 7866
rect 22166 7469 22172 7866
rect 22054 7457 22172 7469
rect 22288 7866 22406 7878
rect 22288 7469 22294 7866
rect 22400 7469 22406 7866
rect 22288 7457 22406 7469
rect 22522 7866 22640 7878
rect 22522 7469 22528 7866
rect 22634 7469 22640 7866
rect 22522 7457 22640 7469
rect 22756 7866 22874 7878
rect 22756 7469 22762 7866
rect 22868 7469 22874 7866
rect 22756 7457 22874 7469
rect 22990 7866 23108 7878
rect 22990 7469 22996 7866
rect 23102 7469 23108 7866
rect 22990 7457 23108 7469
rect 23224 7866 23342 7878
rect 23224 7469 23230 7866
rect 23336 7469 23342 7866
rect 23224 7457 23342 7469
rect 23458 7866 23576 7878
rect 23458 7469 23464 7866
rect 23570 7469 23576 7866
rect 23458 7457 23576 7469
rect 23692 7866 23810 7878
rect 23692 7469 23698 7866
rect 23804 7469 23810 7866
rect 23692 7457 23810 7469
rect 23926 7866 24044 7878
rect 23926 7469 23932 7866
rect 24038 7469 24044 7866
rect 23926 7457 24044 7469
rect 24160 7866 24278 7878
rect 24160 7469 24166 7866
rect 24272 7469 24278 7866
rect 24160 7457 24278 7469
rect 24394 7866 24512 7878
rect 24394 7469 24400 7866
rect 24506 7469 24512 7866
rect 24394 7457 24512 7469
rect 24628 7866 24746 7878
rect 24628 7469 24634 7866
rect 24740 7469 24746 7866
rect 24628 7457 24746 7469
rect 24862 7866 24980 7878
rect 24862 7469 24868 7866
rect 24974 7469 24980 7866
rect 24862 7457 24980 7469
rect 25096 7866 25214 7878
rect 25096 7469 25102 7866
rect 25208 7469 25214 7866
rect 25096 7457 25214 7469
rect 25330 7866 25448 7878
rect 25330 7469 25336 7866
rect 25442 7469 25448 7866
rect 25330 7457 25448 7469
rect 25564 7866 25682 7878
rect 25564 7469 25570 7866
rect 25676 7469 25682 7866
rect 25564 7457 25682 7469
rect 25798 7866 25916 7878
rect 25798 7469 25804 7866
rect 25910 7469 25916 7866
rect 25798 7457 25916 7469
rect 26032 7866 26150 7878
rect 26032 7469 26038 7866
rect 26144 7469 26150 7866
rect 26032 7457 26150 7469
rect 26266 7866 26384 7878
rect 26266 7469 26272 7866
rect 26378 7469 26384 7866
rect 26266 7457 26384 7469
rect 26500 7866 26618 7878
rect 26500 7469 26506 7866
rect 26612 7469 26618 7866
rect 26500 7457 26618 7469
rect 26734 7866 26852 7878
rect 26734 7469 26740 7866
rect 26846 7469 26852 7866
rect 26734 7457 26852 7469
rect 26968 7866 27086 7878
rect 26968 7469 26974 7866
rect 27080 7469 27086 7866
rect 26968 7457 27086 7469
rect 27202 7866 27320 7878
rect 27202 7469 27208 7866
rect 27314 7469 27320 7866
rect 27202 7457 27320 7469
rect 27436 7866 27554 7878
rect 27436 7469 27442 7866
rect 27548 7469 27554 7866
rect 27436 7457 27554 7469
rect 27670 7866 27788 7878
rect 27670 7469 27676 7866
rect 27782 7469 27788 7866
rect 27670 7457 27788 7469
rect 27904 7866 28022 7878
rect 27904 7469 27910 7866
rect 28016 7469 28022 7866
rect 27904 7457 28022 7469
rect 28138 7866 28256 7878
rect 28138 7469 28144 7866
rect 28250 7469 28256 7866
rect 28138 7457 28256 7469
rect 28372 7866 28490 7878
rect 28372 7469 28378 7866
rect 28484 7469 28490 7866
rect 28372 7457 28490 7469
rect 28606 7866 28724 7878
rect 28606 7469 28612 7866
rect 28718 7469 28724 7866
rect 28606 7457 28724 7469
rect 28840 7866 28958 7878
rect 28840 7469 28846 7866
rect 28952 7469 28958 7866
rect 28840 7457 28958 7469
rect 29074 7866 29192 7878
rect 29074 7469 29080 7866
rect 29186 7469 29192 7866
rect 29074 7457 29192 7469
rect 29308 7866 29426 7878
rect 29308 7469 29314 7866
rect 29420 7469 29426 7866
rect 29308 7457 29426 7469
rect 29542 7866 29660 7878
rect 29542 7469 29548 7866
rect 29654 7469 29660 7866
rect 29542 7457 29660 7469
rect 29776 7866 29894 7878
rect 29776 7469 29782 7866
rect 29888 7469 29894 7866
rect 29776 7457 29894 7469
rect -29894 467 -29776 479
rect -29894 70 -29888 467
rect -29782 70 -29776 467
rect -29894 58 -29776 70
rect -29660 467 -29542 479
rect -29660 70 -29654 467
rect -29548 70 -29542 467
rect -29660 58 -29542 70
rect -29426 467 -29308 479
rect -29426 70 -29420 467
rect -29314 70 -29308 467
rect -29426 58 -29308 70
rect -29192 467 -29074 479
rect -29192 70 -29186 467
rect -29080 70 -29074 467
rect -29192 58 -29074 70
rect -28958 467 -28840 479
rect -28958 70 -28952 467
rect -28846 70 -28840 467
rect -28958 58 -28840 70
rect -28724 467 -28606 479
rect -28724 70 -28718 467
rect -28612 70 -28606 467
rect -28724 58 -28606 70
rect -28490 467 -28372 479
rect -28490 70 -28484 467
rect -28378 70 -28372 467
rect -28490 58 -28372 70
rect -28256 467 -28138 479
rect -28256 70 -28250 467
rect -28144 70 -28138 467
rect -28256 58 -28138 70
rect -28022 467 -27904 479
rect -28022 70 -28016 467
rect -27910 70 -27904 467
rect -28022 58 -27904 70
rect -27788 467 -27670 479
rect -27788 70 -27782 467
rect -27676 70 -27670 467
rect -27788 58 -27670 70
rect -27554 467 -27436 479
rect -27554 70 -27548 467
rect -27442 70 -27436 467
rect -27554 58 -27436 70
rect -27320 467 -27202 479
rect -27320 70 -27314 467
rect -27208 70 -27202 467
rect -27320 58 -27202 70
rect -27086 467 -26968 479
rect -27086 70 -27080 467
rect -26974 70 -26968 467
rect -27086 58 -26968 70
rect -26852 467 -26734 479
rect -26852 70 -26846 467
rect -26740 70 -26734 467
rect -26852 58 -26734 70
rect -26618 467 -26500 479
rect -26618 70 -26612 467
rect -26506 70 -26500 467
rect -26618 58 -26500 70
rect -26384 467 -26266 479
rect -26384 70 -26378 467
rect -26272 70 -26266 467
rect -26384 58 -26266 70
rect -26150 467 -26032 479
rect -26150 70 -26144 467
rect -26038 70 -26032 467
rect -26150 58 -26032 70
rect -25916 467 -25798 479
rect -25916 70 -25910 467
rect -25804 70 -25798 467
rect -25916 58 -25798 70
rect -25682 467 -25564 479
rect -25682 70 -25676 467
rect -25570 70 -25564 467
rect -25682 58 -25564 70
rect -25448 467 -25330 479
rect -25448 70 -25442 467
rect -25336 70 -25330 467
rect -25448 58 -25330 70
rect -25214 467 -25096 479
rect -25214 70 -25208 467
rect -25102 70 -25096 467
rect -25214 58 -25096 70
rect -24980 467 -24862 479
rect -24980 70 -24974 467
rect -24868 70 -24862 467
rect -24980 58 -24862 70
rect -24746 467 -24628 479
rect -24746 70 -24740 467
rect -24634 70 -24628 467
rect -24746 58 -24628 70
rect -24512 467 -24394 479
rect -24512 70 -24506 467
rect -24400 70 -24394 467
rect -24512 58 -24394 70
rect -24278 467 -24160 479
rect -24278 70 -24272 467
rect -24166 70 -24160 467
rect -24278 58 -24160 70
rect -24044 467 -23926 479
rect -24044 70 -24038 467
rect -23932 70 -23926 467
rect -24044 58 -23926 70
rect -23810 467 -23692 479
rect -23810 70 -23804 467
rect -23698 70 -23692 467
rect -23810 58 -23692 70
rect -23576 467 -23458 479
rect -23576 70 -23570 467
rect -23464 70 -23458 467
rect -23576 58 -23458 70
rect -23342 467 -23224 479
rect -23342 70 -23336 467
rect -23230 70 -23224 467
rect -23342 58 -23224 70
rect -23108 467 -22990 479
rect -23108 70 -23102 467
rect -22996 70 -22990 467
rect -23108 58 -22990 70
rect -22874 467 -22756 479
rect -22874 70 -22868 467
rect -22762 70 -22756 467
rect -22874 58 -22756 70
rect -22640 467 -22522 479
rect -22640 70 -22634 467
rect -22528 70 -22522 467
rect -22640 58 -22522 70
rect -22406 467 -22288 479
rect -22406 70 -22400 467
rect -22294 70 -22288 467
rect -22406 58 -22288 70
rect -22172 467 -22054 479
rect -22172 70 -22166 467
rect -22060 70 -22054 467
rect -22172 58 -22054 70
rect -21938 467 -21820 479
rect -21938 70 -21932 467
rect -21826 70 -21820 467
rect -21938 58 -21820 70
rect -21704 467 -21586 479
rect -21704 70 -21698 467
rect -21592 70 -21586 467
rect -21704 58 -21586 70
rect -21470 467 -21352 479
rect -21470 70 -21464 467
rect -21358 70 -21352 467
rect -21470 58 -21352 70
rect -21236 467 -21118 479
rect -21236 70 -21230 467
rect -21124 70 -21118 467
rect -21236 58 -21118 70
rect -21002 467 -20884 479
rect -21002 70 -20996 467
rect -20890 70 -20884 467
rect -21002 58 -20884 70
rect -20768 467 -20650 479
rect -20768 70 -20762 467
rect -20656 70 -20650 467
rect -20768 58 -20650 70
rect -20534 467 -20416 479
rect -20534 70 -20528 467
rect -20422 70 -20416 467
rect -20534 58 -20416 70
rect -20300 467 -20182 479
rect -20300 70 -20294 467
rect -20188 70 -20182 467
rect -20300 58 -20182 70
rect -20066 467 -19948 479
rect -20066 70 -20060 467
rect -19954 70 -19948 467
rect -20066 58 -19948 70
rect -19832 467 -19714 479
rect -19832 70 -19826 467
rect -19720 70 -19714 467
rect -19832 58 -19714 70
rect -19598 467 -19480 479
rect -19598 70 -19592 467
rect -19486 70 -19480 467
rect -19598 58 -19480 70
rect -19364 467 -19246 479
rect -19364 70 -19358 467
rect -19252 70 -19246 467
rect -19364 58 -19246 70
rect -19130 467 -19012 479
rect -19130 70 -19124 467
rect -19018 70 -19012 467
rect -19130 58 -19012 70
rect -18896 467 -18778 479
rect -18896 70 -18890 467
rect -18784 70 -18778 467
rect -18896 58 -18778 70
rect -18662 467 -18544 479
rect -18662 70 -18656 467
rect -18550 70 -18544 467
rect -18662 58 -18544 70
rect -18428 467 -18310 479
rect -18428 70 -18422 467
rect -18316 70 -18310 467
rect -18428 58 -18310 70
rect -18194 467 -18076 479
rect -18194 70 -18188 467
rect -18082 70 -18076 467
rect -18194 58 -18076 70
rect -17960 467 -17842 479
rect -17960 70 -17954 467
rect -17848 70 -17842 467
rect -17960 58 -17842 70
rect -17726 467 -17608 479
rect -17726 70 -17720 467
rect -17614 70 -17608 467
rect -17726 58 -17608 70
rect -17492 467 -17374 479
rect -17492 70 -17486 467
rect -17380 70 -17374 467
rect -17492 58 -17374 70
rect -17258 467 -17140 479
rect -17258 70 -17252 467
rect -17146 70 -17140 467
rect -17258 58 -17140 70
rect -17024 467 -16906 479
rect -17024 70 -17018 467
rect -16912 70 -16906 467
rect -17024 58 -16906 70
rect -16790 467 -16672 479
rect -16790 70 -16784 467
rect -16678 70 -16672 467
rect -16790 58 -16672 70
rect -16556 467 -16438 479
rect -16556 70 -16550 467
rect -16444 70 -16438 467
rect -16556 58 -16438 70
rect -16322 467 -16204 479
rect -16322 70 -16316 467
rect -16210 70 -16204 467
rect -16322 58 -16204 70
rect -16088 467 -15970 479
rect -16088 70 -16082 467
rect -15976 70 -15970 467
rect -16088 58 -15970 70
rect -15854 467 -15736 479
rect -15854 70 -15848 467
rect -15742 70 -15736 467
rect -15854 58 -15736 70
rect -15620 467 -15502 479
rect -15620 70 -15614 467
rect -15508 70 -15502 467
rect -15620 58 -15502 70
rect -15386 467 -15268 479
rect -15386 70 -15380 467
rect -15274 70 -15268 467
rect -15386 58 -15268 70
rect -15152 467 -15034 479
rect -15152 70 -15146 467
rect -15040 70 -15034 467
rect -15152 58 -15034 70
rect -14918 467 -14800 479
rect -14918 70 -14912 467
rect -14806 70 -14800 467
rect -14918 58 -14800 70
rect -14684 467 -14566 479
rect -14684 70 -14678 467
rect -14572 70 -14566 467
rect -14684 58 -14566 70
rect -14450 467 -14332 479
rect -14450 70 -14444 467
rect -14338 70 -14332 467
rect -14450 58 -14332 70
rect -14216 467 -14098 479
rect -14216 70 -14210 467
rect -14104 70 -14098 467
rect -14216 58 -14098 70
rect -13982 467 -13864 479
rect -13982 70 -13976 467
rect -13870 70 -13864 467
rect -13982 58 -13864 70
rect -13748 467 -13630 479
rect -13748 70 -13742 467
rect -13636 70 -13630 467
rect -13748 58 -13630 70
rect -13514 467 -13396 479
rect -13514 70 -13508 467
rect -13402 70 -13396 467
rect -13514 58 -13396 70
rect -13280 467 -13162 479
rect -13280 70 -13274 467
rect -13168 70 -13162 467
rect -13280 58 -13162 70
rect -13046 467 -12928 479
rect -13046 70 -13040 467
rect -12934 70 -12928 467
rect -13046 58 -12928 70
rect -12812 467 -12694 479
rect -12812 70 -12806 467
rect -12700 70 -12694 467
rect -12812 58 -12694 70
rect -12578 467 -12460 479
rect -12578 70 -12572 467
rect -12466 70 -12460 467
rect -12578 58 -12460 70
rect -12344 467 -12226 479
rect -12344 70 -12338 467
rect -12232 70 -12226 467
rect -12344 58 -12226 70
rect -12110 467 -11992 479
rect -12110 70 -12104 467
rect -11998 70 -11992 467
rect -12110 58 -11992 70
rect -11876 467 -11758 479
rect -11876 70 -11870 467
rect -11764 70 -11758 467
rect -11876 58 -11758 70
rect -11642 467 -11524 479
rect -11642 70 -11636 467
rect -11530 70 -11524 467
rect -11642 58 -11524 70
rect -11408 467 -11290 479
rect -11408 70 -11402 467
rect -11296 70 -11290 467
rect -11408 58 -11290 70
rect -11174 467 -11056 479
rect -11174 70 -11168 467
rect -11062 70 -11056 467
rect -11174 58 -11056 70
rect -10940 467 -10822 479
rect -10940 70 -10934 467
rect -10828 70 -10822 467
rect -10940 58 -10822 70
rect -10706 467 -10588 479
rect -10706 70 -10700 467
rect -10594 70 -10588 467
rect -10706 58 -10588 70
rect -10472 467 -10354 479
rect -10472 70 -10466 467
rect -10360 70 -10354 467
rect -10472 58 -10354 70
rect -10238 467 -10120 479
rect -10238 70 -10232 467
rect -10126 70 -10120 467
rect -10238 58 -10120 70
rect -10004 467 -9886 479
rect -10004 70 -9998 467
rect -9892 70 -9886 467
rect -10004 58 -9886 70
rect -9770 467 -9652 479
rect -9770 70 -9764 467
rect -9658 70 -9652 467
rect -9770 58 -9652 70
rect -9536 467 -9418 479
rect -9536 70 -9530 467
rect -9424 70 -9418 467
rect -9536 58 -9418 70
rect -9302 467 -9184 479
rect -9302 70 -9296 467
rect -9190 70 -9184 467
rect -9302 58 -9184 70
rect -9068 467 -8950 479
rect -9068 70 -9062 467
rect -8956 70 -8950 467
rect -9068 58 -8950 70
rect -8834 467 -8716 479
rect -8834 70 -8828 467
rect -8722 70 -8716 467
rect -8834 58 -8716 70
rect -8600 467 -8482 479
rect -8600 70 -8594 467
rect -8488 70 -8482 467
rect -8600 58 -8482 70
rect -8366 467 -8248 479
rect -8366 70 -8360 467
rect -8254 70 -8248 467
rect -8366 58 -8248 70
rect -8132 467 -8014 479
rect -8132 70 -8126 467
rect -8020 70 -8014 467
rect -8132 58 -8014 70
rect -7898 467 -7780 479
rect -7898 70 -7892 467
rect -7786 70 -7780 467
rect -7898 58 -7780 70
rect -7664 467 -7546 479
rect -7664 70 -7658 467
rect -7552 70 -7546 467
rect -7664 58 -7546 70
rect -7430 467 -7312 479
rect -7430 70 -7424 467
rect -7318 70 -7312 467
rect -7430 58 -7312 70
rect -7196 467 -7078 479
rect -7196 70 -7190 467
rect -7084 70 -7078 467
rect -7196 58 -7078 70
rect -6962 467 -6844 479
rect -6962 70 -6956 467
rect -6850 70 -6844 467
rect -6962 58 -6844 70
rect -6728 467 -6610 479
rect -6728 70 -6722 467
rect -6616 70 -6610 467
rect -6728 58 -6610 70
rect -6494 467 -6376 479
rect -6494 70 -6488 467
rect -6382 70 -6376 467
rect -6494 58 -6376 70
rect -6260 467 -6142 479
rect -6260 70 -6254 467
rect -6148 70 -6142 467
rect -6260 58 -6142 70
rect -6026 467 -5908 479
rect -6026 70 -6020 467
rect -5914 70 -5908 467
rect -6026 58 -5908 70
rect -5792 467 -5674 479
rect -5792 70 -5786 467
rect -5680 70 -5674 467
rect -5792 58 -5674 70
rect -5558 467 -5440 479
rect -5558 70 -5552 467
rect -5446 70 -5440 467
rect -5558 58 -5440 70
rect -5324 467 -5206 479
rect -5324 70 -5318 467
rect -5212 70 -5206 467
rect -5324 58 -5206 70
rect -5090 467 -4972 479
rect -5090 70 -5084 467
rect -4978 70 -4972 467
rect -5090 58 -4972 70
rect -4856 467 -4738 479
rect -4856 70 -4850 467
rect -4744 70 -4738 467
rect -4856 58 -4738 70
rect -4622 467 -4504 479
rect -4622 70 -4616 467
rect -4510 70 -4504 467
rect -4622 58 -4504 70
rect -4388 467 -4270 479
rect -4388 70 -4382 467
rect -4276 70 -4270 467
rect -4388 58 -4270 70
rect -4154 467 -4036 479
rect -4154 70 -4148 467
rect -4042 70 -4036 467
rect -4154 58 -4036 70
rect -3920 467 -3802 479
rect -3920 70 -3914 467
rect -3808 70 -3802 467
rect -3920 58 -3802 70
rect -3686 467 -3568 479
rect -3686 70 -3680 467
rect -3574 70 -3568 467
rect -3686 58 -3568 70
rect -3452 467 -3334 479
rect -3452 70 -3446 467
rect -3340 70 -3334 467
rect -3452 58 -3334 70
rect -3218 467 -3100 479
rect -3218 70 -3212 467
rect -3106 70 -3100 467
rect -3218 58 -3100 70
rect -2984 467 -2866 479
rect -2984 70 -2978 467
rect -2872 70 -2866 467
rect -2984 58 -2866 70
rect -2750 467 -2632 479
rect -2750 70 -2744 467
rect -2638 70 -2632 467
rect -2750 58 -2632 70
rect -2516 467 -2398 479
rect -2516 70 -2510 467
rect -2404 70 -2398 467
rect -2516 58 -2398 70
rect -2282 467 -2164 479
rect -2282 70 -2276 467
rect -2170 70 -2164 467
rect -2282 58 -2164 70
rect -2048 467 -1930 479
rect -2048 70 -2042 467
rect -1936 70 -1930 467
rect -2048 58 -1930 70
rect -1814 467 -1696 479
rect -1814 70 -1808 467
rect -1702 70 -1696 467
rect -1814 58 -1696 70
rect -1580 467 -1462 479
rect -1580 70 -1574 467
rect -1468 70 -1462 467
rect -1580 58 -1462 70
rect -1346 467 -1228 479
rect -1346 70 -1340 467
rect -1234 70 -1228 467
rect -1346 58 -1228 70
rect -1112 467 -994 479
rect -1112 70 -1106 467
rect -1000 70 -994 467
rect -1112 58 -994 70
rect -878 467 -760 479
rect -878 70 -872 467
rect -766 70 -760 467
rect -878 58 -760 70
rect -644 467 -526 479
rect -644 70 -638 467
rect -532 70 -526 467
rect -644 58 -526 70
rect -410 467 -292 479
rect -410 70 -404 467
rect -298 70 -292 467
rect -410 58 -292 70
rect -176 467 -58 479
rect -176 70 -170 467
rect -64 70 -58 467
rect -176 58 -58 70
rect 58 467 176 479
rect 58 70 64 467
rect 170 70 176 467
rect 58 58 176 70
rect 292 467 410 479
rect 292 70 298 467
rect 404 70 410 467
rect 292 58 410 70
rect 526 467 644 479
rect 526 70 532 467
rect 638 70 644 467
rect 526 58 644 70
rect 760 467 878 479
rect 760 70 766 467
rect 872 70 878 467
rect 760 58 878 70
rect 994 467 1112 479
rect 994 70 1000 467
rect 1106 70 1112 467
rect 994 58 1112 70
rect 1228 467 1346 479
rect 1228 70 1234 467
rect 1340 70 1346 467
rect 1228 58 1346 70
rect 1462 467 1580 479
rect 1462 70 1468 467
rect 1574 70 1580 467
rect 1462 58 1580 70
rect 1696 467 1814 479
rect 1696 70 1702 467
rect 1808 70 1814 467
rect 1696 58 1814 70
rect 1930 467 2048 479
rect 1930 70 1936 467
rect 2042 70 2048 467
rect 1930 58 2048 70
rect 2164 467 2282 479
rect 2164 70 2170 467
rect 2276 70 2282 467
rect 2164 58 2282 70
rect 2398 467 2516 479
rect 2398 70 2404 467
rect 2510 70 2516 467
rect 2398 58 2516 70
rect 2632 467 2750 479
rect 2632 70 2638 467
rect 2744 70 2750 467
rect 2632 58 2750 70
rect 2866 467 2984 479
rect 2866 70 2872 467
rect 2978 70 2984 467
rect 2866 58 2984 70
rect 3100 467 3218 479
rect 3100 70 3106 467
rect 3212 70 3218 467
rect 3100 58 3218 70
rect 3334 467 3452 479
rect 3334 70 3340 467
rect 3446 70 3452 467
rect 3334 58 3452 70
rect 3568 467 3686 479
rect 3568 70 3574 467
rect 3680 70 3686 467
rect 3568 58 3686 70
rect 3802 467 3920 479
rect 3802 70 3808 467
rect 3914 70 3920 467
rect 3802 58 3920 70
rect 4036 467 4154 479
rect 4036 70 4042 467
rect 4148 70 4154 467
rect 4036 58 4154 70
rect 4270 467 4388 479
rect 4270 70 4276 467
rect 4382 70 4388 467
rect 4270 58 4388 70
rect 4504 467 4622 479
rect 4504 70 4510 467
rect 4616 70 4622 467
rect 4504 58 4622 70
rect 4738 467 4856 479
rect 4738 70 4744 467
rect 4850 70 4856 467
rect 4738 58 4856 70
rect 4972 467 5090 479
rect 4972 70 4978 467
rect 5084 70 5090 467
rect 4972 58 5090 70
rect 5206 467 5324 479
rect 5206 70 5212 467
rect 5318 70 5324 467
rect 5206 58 5324 70
rect 5440 467 5558 479
rect 5440 70 5446 467
rect 5552 70 5558 467
rect 5440 58 5558 70
rect 5674 467 5792 479
rect 5674 70 5680 467
rect 5786 70 5792 467
rect 5674 58 5792 70
rect 5908 467 6026 479
rect 5908 70 5914 467
rect 6020 70 6026 467
rect 5908 58 6026 70
rect 6142 467 6260 479
rect 6142 70 6148 467
rect 6254 70 6260 467
rect 6142 58 6260 70
rect 6376 467 6494 479
rect 6376 70 6382 467
rect 6488 70 6494 467
rect 6376 58 6494 70
rect 6610 467 6728 479
rect 6610 70 6616 467
rect 6722 70 6728 467
rect 6610 58 6728 70
rect 6844 467 6962 479
rect 6844 70 6850 467
rect 6956 70 6962 467
rect 6844 58 6962 70
rect 7078 467 7196 479
rect 7078 70 7084 467
rect 7190 70 7196 467
rect 7078 58 7196 70
rect 7312 467 7430 479
rect 7312 70 7318 467
rect 7424 70 7430 467
rect 7312 58 7430 70
rect 7546 467 7664 479
rect 7546 70 7552 467
rect 7658 70 7664 467
rect 7546 58 7664 70
rect 7780 467 7898 479
rect 7780 70 7786 467
rect 7892 70 7898 467
rect 7780 58 7898 70
rect 8014 467 8132 479
rect 8014 70 8020 467
rect 8126 70 8132 467
rect 8014 58 8132 70
rect 8248 467 8366 479
rect 8248 70 8254 467
rect 8360 70 8366 467
rect 8248 58 8366 70
rect 8482 467 8600 479
rect 8482 70 8488 467
rect 8594 70 8600 467
rect 8482 58 8600 70
rect 8716 467 8834 479
rect 8716 70 8722 467
rect 8828 70 8834 467
rect 8716 58 8834 70
rect 8950 467 9068 479
rect 8950 70 8956 467
rect 9062 70 9068 467
rect 8950 58 9068 70
rect 9184 467 9302 479
rect 9184 70 9190 467
rect 9296 70 9302 467
rect 9184 58 9302 70
rect 9418 467 9536 479
rect 9418 70 9424 467
rect 9530 70 9536 467
rect 9418 58 9536 70
rect 9652 467 9770 479
rect 9652 70 9658 467
rect 9764 70 9770 467
rect 9652 58 9770 70
rect 9886 467 10004 479
rect 9886 70 9892 467
rect 9998 70 10004 467
rect 9886 58 10004 70
rect 10120 467 10238 479
rect 10120 70 10126 467
rect 10232 70 10238 467
rect 10120 58 10238 70
rect 10354 467 10472 479
rect 10354 70 10360 467
rect 10466 70 10472 467
rect 10354 58 10472 70
rect 10588 467 10706 479
rect 10588 70 10594 467
rect 10700 70 10706 467
rect 10588 58 10706 70
rect 10822 467 10940 479
rect 10822 70 10828 467
rect 10934 70 10940 467
rect 10822 58 10940 70
rect 11056 467 11174 479
rect 11056 70 11062 467
rect 11168 70 11174 467
rect 11056 58 11174 70
rect 11290 467 11408 479
rect 11290 70 11296 467
rect 11402 70 11408 467
rect 11290 58 11408 70
rect 11524 467 11642 479
rect 11524 70 11530 467
rect 11636 70 11642 467
rect 11524 58 11642 70
rect 11758 467 11876 479
rect 11758 70 11764 467
rect 11870 70 11876 467
rect 11758 58 11876 70
rect 11992 467 12110 479
rect 11992 70 11998 467
rect 12104 70 12110 467
rect 11992 58 12110 70
rect 12226 467 12344 479
rect 12226 70 12232 467
rect 12338 70 12344 467
rect 12226 58 12344 70
rect 12460 467 12578 479
rect 12460 70 12466 467
rect 12572 70 12578 467
rect 12460 58 12578 70
rect 12694 467 12812 479
rect 12694 70 12700 467
rect 12806 70 12812 467
rect 12694 58 12812 70
rect 12928 467 13046 479
rect 12928 70 12934 467
rect 13040 70 13046 467
rect 12928 58 13046 70
rect 13162 467 13280 479
rect 13162 70 13168 467
rect 13274 70 13280 467
rect 13162 58 13280 70
rect 13396 467 13514 479
rect 13396 70 13402 467
rect 13508 70 13514 467
rect 13396 58 13514 70
rect 13630 467 13748 479
rect 13630 70 13636 467
rect 13742 70 13748 467
rect 13630 58 13748 70
rect 13864 467 13982 479
rect 13864 70 13870 467
rect 13976 70 13982 467
rect 13864 58 13982 70
rect 14098 467 14216 479
rect 14098 70 14104 467
rect 14210 70 14216 467
rect 14098 58 14216 70
rect 14332 467 14450 479
rect 14332 70 14338 467
rect 14444 70 14450 467
rect 14332 58 14450 70
rect 14566 467 14684 479
rect 14566 70 14572 467
rect 14678 70 14684 467
rect 14566 58 14684 70
rect 14800 467 14918 479
rect 14800 70 14806 467
rect 14912 70 14918 467
rect 14800 58 14918 70
rect 15034 467 15152 479
rect 15034 70 15040 467
rect 15146 70 15152 467
rect 15034 58 15152 70
rect 15268 467 15386 479
rect 15268 70 15274 467
rect 15380 70 15386 467
rect 15268 58 15386 70
rect 15502 467 15620 479
rect 15502 70 15508 467
rect 15614 70 15620 467
rect 15502 58 15620 70
rect 15736 467 15854 479
rect 15736 70 15742 467
rect 15848 70 15854 467
rect 15736 58 15854 70
rect 15970 467 16088 479
rect 15970 70 15976 467
rect 16082 70 16088 467
rect 15970 58 16088 70
rect 16204 467 16322 479
rect 16204 70 16210 467
rect 16316 70 16322 467
rect 16204 58 16322 70
rect 16438 467 16556 479
rect 16438 70 16444 467
rect 16550 70 16556 467
rect 16438 58 16556 70
rect 16672 467 16790 479
rect 16672 70 16678 467
rect 16784 70 16790 467
rect 16672 58 16790 70
rect 16906 467 17024 479
rect 16906 70 16912 467
rect 17018 70 17024 467
rect 16906 58 17024 70
rect 17140 467 17258 479
rect 17140 70 17146 467
rect 17252 70 17258 467
rect 17140 58 17258 70
rect 17374 467 17492 479
rect 17374 70 17380 467
rect 17486 70 17492 467
rect 17374 58 17492 70
rect 17608 467 17726 479
rect 17608 70 17614 467
rect 17720 70 17726 467
rect 17608 58 17726 70
rect 17842 467 17960 479
rect 17842 70 17848 467
rect 17954 70 17960 467
rect 17842 58 17960 70
rect 18076 467 18194 479
rect 18076 70 18082 467
rect 18188 70 18194 467
rect 18076 58 18194 70
rect 18310 467 18428 479
rect 18310 70 18316 467
rect 18422 70 18428 467
rect 18310 58 18428 70
rect 18544 467 18662 479
rect 18544 70 18550 467
rect 18656 70 18662 467
rect 18544 58 18662 70
rect 18778 467 18896 479
rect 18778 70 18784 467
rect 18890 70 18896 467
rect 18778 58 18896 70
rect 19012 467 19130 479
rect 19012 70 19018 467
rect 19124 70 19130 467
rect 19012 58 19130 70
rect 19246 467 19364 479
rect 19246 70 19252 467
rect 19358 70 19364 467
rect 19246 58 19364 70
rect 19480 467 19598 479
rect 19480 70 19486 467
rect 19592 70 19598 467
rect 19480 58 19598 70
rect 19714 467 19832 479
rect 19714 70 19720 467
rect 19826 70 19832 467
rect 19714 58 19832 70
rect 19948 467 20066 479
rect 19948 70 19954 467
rect 20060 70 20066 467
rect 19948 58 20066 70
rect 20182 467 20300 479
rect 20182 70 20188 467
rect 20294 70 20300 467
rect 20182 58 20300 70
rect 20416 467 20534 479
rect 20416 70 20422 467
rect 20528 70 20534 467
rect 20416 58 20534 70
rect 20650 467 20768 479
rect 20650 70 20656 467
rect 20762 70 20768 467
rect 20650 58 20768 70
rect 20884 467 21002 479
rect 20884 70 20890 467
rect 20996 70 21002 467
rect 20884 58 21002 70
rect 21118 467 21236 479
rect 21118 70 21124 467
rect 21230 70 21236 467
rect 21118 58 21236 70
rect 21352 467 21470 479
rect 21352 70 21358 467
rect 21464 70 21470 467
rect 21352 58 21470 70
rect 21586 467 21704 479
rect 21586 70 21592 467
rect 21698 70 21704 467
rect 21586 58 21704 70
rect 21820 467 21938 479
rect 21820 70 21826 467
rect 21932 70 21938 467
rect 21820 58 21938 70
rect 22054 467 22172 479
rect 22054 70 22060 467
rect 22166 70 22172 467
rect 22054 58 22172 70
rect 22288 467 22406 479
rect 22288 70 22294 467
rect 22400 70 22406 467
rect 22288 58 22406 70
rect 22522 467 22640 479
rect 22522 70 22528 467
rect 22634 70 22640 467
rect 22522 58 22640 70
rect 22756 467 22874 479
rect 22756 70 22762 467
rect 22868 70 22874 467
rect 22756 58 22874 70
rect 22990 467 23108 479
rect 22990 70 22996 467
rect 23102 70 23108 467
rect 22990 58 23108 70
rect 23224 467 23342 479
rect 23224 70 23230 467
rect 23336 70 23342 467
rect 23224 58 23342 70
rect 23458 467 23576 479
rect 23458 70 23464 467
rect 23570 70 23576 467
rect 23458 58 23576 70
rect 23692 467 23810 479
rect 23692 70 23698 467
rect 23804 70 23810 467
rect 23692 58 23810 70
rect 23926 467 24044 479
rect 23926 70 23932 467
rect 24038 70 24044 467
rect 23926 58 24044 70
rect 24160 467 24278 479
rect 24160 70 24166 467
rect 24272 70 24278 467
rect 24160 58 24278 70
rect 24394 467 24512 479
rect 24394 70 24400 467
rect 24506 70 24512 467
rect 24394 58 24512 70
rect 24628 467 24746 479
rect 24628 70 24634 467
rect 24740 70 24746 467
rect 24628 58 24746 70
rect 24862 467 24980 479
rect 24862 70 24868 467
rect 24974 70 24980 467
rect 24862 58 24980 70
rect 25096 467 25214 479
rect 25096 70 25102 467
rect 25208 70 25214 467
rect 25096 58 25214 70
rect 25330 467 25448 479
rect 25330 70 25336 467
rect 25442 70 25448 467
rect 25330 58 25448 70
rect 25564 467 25682 479
rect 25564 70 25570 467
rect 25676 70 25682 467
rect 25564 58 25682 70
rect 25798 467 25916 479
rect 25798 70 25804 467
rect 25910 70 25916 467
rect 25798 58 25916 70
rect 26032 467 26150 479
rect 26032 70 26038 467
rect 26144 70 26150 467
rect 26032 58 26150 70
rect 26266 467 26384 479
rect 26266 70 26272 467
rect 26378 70 26384 467
rect 26266 58 26384 70
rect 26500 467 26618 479
rect 26500 70 26506 467
rect 26612 70 26618 467
rect 26500 58 26618 70
rect 26734 467 26852 479
rect 26734 70 26740 467
rect 26846 70 26852 467
rect 26734 58 26852 70
rect 26968 467 27086 479
rect 26968 70 26974 467
rect 27080 70 27086 467
rect 26968 58 27086 70
rect 27202 467 27320 479
rect 27202 70 27208 467
rect 27314 70 27320 467
rect 27202 58 27320 70
rect 27436 467 27554 479
rect 27436 70 27442 467
rect 27548 70 27554 467
rect 27436 58 27554 70
rect 27670 467 27788 479
rect 27670 70 27676 467
rect 27782 70 27788 467
rect 27670 58 27788 70
rect 27904 467 28022 479
rect 27904 70 27910 467
rect 28016 70 28022 467
rect 27904 58 28022 70
rect 28138 467 28256 479
rect 28138 70 28144 467
rect 28250 70 28256 467
rect 28138 58 28256 70
rect 28372 467 28490 479
rect 28372 70 28378 467
rect 28484 70 28490 467
rect 28372 58 28490 70
rect 28606 467 28724 479
rect 28606 70 28612 467
rect 28718 70 28724 467
rect 28606 58 28724 70
rect 28840 467 28958 479
rect 28840 70 28846 467
rect 28952 70 28958 467
rect 28840 58 28958 70
rect 29074 467 29192 479
rect 29074 70 29080 467
rect 29186 70 29192 467
rect 29074 58 29192 70
rect 29308 467 29426 479
rect 29308 70 29314 467
rect 29420 70 29426 467
rect 29308 58 29426 70
rect 29542 467 29660 479
rect 29542 70 29548 467
rect 29654 70 29660 467
rect 29542 58 29660 70
rect 29776 467 29894 479
rect 29776 70 29782 467
rect 29888 70 29894 467
rect 29776 58 29894 70
rect -29894 -70 -29776 -58
rect -29894 -467 -29888 -70
rect -29782 -467 -29776 -70
rect -29894 -479 -29776 -467
rect -29660 -70 -29542 -58
rect -29660 -467 -29654 -70
rect -29548 -467 -29542 -70
rect -29660 -479 -29542 -467
rect -29426 -70 -29308 -58
rect -29426 -467 -29420 -70
rect -29314 -467 -29308 -70
rect -29426 -479 -29308 -467
rect -29192 -70 -29074 -58
rect -29192 -467 -29186 -70
rect -29080 -467 -29074 -70
rect -29192 -479 -29074 -467
rect -28958 -70 -28840 -58
rect -28958 -467 -28952 -70
rect -28846 -467 -28840 -70
rect -28958 -479 -28840 -467
rect -28724 -70 -28606 -58
rect -28724 -467 -28718 -70
rect -28612 -467 -28606 -70
rect -28724 -479 -28606 -467
rect -28490 -70 -28372 -58
rect -28490 -467 -28484 -70
rect -28378 -467 -28372 -70
rect -28490 -479 -28372 -467
rect -28256 -70 -28138 -58
rect -28256 -467 -28250 -70
rect -28144 -467 -28138 -70
rect -28256 -479 -28138 -467
rect -28022 -70 -27904 -58
rect -28022 -467 -28016 -70
rect -27910 -467 -27904 -70
rect -28022 -479 -27904 -467
rect -27788 -70 -27670 -58
rect -27788 -467 -27782 -70
rect -27676 -467 -27670 -70
rect -27788 -479 -27670 -467
rect -27554 -70 -27436 -58
rect -27554 -467 -27548 -70
rect -27442 -467 -27436 -70
rect -27554 -479 -27436 -467
rect -27320 -70 -27202 -58
rect -27320 -467 -27314 -70
rect -27208 -467 -27202 -70
rect -27320 -479 -27202 -467
rect -27086 -70 -26968 -58
rect -27086 -467 -27080 -70
rect -26974 -467 -26968 -70
rect -27086 -479 -26968 -467
rect -26852 -70 -26734 -58
rect -26852 -467 -26846 -70
rect -26740 -467 -26734 -70
rect -26852 -479 -26734 -467
rect -26618 -70 -26500 -58
rect -26618 -467 -26612 -70
rect -26506 -467 -26500 -70
rect -26618 -479 -26500 -467
rect -26384 -70 -26266 -58
rect -26384 -467 -26378 -70
rect -26272 -467 -26266 -70
rect -26384 -479 -26266 -467
rect -26150 -70 -26032 -58
rect -26150 -467 -26144 -70
rect -26038 -467 -26032 -70
rect -26150 -479 -26032 -467
rect -25916 -70 -25798 -58
rect -25916 -467 -25910 -70
rect -25804 -467 -25798 -70
rect -25916 -479 -25798 -467
rect -25682 -70 -25564 -58
rect -25682 -467 -25676 -70
rect -25570 -467 -25564 -70
rect -25682 -479 -25564 -467
rect -25448 -70 -25330 -58
rect -25448 -467 -25442 -70
rect -25336 -467 -25330 -70
rect -25448 -479 -25330 -467
rect -25214 -70 -25096 -58
rect -25214 -467 -25208 -70
rect -25102 -467 -25096 -70
rect -25214 -479 -25096 -467
rect -24980 -70 -24862 -58
rect -24980 -467 -24974 -70
rect -24868 -467 -24862 -70
rect -24980 -479 -24862 -467
rect -24746 -70 -24628 -58
rect -24746 -467 -24740 -70
rect -24634 -467 -24628 -70
rect -24746 -479 -24628 -467
rect -24512 -70 -24394 -58
rect -24512 -467 -24506 -70
rect -24400 -467 -24394 -70
rect -24512 -479 -24394 -467
rect -24278 -70 -24160 -58
rect -24278 -467 -24272 -70
rect -24166 -467 -24160 -70
rect -24278 -479 -24160 -467
rect -24044 -70 -23926 -58
rect -24044 -467 -24038 -70
rect -23932 -467 -23926 -70
rect -24044 -479 -23926 -467
rect -23810 -70 -23692 -58
rect -23810 -467 -23804 -70
rect -23698 -467 -23692 -70
rect -23810 -479 -23692 -467
rect -23576 -70 -23458 -58
rect -23576 -467 -23570 -70
rect -23464 -467 -23458 -70
rect -23576 -479 -23458 -467
rect -23342 -70 -23224 -58
rect -23342 -467 -23336 -70
rect -23230 -467 -23224 -70
rect -23342 -479 -23224 -467
rect -23108 -70 -22990 -58
rect -23108 -467 -23102 -70
rect -22996 -467 -22990 -70
rect -23108 -479 -22990 -467
rect -22874 -70 -22756 -58
rect -22874 -467 -22868 -70
rect -22762 -467 -22756 -70
rect -22874 -479 -22756 -467
rect -22640 -70 -22522 -58
rect -22640 -467 -22634 -70
rect -22528 -467 -22522 -70
rect -22640 -479 -22522 -467
rect -22406 -70 -22288 -58
rect -22406 -467 -22400 -70
rect -22294 -467 -22288 -70
rect -22406 -479 -22288 -467
rect -22172 -70 -22054 -58
rect -22172 -467 -22166 -70
rect -22060 -467 -22054 -70
rect -22172 -479 -22054 -467
rect -21938 -70 -21820 -58
rect -21938 -467 -21932 -70
rect -21826 -467 -21820 -70
rect -21938 -479 -21820 -467
rect -21704 -70 -21586 -58
rect -21704 -467 -21698 -70
rect -21592 -467 -21586 -70
rect -21704 -479 -21586 -467
rect -21470 -70 -21352 -58
rect -21470 -467 -21464 -70
rect -21358 -467 -21352 -70
rect -21470 -479 -21352 -467
rect -21236 -70 -21118 -58
rect -21236 -467 -21230 -70
rect -21124 -467 -21118 -70
rect -21236 -479 -21118 -467
rect -21002 -70 -20884 -58
rect -21002 -467 -20996 -70
rect -20890 -467 -20884 -70
rect -21002 -479 -20884 -467
rect -20768 -70 -20650 -58
rect -20768 -467 -20762 -70
rect -20656 -467 -20650 -70
rect -20768 -479 -20650 -467
rect -20534 -70 -20416 -58
rect -20534 -467 -20528 -70
rect -20422 -467 -20416 -70
rect -20534 -479 -20416 -467
rect -20300 -70 -20182 -58
rect -20300 -467 -20294 -70
rect -20188 -467 -20182 -70
rect -20300 -479 -20182 -467
rect -20066 -70 -19948 -58
rect -20066 -467 -20060 -70
rect -19954 -467 -19948 -70
rect -20066 -479 -19948 -467
rect -19832 -70 -19714 -58
rect -19832 -467 -19826 -70
rect -19720 -467 -19714 -70
rect -19832 -479 -19714 -467
rect -19598 -70 -19480 -58
rect -19598 -467 -19592 -70
rect -19486 -467 -19480 -70
rect -19598 -479 -19480 -467
rect -19364 -70 -19246 -58
rect -19364 -467 -19358 -70
rect -19252 -467 -19246 -70
rect -19364 -479 -19246 -467
rect -19130 -70 -19012 -58
rect -19130 -467 -19124 -70
rect -19018 -467 -19012 -70
rect -19130 -479 -19012 -467
rect -18896 -70 -18778 -58
rect -18896 -467 -18890 -70
rect -18784 -467 -18778 -70
rect -18896 -479 -18778 -467
rect -18662 -70 -18544 -58
rect -18662 -467 -18656 -70
rect -18550 -467 -18544 -70
rect -18662 -479 -18544 -467
rect -18428 -70 -18310 -58
rect -18428 -467 -18422 -70
rect -18316 -467 -18310 -70
rect -18428 -479 -18310 -467
rect -18194 -70 -18076 -58
rect -18194 -467 -18188 -70
rect -18082 -467 -18076 -70
rect -18194 -479 -18076 -467
rect -17960 -70 -17842 -58
rect -17960 -467 -17954 -70
rect -17848 -467 -17842 -70
rect -17960 -479 -17842 -467
rect -17726 -70 -17608 -58
rect -17726 -467 -17720 -70
rect -17614 -467 -17608 -70
rect -17726 -479 -17608 -467
rect -17492 -70 -17374 -58
rect -17492 -467 -17486 -70
rect -17380 -467 -17374 -70
rect -17492 -479 -17374 -467
rect -17258 -70 -17140 -58
rect -17258 -467 -17252 -70
rect -17146 -467 -17140 -70
rect -17258 -479 -17140 -467
rect -17024 -70 -16906 -58
rect -17024 -467 -17018 -70
rect -16912 -467 -16906 -70
rect -17024 -479 -16906 -467
rect -16790 -70 -16672 -58
rect -16790 -467 -16784 -70
rect -16678 -467 -16672 -70
rect -16790 -479 -16672 -467
rect -16556 -70 -16438 -58
rect -16556 -467 -16550 -70
rect -16444 -467 -16438 -70
rect -16556 -479 -16438 -467
rect -16322 -70 -16204 -58
rect -16322 -467 -16316 -70
rect -16210 -467 -16204 -70
rect -16322 -479 -16204 -467
rect -16088 -70 -15970 -58
rect -16088 -467 -16082 -70
rect -15976 -467 -15970 -70
rect -16088 -479 -15970 -467
rect -15854 -70 -15736 -58
rect -15854 -467 -15848 -70
rect -15742 -467 -15736 -70
rect -15854 -479 -15736 -467
rect -15620 -70 -15502 -58
rect -15620 -467 -15614 -70
rect -15508 -467 -15502 -70
rect -15620 -479 -15502 -467
rect -15386 -70 -15268 -58
rect -15386 -467 -15380 -70
rect -15274 -467 -15268 -70
rect -15386 -479 -15268 -467
rect -15152 -70 -15034 -58
rect -15152 -467 -15146 -70
rect -15040 -467 -15034 -70
rect -15152 -479 -15034 -467
rect -14918 -70 -14800 -58
rect -14918 -467 -14912 -70
rect -14806 -467 -14800 -70
rect -14918 -479 -14800 -467
rect -14684 -70 -14566 -58
rect -14684 -467 -14678 -70
rect -14572 -467 -14566 -70
rect -14684 -479 -14566 -467
rect -14450 -70 -14332 -58
rect -14450 -467 -14444 -70
rect -14338 -467 -14332 -70
rect -14450 -479 -14332 -467
rect -14216 -70 -14098 -58
rect -14216 -467 -14210 -70
rect -14104 -467 -14098 -70
rect -14216 -479 -14098 -467
rect -13982 -70 -13864 -58
rect -13982 -467 -13976 -70
rect -13870 -467 -13864 -70
rect -13982 -479 -13864 -467
rect -13748 -70 -13630 -58
rect -13748 -467 -13742 -70
rect -13636 -467 -13630 -70
rect -13748 -479 -13630 -467
rect -13514 -70 -13396 -58
rect -13514 -467 -13508 -70
rect -13402 -467 -13396 -70
rect -13514 -479 -13396 -467
rect -13280 -70 -13162 -58
rect -13280 -467 -13274 -70
rect -13168 -467 -13162 -70
rect -13280 -479 -13162 -467
rect -13046 -70 -12928 -58
rect -13046 -467 -13040 -70
rect -12934 -467 -12928 -70
rect -13046 -479 -12928 -467
rect -12812 -70 -12694 -58
rect -12812 -467 -12806 -70
rect -12700 -467 -12694 -70
rect -12812 -479 -12694 -467
rect -12578 -70 -12460 -58
rect -12578 -467 -12572 -70
rect -12466 -467 -12460 -70
rect -12578 -479 -12460 -467
rect -12344 -70 -12226 -58
rect -12344 -467 -12338 -70
rect -12232 -467 -12226 -70
rect -12344 -479 -12226 -467
rect -12110 -70 -11992 -58
rect -12110 -467 -12104 -70
rect -11998 -467 -11992 -70
rect -12110 -479 -11992 -467
rect -11876 -70 -11758 -58
rect -11876 -467 -11870 -70
rect -11764 -467 -11758 -70
rect -11876 -479 -11758 -467
rect -11642 -70 -11524 -58
rect -11642 -467 -11636 -70
rect -11530 -467 -11524 -70
rect -11642 -479 -11524 -467
rect -11408 -70 -11290 -58
rect -11408 -467 -11402 -70
rect -11296 -467 -11290 -70
rect -11408 -479 -11290 -467
rect -11174 -70 -11056 -58
rect -11174 -467 -11168 -70
rect -11062 -467 -11056 -70
rect -11174 -479 -11056 -467
rect -10940 -70 -10822 -58
rect -10940 -467 -10934 -70
rect -10828 -467 -10822 -70
rect -10940 -479 -10822 -467
rect -10706 -70 -10588 -58
rect -10706 -467 -10700 -70
rect -10594 -467 -10588 -70
rect -10706 -479 -10588 -467
rect -10472 -70 -10354 -58
rect -10472 -467 -10466 -70
rect -10360 -467 -10354 -70
rect -10472 -479 -10354 -467
rect -10238 -70 -10120 -58
rect -10238 -467 -10232 -70
rect -10126 -467 -10120 -70
rect -10238 -479 -10120 -467
rect -10004 -70 -9886 -58
rect -10004 -467 -9998 -70
rect -9892 -467 -9886 -70
rect -10004 -479 -9886 -467
rect -9770 -70 -9652 -58
rect -9770 -467 -9764 -70
rect -9658 -467 -9652 -70
rect -9770 -479 -9652 -467
rect -9536 -70 -9418 -58
rect -9536 -467 -9530 -70
rect -9424 -467 -9418 -70
rect -9536 -479 -9418 -467
rect -9302 -70 -9184 -58
rect -9302 -467 -9296 -70
rect -9190 -467 -9184 -70
rect -9302 -479 -9184 -467
rect -9068 -70 -8950 -58
rect -9068 -467 -9062 -70
rect -8956 -467 -8950 -70
rect -9068 -479 -8950 -467
rect -8834 -70 -8716 -58
rect -8834 -467 -8828 -70
rect -8722 -467 -8716 -70
rect -8834 -479 -8716 -467
rect -8600 -70 -8482 -58
rect -8600 -467 -8594 -70
rect -8488 -467 -8482 -70
rect -8600 -479 -8482 -467
rect -8366 -70 -8248 -58
rect -8366 -467 -8360 -70
rect -8254 -467 -8248 -70
rect -8366 -479 -8248 -467
rect -8132 -70 -8014 -58
rect -8132 -467 -8126 -70
rect -8020 -467 -8014 -70
rect -8132 -479 -8014 -467
rect -7898 -70 -7780 -58
rect -7898 -467 -7892 -70
rect -7786 -467 -7780 -70
rect -7898 -479 -7780 -467
rect -7664 -70 -7546 -58
rect -7664 -467 -7658 -70
rect -7552 -467 -7546 -70
rect -7664 -479 -7546 -467
rect -7430 -70 -7312 -58
rect -7430 -467 -7424 -70
rect -7318 -467 -7312 -70
rect -7430 -479 -7312 -467
rect -7196 -70 -7078 -58
rect -7196 -467 -7190 -70
rect -7084 -467 -7078 -70
rect -7196 -479 -7078 -467
rect -6962 -70 -6844 -58
rect -6962 -467 -6956 -70
rect -6850 -467 -6844 -70
rect -6962 -479 -6844 -467
rect -6728 -70 -6610 -58
rect -6728 -467 -6722 -70
rect -6616 -467 -6610 -70
rect -6728 -479 -6610 -467
rect -6494 -70 -6376 -58
rect -6494 -467 -6488 -70
rect -6382 -467 -6376 -70
rect -6494 -479 -6376 -467
rect -6260 -70 -6142 -58
rect -6260 -467 -6254 -70
rect -6148 -467 -6142 -70
rect -6260 -479 -6142 -467
rect -6026 -70 -5908 -58
rect -6026 -467 -6020 -70
rect -5914 -467 -5908 -70
rect -6026 -479 -5908 -467
rect -5792 -70 -5674 -58
rect -5792 -467 -5786 -70
rect -5680 -467 -5674 -70
rect -5792 -479 -5674 -467
rect -5558 -70 -5440 -58
rect -5558 -467 -5552 -70
rect -5446 -467 -5440 -70
rect -5558 -479 -5440 -467
rect -5324 -70 -5206 -58
rect -5324 -467 -5318 -70
rect -5212 -467 -5206 -70
rect -5324 -479 -5206 -467
rect -5090 -70 -4972 -58
rect -5090 -467 -5084 -70
rect -4978 -467 -4972 -70
rect -5090 -479 -4972 -467
rect -4856 -70 -4738 -58
rect -4856 -467 -4850 -70
rect -4744 -467 -4738 -70
rect -4856 -479 -4738 -467
rect -4622 -70 -4504 -58
rect -4622 -467 -4616 -70
rect -4510 -467 -4504 -70
rect -4622 -479 -4504 -467
rect -4388 -70 -4270 -58
rect -4388 -467 -4382 -70
rect -4276 -467 -4270 -70
rect -4388 -479 -4270 -467
rect -4154 -70 -4036 -58
rect -4154 -467 -4148 -70
rect -4042 -467 -4036 -70
rect -4154 -479 -4036 -467
rect -3920 -70 -3802 -58
rect -3920 -467 -3914 -70
rect -3808 -467 -3802 -70
rect -3920 -479 -3802 -467
rect -3686 -70 -3568 -58
rect -3686 -467 -3680 -70
rect -3574 -467 -3568 -70
rect -3686 -479 -3568 -467
rect -3452 -70 -3334 -58
rect -3452 -467 -3446 -70
rect -3340 -467 -3334 -70
rect -3452 -479 -3334 -467
rect -3218 -70 -3100 -58
rect -3218 -467 -3212 -70
rect -3106 -467 -3100 -70
rect -3218 -479 -3100 -467
rect -2984 -70 -2866 -58
rect -2984 -467 -2978 -70
rect -2872 -467 -2866 -70
rect -2984 -479 -2866 -467
rect -2750 -70 -2632 -58
rect -2750 -467 -2744 -70
rect -2638 -467 -2632 -70
rect -2750 -479 -2632 -467
rect -2516 -70 -2398 -58
rect -2516 -467 -2510 -70
rect -2404 -467 -2398 -70
rect -2516 -479 -2398 -467
rect -2282 -70 -2164 -58
rect -2282 -467 -2276 -70
rect -2170 -467 -2164 -70
rect -2282 -479 -2164 -467
rect -2048 -70 -1930 -58
rect -2048 -467 -2042 -70
rect -1936 -467 -1930 -70
rect -2048 -479 -1930 -467
rect -1814 -70 -1696 -58
rect -1814 -467 -1808 -70
rect -1702 -467 -1696 -70
rect -1814 -479 -1696 -467
rect -1580 -70 -1462 -58
rect -1580 -467 -1574 -70
rect -1468 -467 -1462 -70
rect -1580 -479 -1462 -467
rect -1346 -70 -1228 -58
rect -1346 -467 -1340 -70
rect -1234 -467 -1228 -70
rect -1346 -479 -1228 -467
rect -1112 -70 -994 -58
rect -1112 -467 -1106 -70
rect -1000 -467 -994 -70
rect -1112 -479 -994 -467
rect -878 -70 -760 -58
rect -878 -467 -872 -70
rect -766 -467 -760 -70
rect -878 -479 -760 -467
rect -644 -70 -526 -58
rect -644 -467 -638 -70
rect -532 -467 -526 -70
rect -644 -479 -526 -467
rect -410 -70 -292 -58
rect -410 -467 -404 -70
rect -298 -467 -292 -70
rect -410 -479 -292 -467
rect -176 -70 -58 -58
rect -176 -467 -170 -70
rect -64 -467 -58 -70
rect -176 -479 -58 -467
rect 58 -70 176 -58
rect 58 -467 64 -70
rect 170 -467 176 -70
rect 58 -479 176 -467
rect 292 -70 410 -58
rect 292 -467 298 -70
rect 404 -467 410 -70
rect 292 -479 410 -467
rect 526 -70 644 -58
rect 526 -467 532 -70
rect 638 -467 644 -70
rect 526 -479 644 -467
rect 760 -70 878 -58
rect 760 -467 766 -70
rect 872 -467 878 -70
rect 760 -479 878 -467
rect 994 -70 1112 -58
rect 994 -467 1000 -70
rect 1106 -467 1112 -70
rect 994 -479 1112 -467
rect 1228 -70 1346 -58
rect 1228 -467 1234 -70
rect 1340 -467 1346 -70
rect 1228 -479 1346 -467
rect 1462 -70 1580 -58
rect 1462 -467 1468 -70
rect 1574 -467 1580 -70
rect 1462 -479 1580 -467
rect 1696 -70 1814 -58
rect 1696 -467 1702 -70
rect 1808 -467 1814 -70
rect 1696 -479 1814 -467
rect 1930 -70 2048 -58
rect 1930 -467 1936 -70
rect 2042 -467 2048 -70
rect 1930 -479 2048 -467
rect 2164 -70 2282 -58
rect 2164 -467 2170 -70
rect 2276 -467 2282 -70
rect 2164 -479 2282 -467
rect 2398 -70 2516 -58
rect 2398 -467 2404 -70
rect 2510 -467 2516 -70
rect 2398 -479 2516 -467
rect 2632 -70 2750 -58
rect 2632 -467 2638 -70
rect 2744 -467 2750 -70
rect 2632 -479 2750 -467
rect 2866 -70 2984 -58
rect 2866 -467 2872 -70
rect 2978 -467 2984 -70
rect 2866 -479 2984 -467
rect 3100 -70 3218 -58
rect 3100 -467 3106 -70
rect 3212 -467 3218 -70
rect 3100 -479 3218 -467
rect 3334 -70 3452 -58
rect 3334 -467 3340 -70
rect 3446 -467 3452 -70
rect 3334 -479 3452 -467
rect 3568 -70 3686 -58
rect 3568 -467 3574 -70
rect 3680 -467 3686 -70
rect 3568 -479 3686 -467
rect 3802 -70 3920 -58
rect 3802 -467 3808 -70
rect 3914 -467 3920 -70
rect 3802 -479 3920 -467
rect 4036 -70 4154 -58
rect 4036 -467 4042 -70
rect 4148 -467 4154 -70
rect 4036 -479 4154 -467
rect 4270 -70 4388 -58
rect 4270 -467 4276 -70
rect 4382 -467 4388 -70
rect 4270 -479 4388 -467
rect 4504 -70 4622 -58
rect 4504 -467 4510 -70
rect 4616 -467 4622 -70
rect 4504 -479 4622 -467
rect 4738 -70 4856 -58
rect 4738 -467 4744 -70
rect 4850 -467 4856 -70
rect 4738 -479 4856 -467
rect 4972 -70 5090 -58
rect 4972 -467 4978 -70
rect 5084 -467 5090 -70
rect 4972 -479 5090 -467
rect 5206 -70 5324 -58
rect 5206 -467 5212 -70
rect 5318 -467 5324 -70
rect 5206 -479 5324 -467
rect 5440 -70 5558 -58
rect 5440 -467 5446 -70
rect 5552 -467 5558 -70
rect 5440 -479 5558 -467
rect 5674 -70 5792 -58
rect 5674 -467 5680 -70
rect 5786 -467 5792 -70
rect 5674 -479 5792 -467
rect 5908 -70 6026 -58
rect 5908 -467 5914 -70
rect 6020 -467 6026 -70
rect 5908 -479 6026 -467
rect 6142 -70 6260 -58
rect 6142 -467 6148 -70
rect 6254 -467 6260 -70
rect 6142 -479 6260 -467
rect 6376 -70 6494 -58
rect 6376 -467 6382 -70
rect 6488 -467 6494 -70
rect 6376 -479 6494 -467
rect 6610 -70 6728 -58
rect 6610 -467 6616 -70
rect 6722 -467 6728 -70
rect 6610 -479 6728 -467
rect 6844 -70 6962 -58
rect 6844 -467 6850 -70
rect 6956 -467 6962 -70
rect 6844 -479 6962 -467
rect 7078 -70 7196 -58
rect 7078 -467 7084 -70
rect 7190 -467 7196 -70
rect 7078 -479 7196 -467
rect 7312 -70 7430 -58
rect 7312 -467 7318 -70
rect 7424 -467 7430 -70
rect 7312 -479 7430 -467
rect 7546 -70 7664 -58
rect 7546 -467 7552 -70
rect 7658 -467 7664 -70
rect 7546 -479 7664 -467
rect 7780 -70 7898 -58
rect 7780 -467 7786 -70
rect 7892 -467 7898 -70
rect 7780 -479 7898 -467
rect 8014 -70 8132 -58
rect 8014 -467 8020 -70
rect 8126 -467 8132 -70
rect 8014 -479 8132 -467
rect 8248 -70 8366 -58
rect 8248 -467 8254 -70
rect 8360 -467 8366 -70
rect 8248 -479 8366 -467
rect 8482 -70 8600 -58
rect 8482 -467 8488 -70
rect 8594 -467 8600 -70
rect 8482 -479 8600 -467
rect 8716 -70 8834 -58
rect 8716 -467 8722 -70
rect 8828 -467 8834 -70
rect 8716 -479 8834 -467
rect 8950 -70 9068 -58
rect 8950 -467 8956 -70
rect 9062 -467 9068 -70
rect 8950 -479 9068 -467
rect 9184 -70 9302 -58
rect 9184 -467 9190 -70
rect 9296 -467 9302 -70
rect 9184 -479 9302 -467
rect 9418 -70 9536 -58
rect 9418 -467 9424 -70
rect 9530 -467 9536 -70
rect 9418 -479 9536 -467
rect 9652 -70 9770 -58
rect 9652 -467 9658 -70
rect 9764 -467 9770 -70
rect 9652 -479 9770 -467
rect 9886 -70 10004 -58
rect 9886 -467 9892 -70
rect 9998 -467 10004 -70
rect 9886 -479 10004 -467
rect 10120 -70 10238 -58
rect 10120 -467 10126 -70
rect 10232 -467 10238 -70
rect 10120 -479 10238 -467
rect 10354 -70 10472 -58
rect 10354 -467 10360 -70
rect 10466 -467 10472 -70
rect 10354 -479 10472 -467
rect 10588 -70 10706 -58
rect 10588 -467 10594 -70
rect 10700 -467 10706 -70
rect 10588 -479 10706 -467
rect 10822 -70 10940 -58
rect 10822 -467 10828 -70
rect 10934 -467 10940 -70
rect 10822 -479 10940 -467
rect 11056 -70 11174 -58
rect 11056 -467 11062 -70
rect 11168 -467 11174 -70
rect 11056 -479 11174 -467
rect 11290 -70 11408 -58
rect 11290 -467 11296 -70
rect 11402 -467 11408 -70
rect 11290 -479 11408 -467
rect 11524 -70 11642 -58
rect 11524 -467 11530 -70
rect 11636 -467 11642 -70
rect 11524 -479 11642 -467
rect 11758 -70 11876 -58
rect 11758 -467 11764 -70
rect 11870 -467 11876 -70
rect 11758 -479 11876 -467
rect 11992 -70 12110 -58
rect 11992 -467 11998 -70
rect 12104 -467 12110 -70
rect 11992 -479 12110 -467
rect 12226 -70 12344 -58
rect 12226 -467 12232 -70
rect 12338 -467 12344 -70
rect 12226 -479 12344 -467
rect 12460 -70 12578 -58
rect 12460 -467 12466 -70
rect 12572 -467 12578 -70
rect 12460 -479 12578 -467
rect 12694 -70 12812 -58
rect 12694 -467 12700 -70
rect 12806 -467 12812 -70
rect 12694 -479 12812 -467
rect 12928 -70 13046 -58
rect 12928 -467 12934 -70
rect 13040 -467 13046 -70
rect 12928 -479 13046 -467
rect 13162 -70 13280 -58
rect 13162 -467 13168 -70
rect 13274 -467 13280 -70
rect 13162 -479 13280 -467
rect 13396 -70 13514 -58
rect 13396 -467 13402 -70
rect 13508 -467 13514 -70
rect 13396 -479 13514 -467
rect 13630 -70 13748 -58
rect 13630 -467 13636 -70
rect 13742 -467 13748 -70
rect 13630 -479 13748 -467
rect 13864 -70 13982 -58
rect 13864 -467 13870 -70
rect 13976 -467 13982 -70
rect 13864 -479 13982 -467
rect 14098 -70 14216 -58
rect 14098 -467 14104 -70
rect 14210 -467 14216 -70
rect 14098 -479 14216 -467
rect 14332 -70 14450 -58
rect 14332 -467 14338 -70
rect 14444 -467 14450 -70
rect 14332 -479 14450 -467
rect 14566 -70 14684 -58
rect 14566 -467 14572 -70
rect 14678 -467 14684 -70
rect 14566 -479 14684 -467
rect 14800 -70 14918 -58
rect 14800 -467 14806 -70
rect 14912 -467 14918 -70
rect 14800 -479 14918 -467
rect 15034 -70 15152 -58
rect 15034 -467 15040 -70
rect 15146 -467 15152 -70
rect 15034 -479 15152 -467
rect 15268 -70 15386 -58
rect 15268 -467 15274 -70
rect 15380 -467 15386 -70
rect 15268 -479 15386 -467
rect 15502 -70 15620 -58
rect 15502 -467 15508 -70
rect 15614 -467 15620 -70
rect 15502 -479 15620 -467
rect 15736 -70 15854 -58
rect 15736 -467 15742 -70
rect 15848 -467 15854 -70
rect 15736 -479 15854 -467
rect 15970 -70 16088 -58
rect 15970 -467 15976 -70
rect 16082 -467 16088 -70
rect 15970 -479 16088 -467
rect 16204 -70 16322 -58
rect 16204 -467 16210 -70
rect 16316 -467 16322 -70
rect 16204 -479 16322 -467
rect 16438 -70 16556 -58
rect 16438 -467 16444 -70
rect 16550 -467 16556 -70
rect 16438 -479 16556 -467
rect 16672 -70 16790 -58
rect 16672 -467 16678 -70
rect 16784 -467 16790 -70
rect 16672 -479 16790 -467
rect 16906 -70 17024 -58
rect 16906 -467 16912 -70
rect 17018 -467 17024 -70
rect 16906 -479 17024 -467
rect 17140 -70 17258 -58
rect 17140 -467 17146 -70
rect 17252 -467 17258 -70
rect 17140 -479 17258 -467
rect 17374 -70 17492 -58
rect 17374 -467 17380 -70
rect 17486 -467 17492 -70
rect 17374 -479 17492 -467
rect 17608 -70 17726 -58
rect 17608 -467 17614 -70
rect 17720 -467 17726 -70
rect 17608 -479 17726 -467
rect 17842 -70 17960 -58
rect 17842 -467 17848 -70
rect 17954 -467 17960 -70
rect 17842 -479 17960 -467
rect 18076 -70 18194 -58
rect 18076 -467 18082 -70
rect 18188 -467 18194 -70
rect 18076 -479 18194 -467
rect 18310 -70 18428 -58
rect 18310 -467 18316 -70
rect 18422 -467 18428 -70
rect 18310 -479 18428 -467
rect 18544 -70 18662 -58
rect 18544 -467 18550 -70
rect 18656 -467 18662 -70
rect 18544 -479 18662 -467
rect 18778 -70 18896 -58
rect 18778 -467 18784 -70
rect 18890 -467 18896 -70
rect 18778 -479 18896 -467
rect 19012 -70 19130 -58
rect 19012 -467 19018 -70
rect 19124 -467 19130 -70
rect 19012 -479 19130 -467
rect 19246 -70 19364 -58
rect 19246 -467 19252 -70
rect 19358 -467 19364 -70
rect 19246 -479 19364 -467
rect 19480 -70 19598 -58
rect 19480 -467 19486 -70
rect 19592 -467 19598 -70
rect 19480 -479 19598 -467
rect 19714 -70 19832 -58
rect 19714 -467 19720 -70
rect 19826 -467 19832 -70
rect 19714 -479 19832 -467
rect 19948 -70 20066 -58
rect 19948 -467 19954 -70
rect 20060 -467 20066 -70
rect 19948 -479 20066 -467
rect 20182 -70 20300 -58
rect 20182 -467 20188 -70
rect 20294 -467 20300 -70
rect 20182 -479 20300 -467
rect 20416 -70 20534 -58
rect 20416 -467 20422 -70
rect 20528 -467 20534 -70
rect 20416 -479 20534 -467
rect 20650 -70 20768 -58
rect 20650 -467 20656 -70
rect 20762 -467 20768 -70
rect 20650 -479 20768 -467
rect 20884 -70 21002 -58
rect 20884 -467 20890 -70
rect 20996 -467 21002 -70
rect 20884 -479 21002 -467
rect 21118 -70 21236 -58
rect 21118 -467 21124 -70
rect 21230 -467 21236 -70
rect 21118 -479 21236 -467
rect 21352 -70 21470 -58
rect 21352 -467 21358 -70
rect 21464 -467 21470 -70
rect 21352 -479 21470 -467
rect 21586 -70 21704 -58
rect 21586 -467 21592 -70
rect 21698 -467 21704 -70
rect 21586 -479 21704 -467
rect 21820 -70 21938 -58
rect 21820 -467 21826 -70
rect 21932 -467 21938 -70
rect 21820 -479 21938 -467
rect 22054 -70 22172 -58
rect 22054 -467 22060 -70
rect 22166 -467 22172 -70
rect 22054 -479 22172 -467
rect 22288 -70 22406 -58
rect 22288 -467 22294 -70
rect 22400 -467 22406 -70
rect 22288 -479 22406 -467
rect 22522 -70 22640 -58
rect 22522 -467 22528 -70
rect 22634 -467 22640 -70
rect 22522 -479 22640 -467
rect 22756 -70 22874 -58
rect 22756 -467 22762 -70
rect 22868 -467 22874 -70
rect 22756 -479 22874 -467
rect 22990 -70 23108 -58
rect 22990 -467 22996 -70
rect 23102 -467 23108 -70
rect 22990 -479 23108 -467
rect 23224 -70 23342 -58
rect 23224 -467 23230 -70
rect 23336 -467 23342 -70
rect 23224 -479 23342 -467
rect 23458 -70 23576 -58
rect 23458 -467 23464 -70
rect 23570 -467 23576 -70
rect 23458 -479 23576 -467
rect 23692 -70 23810 -58
rect 23692 -467 23698 -70
rect 23804 -467 23810 -70
rect 23692 -479 23810 -467
rect 23926 -70 24044 -58
rect 23926 -467 23932 -70
rect 24038 -467 24044 -70
rect 23926 -479 24044 -467
rect 24160 -70 24278 -58
rect 24160 -467 24166 -70
rect 24272 -467 24278 -70
rect 24160 -479 24278 -467
rect 24394 -70 24512 -58
rect 24394 -467 24400 -70
rect 24506 -467 24512 -70
rect 24394 -479 24512 -467
rect 24628 -70 24746 -58
rect 24628 -467 24634 -70
rect 24740 -467 24746 -70
rect 24628 -479 24746 -467
rect 24862 -70 24980 -58
rect 24862 -467 24868 -70
rect 24974 -467 24980 -70
rect 24862 -479 24980 -467
rect 25096 -70 25214 -58
rect 25096 -467 25102 -70
rect 25208 -467 25214 -70
rect 25096 -479 25214 -467
rect 25330 -70 25448 -58
rect 25330 -467 25336 -70
rect 25442 -467 25448 -70
rect 25330 -479 25448 -467
rect 25564 -70 25682 -58
rect 25564 -467 25570 -70
rect 25676 -467 25682 -70
rect 25564 -479 25682 -467
rect 25798 -70 25916 -58
rect 25798 -467 25804 -70
rect 25910 -467 25916 -70
rect 25798 -479 25916 -467
rect 26032 -70 26150 -58
rect 26032 -467 26038 -70
rect 26144 -467 26150 -70
rect 26032 -479 26150 -467
rect 26266 -70 26384 -58
rect 26266 -467 26272 -70
rect 26378 -467 26384 -70
rect 26266 -479 26384 -467
rect 26500 -70 26618 -58
rect 26500 -467 26506 -70
rect 26612 -467 26618 -70
rect 26500 -479 26618 -467
rect 26734 -70 26852 -58
rect 26734 -467 26740 -70
rect 26846 -467 26852 -70
rect 26734 -479 26852 -467
rect 26968 -70 27086 -58
rect 26968 -467 26974 -70
rect 27080 -467 27086 -70
rect 26968 -479 27086 -467
rect 27202 -70 27320 -58
rect 27202 -467 27208 -70
rect 27314 -467 27320 -70
rect 27202 -479 27320 -467
rect 27436 -70 27554 -58
rect 27436 -467 27442 -70
rect 27548 -467 27554 -70
rect 27436 -479 27554 -467
rect 27670 -70 27788 -58
rect 27670 -467 27676 -70
rect 27782 -467 27788 -70
rect 27670 -479 27788 -467
rect 27904 -70 28022 -58
rect 27904 -467 27910 -70
rect 28016 -467 28022 -70
rect 27904 -479 28022 -467
rect 28138 -70 28256 -58
rect 28138 -467 28144 -70
rect 28250 -467 28256 -70
rect 28138 -479 28256 -467
rect 28372 -70 28490 -58
rect 28372 -467 28378 -70
rect 28484 -467 28490 -70
rect 28372 -479 28490 -467
rect 28606 -70 28724 -58
rect 28606 -467 28612 -70
rect 28718 -467 28724 -70
rect 28606 -479 28724 -467
rect 28840 -70 28958 -58
rect 28840 -467 28846 -70
rect 28952 -467 28958 -70
rect 28840 -479 28958 -467
rect 29074 -70 29192 -58
rect 29074 -467 29080 -70
rect 29186 -467 29192 -70
rect 29074 -479 29192 -467
rect 29308 -70 29426 -58
rect 29308 -467 29314 -70
rect 29420 -467 29426 -70
rect 29308 -479 29426 -467
rect 29542 -70 29660 -58
rect 29542 -467 29548 -70
rect 29654 -467 29660 -70
rect 29542 -479 29660 -467
rect 29776 -70 29894 -58
rect 29776 -467 29782 -70
rect 29888 -467 29894 -70
rect 29776 -479 29894 -467
rect -29894 -7469 -29776 -7457
rect -29894 -7866 -29888 -7469
rect -29782 -7866 -29776 -7469
rect -29894 -7878 -29776 -7866
rect -29660 -7469 -29542 -7457
rect -29660 -7866 -29654 -7469
rect -29548 -7866 -29542 -7469
rect -29660 -7878 -29542 -7866
rect -29426 -7469 -29308 -7457
rect -29426 -7866 -29420 -7469
rect -29314 -7866 -29308 -7469
rect -29426 -7878 -29308 -7866
rect -29192 -7469 -29074 -7457
rect -29192 -7866 -29186 -7469
rect -29080 -7866 -29074 -7469
rect -29192 -7878 -29074 -7866
rect -28958 -7469 -28840 -7457
rect -28958 -7866 -28952 -7469
rect -28846 -7866 -28840 -7469
rect -28958 -7878 -28840 -7866
rect -28724 -7469 -28606 -7457
rect -28724 -7866 -28718 -7469
rect -28612 -7866 -28606 -7469
rect -28724 -7878 -28606 -7866
rect -28490 -7469 -28372 -7457
rect -28490 -7866 -28484 -7469
rect -28378 -7866 -28372 -7469
rect -28490 -7878 -28372 -7866
rect -28256 -7469 -28138 -7457
rect -28256 -7866 -28250 -7469
rect -28144 -7866 -28138 -7469
rect -28256 -7878 -28138 -7866
rect -28022 -7469 -27904 -7457
rect -28022 -7866 -28016 -7469
rect -27910 -7866 -27904 -7469
rect -28022 -7878 -27904 -7866
rect -27788 -7469 -27670 -7457
rect -27788 -7866 -27782 -7469
rect -27676 -7866 -27670 -7469
rect -27788 -7878 -27670 -7866
rect -27554 -7469 -27436 -7457
rect -27554 -7866 -27548 -7469
rect -27442 -7866 -27436 -7469
rect -27554 -7878 -27436 -7866
rect -27320 -7469 -27202 -7457
rect -27320 -7866 -27314 -7469
rect -27208 -7866 -27202 -7469
rect -27320 -7878 -27202 -7866
rect -27086 -7469 -26968 -7457
rect -27086 -7866 -27080 -7469
rect -26974 -7866 -26968 -7469
rect -27086 -7878 -26968 -7866
rect -26852 -7469 -26734 -7457
rect -26852 -7866 -26846 -7469
rect -26740 -7866 -26734 -7469
rect -26852 -7878 -26734 -7866
rect -26618 -7469 -26500 -7457
rect -26618 -7866 -26612 -7469
rect -26506 -7866 -26500 -7469
rect -26618 -7878 -26500 -7866
rect -26384 -7469 -26266 -7457
rect -26384 -7866 -26378 -7469
rect -26272 -7866 -26266 -7469
rect -26384 -7878 -26266 -7866
rect -26150 -7469 -26032 -7457
rect -26150 -7866 -26144 -7469
rect -26038 -7866 -26032 -7469
rect -26150 -7878 -26032 -7866
rect -25916 -7469 -25798 -7457
rect -25916 -7866 -25910 -7469
rect -25804 -7866 -25798 -7469
rect -25916 -7878 -25798 -7866
rect -25682 -7469 -25564 -7457
rect -25682 -7866 -25676 -7469
rect -25570 -7866 -25564 -7469
rect -25682 -7878 -25564 -7866
rect -25448 -7469 -25330 -7457
rect -25448 -7866 -25442 -7469
rect -25336 -7866 -25330 -7469
rect -25448 -7878 -25330 -7866
rect -25214 -7469 -25096 -7457
rect -25214 -7866 -25208 -7469
rect -25102 -7866 -25096 -7469
rect -25214 -7878 -25096 -7866
rect -24980 -7469 -24862 -7457
rect -24980 -7866 -24974 -7469
rect -24868 -7866 -24862 -7469
rect -24980 -7878 -24862 -7866
rect -24746 -7469 -24628 -7457
rect -24746 -7866 -24740 -7469
rect -24634 -7866 -24628 -7469
rect -24746 -7878 -24628 -7866
rect -24512 -7469 -24394 -7457
rect -24512 -7866 -24506 -7469
rect -24400 -7866 -24394 -7469
rect -24512 -7878 -24394 -7866
rect -24278 -7469 -24160 -7457
rect -24278 -7866 -24272 -7469
rect -24166 -7866 -24160 -7469
rect -24278 -7878 -24160 -7866
rect -24044 -7469 -23926 -7457
rect -24044 -7866 -24038 -7469
rect -23932 -7866 -23926 -7469
rect -24044 -7878 -23926 -7866
rect -23810 -7469 -23692 -7457
rect -23810 -7866 -23804 -7469
rect -23698 -7866 -23692 -7469
rect -23810 -7878 -23692 -7866
rect -23576 -7469 -23458 -7457
rect -23576 -7866 -23570 -7469
rect -23464 -7866 -23458 -7469
rect -23576 -7878 -23458 -7866
rect -23342 -7469 -23224 -7457
rect -23342 -7866 -23336 -7469
rect -23230 -7866 -23224 -7469
rect -23342 -7878 -23224 -7866
rect -23108 -7469 -22990 -7457
rect -23108 -7866 -23102 -7469
rect -22996 -7866 -22990 -7469
rect -23108 -7878 -22990 -7866
rect -22874 -7469 -22756 -7457
rect -22874 -7866 -22868 -7469
rect -22762 -7866 -22756 -7469
rect -22874 -7878 -22756 -7866
rect -22640 -7469 -22522 -7457
rect -22640 -7866 -22634 -7469
rect -22528 -7866 -22522 -7469
rect -22640 -7878 -22522 -7866
rect -22406 -7469 -22288 -7457
rect -22406 -7866 -22400 -7469
rect -22294 -7866 -22288 -7469
rect -22406 -7878 -22288 -7866
rect -22172 -7469 -22054 -7457
rect -22172 -7866 -22166 -7469
rect -22060 -7866 -22054 -7469
rect -22172 -7878 -22054 -7866
rect -21938 -7469 -21820 -7457
rect -21938 -7866 -21932 -7469
rect -21826 -7866 -21820 -7469
rect -21938 -7878 -21820 -7866
rect -21704 -7469 -21586 -7457
rect -21704 -7866 -21698 -7469
rect -21592 -7866 -21586 -7469
rect -21704 -7878 -21586 -7866
rect -21470 -7469 -21352 -7457
rect -21470 -7866 -21464 -7469
rect -21358 -7866 -21352 -7469
rect -21470 -7878 -21352 -7866
rect -21236 -7469 -21118 -7457
rect -21236 -7866 -21230 -7469
rect -21124 -7866 -21118 -7469
rect -21236 -7878 -21118 -7866
rect -21002 -7469 -20884 -7457
rect -21002 -7866 -20996 -7469
rect -20890 -7866 -20884 -7469
rect -21002 -7878 -20884 -7866
rect -20768 -7469 -20650 -7457
rect -20768 -7866 -20762 -7469
rect -20656 -7866 -20650 -7469
rect -20768 -7878 -20650 -7866
rect -20534 -7469 -20416 -7457
rect -20534 -7866 -20528 -7469
rect -20422 -7866 -20416 -7469
rect -20534 -7878 -20416 -7866
rect -20300 -7469 -20182 -7457
rect -20300 -7866 -20294 -7469
rect -20188 -7866 -20182 -7469
rect -20300 -7878 -20182 -7866
rect -20066 -7469 -19948 -7457
rect -20066 -7866 -20060 -7469
rect -19954 -7866 -19948 -7469
rect -20066 -7878 -19948 -7866
rect -19832 -7469 -19714 -7457
rect -19832 -7866 -19826 -7469
rect -19720 -7866 -19714 -7469
rect -19832 -7878 -19714 -7866
rect -19598 -7469 -19480 -7457
rect -19598 -7866 -19592 -7469
rect -19486 -7866 -19480 -7469
rect -19598 -7878 -19480 -7866
rect -19364 -7469 -19246 -7457
rect -19364 -7866 -19358 -7469
rect -19252 -7866 -19246 -7469
rect -19364 -7878 -19246 -7866
rect -19130 -7469 -19012 -7457
rect -19130 -7866 -19124 -7469
rect -19018 -7866 -19012 -7469
rect -19130 -7878 -19012 -7866
rect -18896 -7469 -18778 -7457
rect -18896 -7866 -18890 -7469
rect -18784 -7866 -18778 -7469
rect -18896 -7878 -18778 -7866
rect -18662 -7469 -18544 -7457
rect -18662 -7866 -18656 -7469
rect -18550 -7866 -18544 -7469
rect -18662 -7878 -18544 -7866
rect -18428 -7469 -18310 -7457
rect -18428 -7866 -18422 -7469
rect -18316 -7866 -18310 -7469
rect -18428 -7878 -18310 -7866
rect -18194 -7469 -18076 -7457
rect -18194 -7866 -18188 -7469
rect -18082 -7866 -18076 -7469
rect -18194 -7878 -18076 -7866
rect -17960 -7469 -17842 -7457
rect -17960 -7866 -17954 -7469
rect -17848 -7866 -17842 -7469
rect -17960 -7878 -17842 -7866
rect -17726 -7469 -17608 -7457
rect -17726 -7866 -17720 -7469
rect -17614 -7866 -17608 -7469
rect -17726 -7878 -17608 -7866
rect -17492 -7469 -17374 -7457
rect -17492 -7866 -17486 -7469
rect -17380 -7866 -17374 -7469
rect -17492 -7878 -17374 -7866
rect -17258 -7469 -17140 -7457
rect -17258 -7866 -17252 -7469
rect -17146 -7866 -17140 -7469
rect -17258 -7878 -17140 -7866
rect -17024 -7469 -16906 -7457
rect -17024 -7866 -17018 -7469
rect -16912 -7866 -16906 -7469
rect -17024 -7878 -16906 -7866
rect -16790 -7469 -16672 -7457
rect -16790 -7866 -16784 -7469
rect -16678 -7866 -16672 -7469
rect -16790 -7878 -16672 -7866
rect -16556 -7469 -16438 -7457
rect -16556 -7866 -16550 -7469
rect -16444 -7866 -16438 -7469
rect -16556 -7878 -16438 -7866
rect -16322 -7469 -16204 -7457
rect -16322 -7866 -16316 -7469
rect -16210 -7866 -16204 -7469
rect -16322 -7878 -16204 -7866
rect -16088 -7469 -15970 -7457
rect -16088 -7866 -16082 -7469
rect -15976 -7866 -15970 -7469
rect -16088 -7878 -15970 -7866
rect -15854 -7469 -15736 -7457
rect -15854 -7866 -15848 -7469
rect -15742 -7866 -15736 -7469
rect -15854 -7878 -15736 -7866
rect -15620 -7469 -15502 -7457
rect -15620 -7866 -15614 -7469
rect -15508 -7866 -15502 -7469
rect -15620 -7878 -15502 -7866
rect -15386 -7469 -15268 -7457
rect -15386 -7866 -15380 -7469
rect -15274 -7866 -15268 -7469
rect -15386 -7878 -15268 -7866
rect -15152 -7469 -15034 -7457
rect -15152 -7866 -15146 -7469
rect -15040 -7866 -15034 -7469
rect -15152 -7878 -15034 -7866
rect -14918 -7469 -14800 -7457
rect -14918 -7866 -14912 -7469
rect -14806 -7866 -14800 -7469
rect -14918 -7878 -14800 -7866
rect -14684 -7469 -14566 -7457
rect -14684 -7866 -14678 -7469
rect -14572 -7866 -14566 -7469
rect -14684 -7878 -14566 -7866
rect -14450 -7469 -14332 -7457
rect -14450 -7866 -14444 -7469
rect -14338 -7866 -14332 -7469
rect -14450 -7878 -14332 -7866
rect -14216 -7469 -14098 -7457
rect -14216 -7866 -14210 -7469
rect -14104 -7866 -14098 -7469
rect -14216 -7878 -14098 -7866
rect -13982 -7469 -13864 -7457
rect -13982 -7866 -13976 -7469
rect -13870 -7866 -13864 -7469
rect -13982 -7878 -13864 -7866
rect -13748 -7469 -13630 -7457
rect -13748 -7866 -13742 -7469
rect -13636 -7866 -13630 -7469
rect -13748 -7878 -13630 -7866
rect -13514 -7469 -13396 -7457
rect -13514 -7866 -13508 -7469
rect -13402 -7866 -13396 -7469
rect -13514 -7878 -13396 -7866
rect -13280 -7469 -13162 -7457
rect -13280 -7866 -13274 -7469
rect -13168 -7866 -13162 -7469
rect -13280 -7878 -13162 -7866
rect -13046 -7469 -12928 -7457
rect -13046 -7866 -13040 -7469
rect -12934 -7866 -12928 -7469
rect -13046 -7878 -12928 -7866
rect -12812 -7469 -12694 -7457
rect -12812 -7866 -12806 -7469
rect -12700 -7866 -12694 -7469
rect -12812 -7878 -12694 -7866
rect -12578 -7469 -12460 -7457
rect -12578 -7866 -12572 -7469
rect -12466 -7866 -12460 -7469
rect -12578 -7878 -12460 -7866
rect -12344 -7469 -12226 -7457
rect -12344 -7866 -12338 -7469
rect -12232 -7866 -12226 -7469
rect -12344 -7878 -12226 -7866
rect -12110 -7469 -11992 -7457
rect -12110 -7866 -12104 -7469
rect -11998 -7866 -11992 -7469
rect -12110 -7878 -11992 -7866
rect -11876 -7469 -11758 -7457
rect -11876 -7866 -11870 -7469
rect -11764 -7866 -11758 -7469
rect -11876 -7878 -11758 -7866
rect -11642 -7469 -11524 -7457
rect -11642 -7866 -11636 -7469
rect -11530 -7866 -11524 -7469
rect -11642 -7878 -11524 -7866
rect -11408 -7469 -11290 -7457
rect -11408 -7866 -11402 -7469
rect -11296 -7866 -11290 -7469
rect -11408 -7878 -11290 -7866
rect -11174 -7469 -11056 -7457
rect -11174 -7866 -11168 -7469
rect -11062 -7866 -11056 -7469
rect -11174 -7878 -11056 -7866
rect -10940 -7469 -10822 -7457
rect -10940 -7866 -10934 -7469
rect -10828 -7866 -10822 -7469
rect -10940 -7878 -10822 -7866
rect -10706 -7469 -10588 -7457
rect -10706 -7866 -10700 -7469
rect -10594 -7866 -10588 -7469
rect -10706 -7878 -10588 -7866
rect -10472 -7469 -10354 -7457
rect -10472 -7866 -10466 -7469
rect -10360 -7866 -10354 -7469
rect -10472 -7878 -10354 -7866
rect -10238 -7469 -10120 -7457
rect -10238 -7866 -10232 -7469
rect -10126 -7866 -10120 -7469
rect -10238 -7878 -10120 -7866
rect -10004 -7469 -9886 -7457
rect -10004 -7866 -9998 -7469
rect -9892 -7866 -9886 -7469
rect -10004 -7878 -9886 -7866
rect -9770 -7469 -9652 -7457
rect -9770 -7866 -9764 -7469
rect -9658 -7866 -9652 -7469
rect -9770 -7878 -9652 -7866
rect -9536 -7469 -9418 -7457
rect -9536 -7866 -9530 -7469
rect -9424 -7866 -9418 -7469
rect -9536 -7878 -9418 -7866
rect -9302 -7469 -9184 -7457
rect -9302 -7866 -9296 -7469
rect -9190 -7866 -9184 -7469
rect -9302 -7878 -9184 -7866
rect -9068 -7469 -8950 -7457
rect -9068 -7866 -9062 -7469
rect -8956 -7866 -8950 -7469
rect -9068 -7878 -8950 -7866
rect -8834 -7469 -8716 -7457
rect -8834 -7866 -8828 -7469
rect -8722 -7866 -8716 -7469
rect -8834 -7878 -8716 -7866
rect -8600 -7469 -8482 -7457
rect -8600 -7866 -8594 -7469
rect -8488 -7866 -8482 -7469
rect -8600 -7878 -8482 -7866
rect -8366 -7469 -8248 -7457
rect -8366 -7866 -8360 -7469
rect -8254 -7866 -8248 -7469
rect -8366 -7878 -8248 -7866
rect -8132 -7469 -8014 -7457
rect -8132 -7866 -8126 -7469
rect -8020 -7866 -8014 -7469
rect -8132 -7878 -8014 -7866
rect -7898 -7469 -7780 -7457
rect -7898 -7866 -7892 -7469
rect -7786 -7866 -7780 -7469
rect -7898 -7878 -7780 -7866
rect -7664 -7469 -7546 -7457
rect -7664 -7866 -7658 -7469
rect -7552 -7866 -7546 -7469
rect -7664 -7878 -7546 -7866
rect -7430 -7469 -7312 -7457
rect -7430 -7866 -7424 -7469
rect -7318 -7866 -7312 -7469
rect -7430 -7878 -7312 -7866
rect -7196 -7469 -7078 -7457
rect -7196 -7866 -7190 -7469
rect -7084 -7866 -7078 -7469
rect -7196 -7878 -7078 -7866
rect -6962 -7469 -6844 -7457
rect -6962 -7866 -6956 -7469
rect -6850 -7866 -6844 -7469
rect -6962 -7878 -6844 -7866
rect -6728 -7469 -6610 -7457
rect -6728 -7866 -6722 -7469
rect -6616 -7866 -6610 -7469
rect -6728 -7878 -6610 -7866
rect -6494 -7469 -6376 -7457
rect -6494 -7866 -6488 -7469
rect -6382 -7866 -6376 -7469
rect -6494 -7878 -6376 -7866
rect -6260 -7469 -6142 -7457
rect -6260 -7866 -6254 -7469
rect -6148 -7866 -6142 -7469
rect -6260 -7878 -6142 -7866
rect -6026 -7469 -5908 -7457
rect -6026 -7866 -6020 -7469
rect -5914 -7866 -5908 -7469
rect -6026 -7878 -5908 -7866
rect -5792 -7469 -5674 -7457
rect -5792 -7866 -5786 -7469
rect -5680 -7866 -5674 -7469
rect -5792 -7878 -5674 -7866
rect -5558 -7469 -5440 -7457
rect -5558 -7866 -5552 -7469
rect -5446 -7866 -5440 -7469
rect -5558 -7878 -5440 -7866
rect -5324 -7469 -5206 -7457
rect -5324 -7866 -5318 -7469
rect -5212 -7866 -5206 -7469
rect -5324 -7878 -5206 -7866
rect -5090 -7469 -4972 -7457
rect -5090 -7866 -5084 -7469
rect -4978 -7866 -4972 -7469
rect -5090 -7878 -4972 -7866
rect -4856 -7469 -4738 -7457
rect -4856 -7866 -4850 -7469
rect -4744 -7866 -4738 -7469
rect -4856 -7878 -4738 -7866
rect -4622 -7469 -4504 -7457
rect -4622 -7866 -4616 -7469
rect -4510 -7866 -4504 -7469
rect -4622 -7878 -4504 -7866
rect -4388 -7469 -4270 -7457
rect -4388 -7866 -4382 -7469
rect -4276 -7866 -4270 -7469
rect -4388 -7878 -4270 -7866
rect -4154 -7469 -4036 -7457
rect -4154 -7866 -4148 -7469
rect -4042 -7866 -4036 -7469
rect -4154 -7878 -4036 -7866
rect -3920 -7469 -3802 -7457
rect -3920 -7866 -3914 -7469
rect -3808 -7866 -3802 -7469
rect -3920 -7878 -3802 -7866
rect -3686 -7469 -3568 -7457
rect -3686 -7866 -3680 -7469
rect -3574 -7866 -3568 -7469
rect -3686 -7878 -3568 -7866
rect -3452 -7469 -3334 -7457
rect -3452 -7866 -3446 -7469
rect -3340 -7866 -3334 -7469
rect -3452 -7878 -3334 -7866
rect -3218 -7469 -3100 -7457
rect -3218 -7866 -3212 -7469
rect -3106 -7866 -3100 -7469
rect -3218 -7878 -3100 -7866
rect -2984 -7469 -2866 -7457
rect -2984 -7866 -2978 -7469
rect -2872 -7866 -2866 -7469
rect -2984 -7878 -2866 -7866
rect -2750 -7469 -2632 -7457
rect -2750 -7866 -2744 -7469
rect -2638 -7866 -2632 -7469
rect -2750 -7878 -2632 -7866
rect -2516 -7469 -2398 -7457
rect -2516 -7866 -2510 -7469
rect -2404 -7866 -2398 -7469
rect -2516 -7878 -2398 -7866
rect -2282 -7469 -2164 -7457
rect -2282 -7866 -2276 -7469
rect -2170 -7866 -2164 -7469
rect -2282 -7878 -2164 -7866
rect -2048 -7469 -1930 -7457
rect -2048 -7866 -2042 -7469
rect -1936 -7866 -1930 -7469
rect -2048 -7878 -1930 -7866
rect -1814 -7469 -1696 -7457
rect -1814 -7866 -1808 -7469
rect -1702 -7866 -1696 -7469
rect -1814 -7878 -1696 -7866
rect -1580 -7469 -1462 -7457
rect -1580 -7866 -1574 -7469
rect -1468 -7866 -1462 -7469
rect -1580 -7878 -1462 -7866
rect -1346 -7469 -1228 -7457
rect -1346 -7866 -1340 -7469
rect -1234 -7866 -1228 -7469
rect -1346 -7878 -1228 -7866
rect -1112 -7469 -994 -7457
rect -1112 -7866 -1106 -7469
rect -1000 -7866 -994 -7469
rect -1112 -7878 -994 -7866
rect -878 -7469 -760 -7457
rect -878 -7866 -872 -7469
rect -766 -7866 -760 -7469
rect -878 -7878 -760 -7866
rect -644 -7469 -526 -7457
rect -644 -7866 -638 -7469
rect -532 -7866 -526 -7469
rect -644 -7878 -526 -7866
rect -410 -7469 -292 -7457
rect -410 -7866 -404 -7469
rect -298 -7866 -292 -7469
rect -410 -7878 -292 -7866
rect -176 -7469 -58 -7457
rect -176 -7866 -170 -7469
rect -64 -7866 -58 -7469
rect -176 -7878 -58 -7866
rect 58 -7469 176 -7457
rect 58 -7866 64 -7469
rect 170 -7866 176 -7469
rect 58 -7878 176 -7866
rect 292 -7469 410 -7457
rect 292 -7866 298 -7469
rect 404 -7866 410 -7469
rect 292 -7878 410 -7866
rect 526 -7469 644 -7457
rect 526 -7866 532 -7469
rect 638 -7866 644 -7469
rect 526 -7878 644 -7866
rect 760 -7469 878 -7457
rect 760 -7866 766 -7469
rect 872 -7866 878 -7469
rect 760 -7878 878 -7866
rect 994 -7469 1112 -7457
rect 994 -7866 1000 -7469
rect 1106 -7866 1112 -7469
rect 994 -7878 1112 -7866
rect 1228 -7469 1346 -7457
rect 1228 -7866 1234 -7469
rect 1340 -7866 1346 -7469
rect 1228 -7878 1346 -7866
rect 1462 -7469 1580 -7457
rect 1462 -7866 1468 -7469
rect 1574 -7866 1580 -7469
rect 1462 -7878 1580 -7866
rect 1696 -7469 1814 -7457
rect 1696 -7866 1702 -7469
rect 1808 -7866 1814 -7469
rect 1696 -7878 1814 -7866
rect 1930 -7469 2048 -7457
rect 1930 -7866 1936 -7469
rect 2042 -7866 2048 -7469
rect 1930 -7878 2048 -7866
rect 2164 -7469 2282 -7457
rect 2164 -7866 2170 -7469
rect 2276 -7866 2282 -7469
rect 2164 -7878 2282 -7866
rect 2398 -7469 2516 -7457
rect 2398 -7866 2404 -7469
rect 2510 -7866 2516 -7469
rect 2398 -7878 2516 -7866
rect 2632 -7469 2750 -7457
rect 2632 -7866 2638 -7469
rect 2744 -7866 2750 -7469
rect 2632 -7878 2750 -7866
rect 2866 -7469 2984 -7457
rect 2866 -7866 2872 -7469
rect 2978 -7866 2984 -7469
rect 2866 -7878 2984 -7866
rect 3100 -7469 3218 -7457
rect 3100 -7866 3106 -7469
rect 3212 -7866 3218 -7469
rect 3100 -7878 3218 -7866
rect 3334 -7469 3452 -7457
rect 3334 -7866 3340 -7469
rect 3446 -7866 3452 -7469
rect 3334 -7878 3452 -7866
rect 3568 -7469 3686 -7457
rect 3568 -7866 3574 -7469
rect 3680 -7866 3686 -7469
rect 3568 -7878 3686 -7866
rect 3802 -7469 3920 -7457
rect 3802 -7866 3808 -7469
rect 3914 -7866 3920 -7469
rect 3802 -7878 3920 -7866
rect 4036 -7469 4154 -7457
rect 4036 -7866 4042 -7469
rect 4148 -7866 4154 -7469
rect 4036 -7878 4154 -7866
rect 4270 -7469 4388 -7457
rect 4270 -7866 4276 -7469
rect 4382 -7866 4388 -7469
rect 4270 -7878 4388 -7866
rect 4504 -7469 4622 -7457
rect 4504 -7866 4510 -7469
rect 4616 -7866 4622 -7469
rect 4504 -7878 4622 -7866
rect 4738 -7469 4856 -7457
rect 4738 -7866 4744 -7469
rect 4850 -7866 4856 -7469
rect 4738 -7878 4856 -7866
rect 4972 -7469 5090 -7457
rect 4972 -7866 4978 -7469
rect 5084 -7866 5090 -7469
rect 4972 -7878 5090 -7866
rect 5206 -7469 5324 -7457
rect 5206 -7866 5212 -7469
rect 5318 -7866 5324 -7469
rect 5206 -7878 5324 -7866
rect 5440 -7469 5558 -7457
rect 5440 -7866 5446 -7469
rect 5552 -7866 5558 -7469
rect 5440 -7878 5558 -7866
rect 5674 -7469 5792 -7457
rect 5674 -7866 5680 -7469
rect 5786 -7866 5792 -7469
rect 5674 -7878 5792 -7866
rect 5908 -7469 6026 -7457
rect 5908 -7866 5914 -7469
rect 6020 -7866 6026 -7469
rect 5908 -7878 6026 -7866
rect 6142 -7469 6260 -7457
rect 6142 -7866 6148 -7469
rect 6254 -7866 6260 -7469
rect 6142 -7878 6260 -7866
rect 6376 -7469 6494 -7457
rect 6376 -7866 6382 -7469
rect 6488 -7866 6494 -7469
rect 6376 -7878 6494 -7866
rect 6610 -7469 6728 -7457
rect 6610 -7866 6616 -7469
rect 6722 -7866 6728 -7469
rect 6610 -7878 6728 -7866
rect 6844 -7469 6962 -7457
rect 6844 -7866 6850 -7469
rect 6956 -7866 6962 -7469
rect 6844 -7878 6962 -7866
rect 7078 -7469 7196 -7457
rect 7078 -7866 7084 -7469
rect 7190 -7866 7196 -7469
rect 7078 -7878 7196 -7866
rect 7312 -7469 7430 -7457
rect 7312 -7866 7318 -7469
rect 7424 -7866 7430 -7469
rect 7312 -7878 7430 -7866
rect 7546 -7469 7664 -7457
rect 7546 -7866 7552 -7469
rect 7658 -7866 7664 -7469
rect 7546 -7878 7664 -7866
rect 7780 -7469 7898 -7457
rect 7780 -7866 7786 -7469
rect 7892 -7866 7898 -7469
rect 7780 -7878 7898 -7866
rect 8014 -7469 8132 -7457
rect 8014 -7866 8020 -7469
rect 8126 -7866 8132 -7469
rect 8014 -7878 8132 -7866
rect 8248 -7469 8366 -7457
rect 8248 -7866 8254 -7469
rect 8360 -7866 8366 -7469
rect 8248 -7878 8366 -7866
rect 8482 -7469 8600 -7457
rect 8482 -7866 8488 -7469
rect 8594 -7866 8600 -7469
rect 8482 -7878 8600 -7866
rect 8716 -7469 8834 -7457
rect 8716 -7866 8722 -7469
rect 8828 -7866 8834 -7469
rect 8716 -7878 8834 -7866
rect 8950 -7469 9068 -7457
rect 8950 -7866 8956 -7469
rect 9062 -7866 9068 -7469
rect 8950 -7878 9068 -7866
rect 9184 -7469 9302 -7457
rect 9184 -7866 9190 -7469
rect 9296 -7866 9302 -7469
rect 9184 -7878 9302 -7866
rect 9418 -7469 9536 -7457
rect 9418 -7866 9424 -7469
rect 9530 -7866 9536 -7469
rect 9418 -7878 9536 -7866
rect 9652 -7469 9770 -7457
rect 9652 -7866 9658 -7469
rect 9764 -7866 9770 -7469
rect 9652 -7878 9770 -7866
rect 9886 -7469 10004 -7457
rect 9886 -7866 9892 -7469
rect 9998 -7866 10004 -7469
rect 9886 -7878 10004 -7866
rect 10120 -7469 10238 -7457
rect 10120 -7866 10126 -7469
rect 10232 -7866 10238 -7469
rect 10120 -7878 10238 -7866
rect 10354 -7469 10472 -7457
rect 10354 -7866 10360 -7469
rect 10466 -7866 10472 -7469
rect 10354 -7878 10472 -7866
rect 10588 -7469 10706 -7457
rect 10588 -7866 10594 -7469
rect 10700 -7866 10706 -7469
rect 10588 -7878 10706 -7866
rect 10822 -7469 10940 -7457
rect 10822 -7866 10828 -7469
rect 10934 -7866 10940 -7469
rect 10822 -7878 10940 -7866
rect 11056 -7469 11174 -7457
rect 11056 -7866 11062 -7469
rect 11168 -7866 11174 -7469
rect 11056 -7878 11174 -7866
rect 11290 -7469 11408 -7457
rect 11290 -7866 11296 -7469
rect 11402 -7866 11408 -7469
rect 11290 -7878 11408 -7866
rect 11524 -7469 11642 -7457
rect 11524 -7866 11530 -7469
rect 11636 -7866 11642 -7469
rect 11524 -7878 11642 -7866
rect 11758 -7469 11876 -7457
rect 11758 -7866 11764 -7469
rect 11870 -7866 11876 -7469
rect 11758 -7878 11876 -7866
rect 11992 -7469 12110 -7457
rect 11992 -7866 11998 -7469
rect 12104 -7866 12110 -7469
rect 11992 -7878 12110 -7866
rect 12226 -7469 12344 -7457
rect 12226 -7866 12232 -7469
rect 12338 -7866 12344 -7469
rect 12226 -7878 12344 -7866
rect 12460 -7469 12578 -7457
rect 12460 -7866 12466 -7469
rect 12572 -7866 12578 -7469
rect 12460 -7878 12578 -7866
rect 12694 -7469 12812 -7457
rect 12694 -7866 12700 -7469
rect 12806 -7866 12812 -7469
rect 12694 -7878 12812 -7866
rect 12928 -7469 13046 -7457
rect 12928 -7866 12934 -7469
rect 13040 -7866 13046 -7469
rect 12928 -7878 13046 -7866
rect 13162 -7469 13280 -7457
rect 13162 -7866 13168 -7469
rect 13274 -7866 13280 -7469
rect 13162 -7878 13280 -7866
rect 13396 -7469 13514 -7457
rect 13396 -7866 13402 -7469
rect 13508 -7866 13514 -7469
rect 13396 -7878 13514 -7866
rect 13630 -7469 13748 -7457
rect 13630 -7866 13636 -7469
rect 13742 -7866 13748 -7469
rect 13630 -7878 13748 -7866
rect 13864 -7469 13982 -7457
rect 13864 -7866 13870 -7469
rect 13976 -7866 13982 -7469
rect 13864 -7878 13982 -7866
rect 14098 -7469 14216 -7457
rect 14098 -7866 14104 -7469
rect 14210 -7866 14216 -7469
rect 14098 -7878 14216 -7866
rect 14332 -7469 14450 -7457
rect 14332 -7866 14338 -7469
rect 14444 -7866 14450 -7469
rect 14332 -7878 14450 -7866
rect 14566 -7469 14684 -7457
rect 14566 -7866 14572 -7469
rect 14678 -7866 14684 -7469
rect 14566 -7878 14684 -7866
rect 14800 -7469 14918 -7457
rect 14800 -7866 14806 -7469
rect 14912 -7866 14918 -7469
rect 14800 -7878 14918 -7866
rect 15034 -7469 15152 -7457
rect 15034 -7866 15040 -7469
rect 15146 -7866 15152 -7469
rect 15034 -7878 15152 -7866
rect 15268 -7469 15386 -7457
rect 15268 -7866 15274 -7469
rect 15380 -7866 15386 -7469
rect 15268 -7878 15386 -7866
rect 15502 -7469 15620 -7457
rect 15502 -7866 15508 -7469
rect 15614 -7866 15620 -7469
rect 15502 -7878 15620 -7866
rect 15736 -7469 15854 -7457
rect 15736 -7866 15742 -7469
rect 15848 -7866 15854 -7469
rect 15736 -7878 15854 -7866
rect 15970 -7469 16088 -7457
rect 15970 -7866 15976 -7469
rect 16082 -7866 16088 -7469
rect 15970 -7878 16088 -7866
rect 16204 -7469 16322 -7457
rect 16204 -7866 16210 -7469
rect 16316 -7866 16322 -7469
rect 16204 -7878 16322 -7866
rect 16438 -7469 16556 -7457
rect 16438 -7866 16444 -7469
rect 16550 -7866 16556 -7469
rect 16438 -7878 16556 -7866
rect 16672 -7469 16790 -7457
rect 16672 -7866 16678 -7469
rect 16784 -7866 16790 -7469
rect 16672 -7878 16790 -7866
rect 16906 -7469 17024 -7457
rect 16906 -7866 16912 -7469
rect 17018 -7866 17024 -7469
rect 16906 -7878 17024 -7866
rect 17140 -7469 17258 -7457
rect 17140 -7866 17146 -7469
rect 17252 -7866 17258 -7469
rect 17140 -7878 17258 -7866
rect 17374 -7469 17492 -7457
rect 17374 -7866 17380 -7469
rect 17486 -7866 17492 -7469
rect 17374 -7878 17492 -7866
rect 17608 -7469 17726 -7457
rect 17608 -7866 17614 -7469
rect 17720 -7866 17726 -7469
rect 17608 -7878 17726 -7866
rect 17842 -7469 17960 -7457
rect 17842 -7866 17848 -7469
rect 17954 -7866 17960 -7469
rect 17842 -7878 17960 -7866
rect 18076 -7469 18194 -7457
rect 18076 -7866 18082 -7469
rect 18188 -7866 18194 -7469
rect 18076 -7878 18194 -7866
rect 18310 -7469 18428 -7457
rect 18310 -7866 18316 -7469
rect 18422 -7866 18428 -7469
rect 18310 -7878 18428 -7866
rect 18544 -7469 18662 -7457
rect 18544 -7866 18550 -7469
rect 18656 -7866 18662 -7469
rect 18544 -7878 18662 -7866
rect 18778 -7469 18896 -7457
rect 18778 -7866 18784 -7469
rect 18890 -7866 18896 -7469
rect 18778 -7878 18896 -7866
rect 19012 -7469 19130 -7457
rect 19012 -7866 19018 -7469
rect 19124 -7866 19130 -7469
rect 19012 -7878 19130 -7866
rect 19246 -7469 19364 -7457
rect 19246 -7866 19252 -7469
rect 19358 -7866 19364 -7469
rect 19246 -7878 19364 -7866
rect 19480 -7469 19598 -7457
rect 19480 -7866 19486 -7469
rect 19592 -7866 19598 -7469
rect 19480 -7878 19598 -7866
rect 19714 -7469 19832 -7457
rect 19714 -7866 19720 -7469
rect 19826 -7866 19832 -7469
rect 19714 -7878 19832 -7866
rect 19948 -7469 20066 -7457
rect 19948 -7866 19954 -7469
rect 20060 -7866 20066 -7469
rect 19948 -7878 20066 -7866
rect 20182 -7469 20300 -7457
rect 20182 -7866 20188 -7469
rect 20294 -7866 20300 -7469
rect 20182 -7878 20300 -7866
rect 20416 -7469 20534 -7457
rect 20416 -7866 20422 -7469
rect 20528 -7866 20534 -7469
rect 20416 -7878 20534 -7866
rect 20650 -7469 20768 -7457
rect 20650 -7866 20656 -7469
rect 20762 -7866 20768 -7469
rect 20650 -7878 20768 -7866
rect 20884 -7469 21002 -7457
rect 20884 -7866 20890 -7469
rect 20996 -7866 21002 -7469
rect 20884 -7878 21002 -7866
rect 21118 -7469 21236 -7457
rect 21118 -7866 21124 -7469
rect 21230 -7866 21236 -7469
rect 21118 -7878 21236 -7866
rect 21352 -7469 21470 -7457
rect 21352 -7866 21358 -7469
rect 21464 -7866 21470 -7469
rect 21352 -7878 21470 -7866
rect 21586 -7469 21704 -7457
rect 21586 -7866 21592 -7469
rect 21698 -7866 21704 -7469
rect 21586 -7878 21704 -7866
rect 21820 -7469 21938 -7457
rect 21820 -7866 21826 -7469
rect 21932 -7866 21938 -7469
rect 21820 -7878 21938 -7866
rect 22054 -7469 22172 -7457
rect 22054 -7866 22060 -7469
rect 22166 -7866 22172 -7469
rect 22054 -7878 22172 -7866
rect 22288 -7469 22406 -7457
rect 22288 -7866 22294 -7469
rect 22400 -7866 22406 -7469
rect 22288 -7878 22406 -7866
rect 22522 -7469 22640 -7457
rect 22522 -7866 22528 -7469
rect 22634 -7866 22640 -7469
rect 22522 -7878 22640 -7866
rect 22756 -7469 22874 -7457
rect 22756 -7866 22762 -7469
rect 22868 -7866 22874 -7469
rect 22756 -7878 22874 -7866
rect 22990 -7469 23108 -7457
rect 22990 -7866 22996 -7469
rect 23102 -7866 23108 -7469
rect 22990 -7878 23108 -7866
rect 23224 -7469 23342 -7457
rect 23224 -7866 23230 -7469
rect 23336 -7866 23342 -7469
rect 23224 -7878 23342 -7866
rect 23458 -7469 23576 -7457
rect 23458 -7866 23464 -7469
rect 23570 -7866 23576 -7469
rect 23458 -7878 23576 -7866
rect 23692 -7469 23810 -7457
rect 23692 -7866 23698 -7469
rect 23804 -7866 23810 -7469
rect 23692 -7878 23810 -7866
rect 23926 -7469 24044 -7457
rect 23926 -7866 23932 -7469
rect 24038 -7866 24044 -7469
rect 23926 -7878 24044 -7866
rect 24160 -7469 24278 -7457
rect 24160 -7866 24166 -7469
rect 24272 -7866 24278 -7469
rect 24160 -7878 24278 -7866
rect 24394 -7469 24512 -7457
rect 24394 -7866 24400 -7469
rect 24506 -7866 24512 -7469
rect 24394 -7878 24512 -7866
rect 24628 -7469 24746 -7457
rect 24628 -7866 24634 -7469
rect 24740 -7866 24746 -7469
rect 24628 -7878 24746 -7866
rect 24862 -7469 24980 -7457
rect 24862 -7866 24868 -7469
rect 24974 -7866 24980 -7469
rect 24862 -7878 24980 -7866
rect 25096 -7469 25214 -7457
rect 25096 -7866 25102 -7469
rect 25208 -7866 25214 -7469
rect 25096 -7878 25214 -7866
rect 25330 -7469 25448 -7457
rect 25330 -7866 25336 -7469
rect 25442 -7866 25448 -7469
rect 25330 -7878 25448 -7866
rect 25564 -7469 25682 -7457
rect 25564 -7866 25570 -7469
rect 25676 -7866 25682 -7469
rect 25564 -7878 25682 -7866
rect 25798 -7469 25916 -7457
rect 25798 -7866 25804 -7469
rect 25910 -7866 25916 -7469
rect 25798 -7878 25916 -7866
rect 26032 -7469 26150 -7457
rect 26032 -7866 26038 -7469
rect 26144 -7866 26150 -7469
rect 26032 -7878 26150 -7866
rect 26266 -7469 26384 -7457
rect 26266 -7866 26272 -7469
rect 26378 -7866 26384 -7469
rect 26266 -7878 26384 -7866
rect 26500 -7469 26618 -7457
rect 26500 -7866 26506 -7469
rect 26612 -7866 26618 -7469
rect 26500 -7878 26618 -7866
rect 26734 -7469 26852 -7457
rect 26734 -7866 26740 -7469
rect 26846 -7866 26852 -7469
rect 26734 -7878 26852 -7866
rect 26968 -7469 27086 -7457
rect 26968 -7866 26974 -7469
rect 27080 -7866 27086 -7469
rect 26968 -7878 27086 -7866
rect 27202 -7469 27320 -7457
rect 27202 -7866 27208 -7469
rect 27314 -7866 27320 -7469
rect 27202 -7878 27320 -7866
rect 27436 -7469 27554 -7457
rect 27436 -7866 27442 -7469
rect 27548 -7866 27554 -7469
rect 27436 -7878 27554 -7866
rect 27670 -7469 27788 -7457
rect 27670 -7866 27676 -7469
rect 27782 -7866 27788 -7469
rect 27670 -7878 27788 -7866
rect 27904 -7469 28022 -7457
rect 27904 -7866 27910 -7469
rect 28016 -7866 28022 -7469
rect 27904 -7878 28022 -7866
rect 28138 -7469 28256 -7457
rect 28138 -7866 28144 -7469
rect 28250 -7866 28256 -7469
rect 28138 -7878 28256 -7866
rect 28372 -7469 28490 -7457
rect 28372 -7866 28378 -7469
rect 28484 -7866 28490 -7469
rect 28372 -7878 28490 -7866
rect 28606 -7469 28724 -7457
rect 28606 -7866 28612 -7469
rect 28718 -7866 28724 -7469
rect 28606 -7878 28724 -7866
rect 28840 -7469 28958 -7457
rect 28840 -7866 28846 -7469
rect 28952 -7866 28958 -7469
rect 28840 -7878 28958 -7866
rect 29074 -7469 29192 -7457
rect 29074 -7866 29080 -7469
rect 29186 -7866 29192 -7469
rect 29074 -7878 29192 -7866
rect 29308 -7469 29426 -7457
rect 29308 -7866 29314 -7469
rect 29420 -7866 29426 -7469
rect 29308 -7878 29426 -7866
rect 29542 -7469 29660 -7457
rect 29542 -7866 29548 -7469
rect 29654 -7866 29660 -7469
rect 29542 -7878 29660 -7866
rect 29776 -7469 29894 -7457
rect 29776 -7866 29782 -7469
rect 29888 -7866 29894 -7469
rect 29776 -7878 29894 -7866
<< properties >>
string FIXED_BBOX -30017 -7997 30017 7997
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 35.0 m 2 nx 256 wmin 0.690 lmin 0.50 class resistor rho 319.8 val 16.786k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
