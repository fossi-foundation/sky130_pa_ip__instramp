magic
tech sky130A
magscale 1 2
timestamp 1729620069
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use sky130_fd_pr__nfet_g5v0d10v5_92HZNS  XM1
timestamp 1729620069
transform 1 0 728 0 1 -534
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_TUFYNQ  XM2
timestamp 1729620069
transform 1 0 730 0 1 -1459
box -308 -397 308 397
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 UPPER
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 PGATE
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 NGATE
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 LOWER
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 DVSS
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 DVDD
port 5 nsew
<< end >>
