magic
tech sky130A
magscale 1 2
timestamp 1729620069
<< nwell >>
rect -1282 -2219 1282 2219
<< pmoslvt >>
rect -1086 -2000 -86 2000
rect 86 -2000 1086 2000
<< pdiff >>
rect -1144 1988 -1086 2000
rect -1144 -1988 -1132 1988
rect -1098 -1988 -1086 1988
rect -1144 -2000 -1086 -1988
rect -86 1988 -28 2000
rect -86 -1988 -74 1988
rect -40 -1988 -28 1988
rect -86 -2000 -28 -1988
rect 28 1988 86 2000
rect 28 -1988 40 1988
rect 74 -1988 86 1988
rect 28 -2000 86 -1988
rect 1086 1988 1144 2000
rect 1086 -1988 1098 1988
rect 1132 -1988 1144 1988
rect 1086 -2000 1144 -1988
<< pdiffc >>
rect -1132 -1988 -1098 1988
rect -74 -1988 -40 1988
rect 40 -1988 74 1988
rect 1098 -1988 1132 1988
<< nsubdiff >>
rect -1246 2149 -1150 2183
rect 1150 2149 1246 2183
rect -1246 2087 -1212 2149
rect 1212 2087 1246 2149
rect -1246 -2149 -1212 -2087
rect 1212 -2149 1246 -2087
rect -1246 -2183 -1150 -2149
rect 1150 -2183 1246 -2149
<< nsubdiffcont >>
rect -1150 2149 1150 2183
rect -1246 -2087 -1212 2087
rect 1212 -2087 1246 2087
rect -1150 -2183 1150 -2149
<< poly >>
rect -1086 2081 -86 2097
rect -1086 2047 -1070 2081
rect -102 2047 -86 2081
rect -1086 2000 -86 2047
rect 86 2081 1086 2097
rect 86 2047 102 2081
rect 1070 2047 1086 2081
rect 86 2000 1086 2047
rect -1086 -2047 -86 -2000
rect -1086 -2081 -1070 -2047
rect -102 -2081 -86 -2047
rect -1086 -2097 -86 -2081
rect 86 -2047 1086 -2000
rect 86 -2081 102 -2047
rect 1070 -2081 1086 -2047
rect 86 -2097 1086 -2081
<< polycont >>
rect -1070 2047 -102 2081
rect 102 2047 1070 2081
rect -1070 -2081 -102 -2047
rect 102 -2081 1070 -2047
<< locali >>
rect -1246 2149 -1150 2183
rect 1150 2149 1246 2183
rect -1246 2087 -1212 2149
rect 1212 2087 1246 2149
rect -1086 2047 -1070 2081
rect -102 2047 -86 2081
rect 86 2047 102 2081
rect 1070 2047 1086 2081
rect -1132 1988 -1098 2004
rect -1132 -2004 -1098 -1988
rect -74 1988 -40 2004
rect -74 -2004 -40 -1988
rect 40 1988 74 2004
rect 40 -2004 74 -1988
rect 1098 1988 1132 2004
rect 1098 -2004 1132 -1988
rect -1086 -2081 -1070 -2047
rect -102 -2081 -86 -2047
rect 86 -2081 102 -2047
rect 1070 -2081 1086 -2047
rect -1246 -2149 -1212 -2087
rect 1212 -2149 1246 -2087
rect -1246 -2183 -1150 -2149
rect 1150 -2183 1246 -2149
<< viali >>
rect -1070 2047 -102 2081
rect 102 2047 1070 2081
rect -1132 -1988 -1098 1988
rect -74 -1988 -40 1988
rect 40 -1988 74 1988
rect 1098 -1988 1132 1988
rect -1070 -2081 -102 -2047
rect 102 -2081 1070 -2047
<< metal1 >>
rect -1082 2081 -90 2087
rect -1082 2047 -1070 2081
rect -102 2047 -90 2081
rect -1082 2041 -90 2047
rect 90 2081 1082 2087
rect 90 2047 102 2081
rect 1070 2047 1082 2081
rect 90 2041 1082 2047
rect -1138 1988 -1092 2000
rect -1138 -1988 -1132 1988
rect -1098 -1988 -1092 1988
rect -1138 -2000 -1092 -1988
rect -80 1988 -34 2000
rect -80 -1988 -74 1988
rect -40 -1988 -34 1988
rect -80 -2000 -34 -1988
rect 34 1988 80 2000
rect 34 -1988 40 1988
rect 74 -1988 80 1988
rect 34 -2000 80 -1988
rect 1092 1988 1138 2000
rect 1092 -1988 1098 1988
rect 1132 -1988 1138 1988
rect 1092 -2000 1138 -1988
rect -1082 -2047 -90 -2041
rect -1082 -2081 -1070 -2047
rect -102 -2081 -90 -2047
rect -1082 -2087 -90 -2081
rect 90 -2047 1082 -2041
rect 90 -2081 102 -2047
rect 1070 -2081 1082 -2047
rect 90 -2087 1082 -2081
<< properties >>
string FIXED_BBOX -1229 -2166 1229 2166
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 20.0 l 5.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.35 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
