magic
tech sky130A
timestamp 1729620069
<< pwell >>
rect -1067 -379 1067 379
<< mvnmos >>
rect -953 -250 -853 250
rect -824 -250 -724 250
rect -695 -250 -595 250
rect -566 -250 -466 250
rect -437 -250 -337 250
rect -308 -250 -208 250
rect -179 -250 -79 250
rect -50 -250 50 250
rect 79 -250 179 250
rect 208 -250 308 250
rect 337 -250 437 250
rect 466 -250 566 250
rect 595 -250 695 250
rect 724 -250 824 250
rect 853 -250 953 250
<< mvndiff >>
rect -982 244 -953 250
rect -982 -244 -976 244
rect -959 -244 -953 244
rect -982 -250 -953 -244
rect -853 244 -824 250
rect -853 -244 -847 244
rect -830 -244 -824 244
rect -853 -250 -824 -244
rect -724 244 -695 250
rect -724 -244 -718 244
rect -701 -244 -695 244
rect -724 -250 -695 -244
rect -595 244 -566 250
rect -595 -244 -589 244
rect -572 -244 -566 244
rect -595 -250 -566 -244
rect -466 244 -437 250
rect -466 -244 -460 244
rect -443 -244 -437 244
rect -466 -250 -437 -244
rect -337 244 -308 250
rect -337 -244 -331 244
rect -314 -244 -308 244
rect -337 -250 -308 -244
rect -208 244 -179 250
rect -208 -244 -202 244
rect -185 -244 -179 244
rect -208 -250 -179 -244
rect -79 244 -50 250
rect -79 -244 -73 244
rect -56 -244 -50 244
rect -79 -250 -50 -244
rect 50 244 79 250
rect 50 -244 56 244
rect 73 -244 79 244
rect 50 -250 79 -244
rect 179 244 208 250
rect 179 -244 185 244
rect 202 -244 208 244
rect 179 -250 208 -244
rect 308 244 337 250
rect 308 -244 314 244
rect 331 -244 337 244
rect 308 -250 337 -244
rect 437 244 466 250
rect 437 -244 443 244
rect 460 -244 466 244
rect 437 -250 466 -244
rect 566 244 595 250
rect 566 -244 572 244
rect 589 -244 595 244
rect 566 -250 595 -244
rect 695 244 724 250
rect 695 -244 701 244
rect 718 -244 724 244
rect 695 -250 724 -244
rect 824 244 853 250
rect 824 -244 830 244
rect 847 -244 853 244
rect 824 -250 853 -244
rect 953 244 982 250
rect 953 -244 959 244
rect 976 -244 982 244
rect 953 -250 982 -244
<< mvndiffc >>
rect -976 -244 -959 244
rect -847 -244 -830 244
rect -718 -244 -701 244
rect -589 -244 -572 244
rect -460 -244 -443 244
rect -331 -244 -314 244
rect -202 -244 -185 244
rect -73 -244 -56 244
rect 56 -244 73 244
rect 185 -244 202 244
rect 314 -244 331 244
rect 443 -244 460 244
rect 572 -244 589 244
rect 701 -244 718 244
rect 830 -244 847 244
rect 959 -244 976 244
<< mvpsubdiff >>
rect -1049 355 1049 361
rect -1049 338 -995 355
rect 995 338 1049 355
rect -1049 332 1049 338
rect -1049 307 -1020 332
rect -1049 -307 -1043 307
rect -1026 -307 -1020 307
rect 1020 307 1049 332
rect -1049 -332 -1020 -307
rect 1020 -307 1026 307
rect 1043 -307 1049 307
rect 1020 -332 1049 -307
rect -1049 -338 1049 -332
rect -1049 -355 -995 -338
rect 995 -355 1049 -338
rect -1049 -361 1049 -355
<< mvpsubdiffcont >>
rect -995 338 995 355
rect -1043 -307 -1026 307
rect 1026 -307 1043 307
rect -995 -355 995 -338
<< poly >>
rect -953 286 -853 294
rect -953 269 -945 286
rect -861 269 -853 286
rect -953 250 -853 269
rect -824 286 -724 294
rect -824 269 -816 286
rect -732 269 -724 286
rect -824 250 -724 269
rect -695 286 -595 294
rect -695 269 -687 286
rect -603 269 -595 286
rect -695 250 -595 269
rect -566 286 -466 294
rect -566 269 -558 286
rect -474 269 -466 286
rect -566 250 -466 269
rect -437 286 -337 294
rect -437 269 -429 286
rect -345 269 -337 286
rect -437 250 -337 269
rect -308 286 -208 294
rect -308 269 -300 286
rect -216 269 -208 286
rect -308 250 -208 269
rect -179 286 -79 294
rect -179 269 -171 286
rect -87 269 -79 286
rect -179 250 -79 269
rect -50 286 50 294
rect -50 269 -42 286
rect 42 269 50 286
rect -50 250 50 269
rect 79 286 179 294
rect 79 269 87 286
rect 171 269 179 286
rect 79 250 179 269
rect 208 286 308 294
rect 208 269 216 286
rect 300 269 308 286
rect 208 250 308 269
rect 337 286 437 294
rect 337 269 345 286
rect 429 269 437 286
rect 337 250 437 269
rect 466 286 566 294
rect 466 269 474 286
rect 558 269 566 286
rect 466 250 566 269
rect 595 286 695 294
rect 595 269 603 286
rect 687 269 695 286
rect 595 250 695 269
rect 724 286 824 294
rect 724 269 732 286
rect 816 269 824 286
rect 724 250 824 269
rect 853 286 953 294
rect 853 269 861 286
rect 945 269 953 286
rect 853 250 953 269
rect -953 -269 -853 -250
rect -953 -286 -945 -269
rect -861 -286 -853 -269
rect -953 -294 -853 -286
rect -824 -269 -724 -250
rect -824 -286 -816 -269
rect -732 -286 -724 -269
rect -824 -294 -724 -286
rect -695 -269 -595 -250
rect -695 -286 -687 -269
rect -603 -286 -595 -269
rect -695 -294 -595 -286
rect -566 -269 -466 -250
rect -566 -286 -558 -269
rect -474 -286 -466 -269
rect -566 -294 -466 -286
rect -437 -269 -337 -250
rect -437 -286 -429 -269
rect -345 -286 -337 -269
rect -437 -294 -337 -286
rect -308 -269 -208 -250
rect -308 -286 -300 -269
rect -216 -286 -208 -269
rect -308 -294 -208 -286
rect -179 -269 -79 -250
rect -179 -286 -171 -269
rect -87 -286 -79 -269
rect -179 -294 -79 -286
rect -50 -269 50 -250
rect -50 -286 -42 -269
rect 42 -286 50 -269
rect -50 -294 50 -286
rect 79 -269 179 -250
rect 79 -286 87 -269
rect 171 -286 179 -269
rect 79 -294 179 -286
rect 208 -269 308 -250
rect 208 -286 216 -269
rect 300 -286 308 -269
rect 208 -294 308 -286
rect 337 -269 437 -250
rect 337 -286 345 -269
rect 429 -286 437 -269
rect 337 -294 437 -286
rect 466 -269 566 -250
rect 466 -286 474 -269
rect 558 -286 566 -269
rect 466 -294 566 -286
rect 595 -269 695 -250
rect 595 -286 603 -269
rect 687 -286 695 -269
rect 595 -294 695 -286
rect 724 -269 824 -250
rect 724 -286 732 -269
rect 816 -286 824 -269
rect 724 -294 824 -286
rect 853 -269 953 -250
rect 853 -286 861 -269
rect 945 -286 953 -269
rect 853 -294 953 -286
<< polycont >>
rect -945 269 -861 286
rect -816 269 -732 286
rect -687 269 -603 286
rect -558 269 -474 286
rect -429 269 -345 286
rect -300 269 -216 286
rect -171 269 -87 286
rect -42 269 42 286
rect 87 269 171 286
rect 216 269 300 286
rect 345 269 429 286
rect 474 269 558 286
rect 603 269 687 286
rect 732 269 816 286
rect 861 269 945 286
rect -945 -286 -861 -269
rect -816 -286 -732 -269
rect -687 -286 -603 -269
rect -558 -286 -474 -269
rect -429 -286 -345 -269
rect -300 -286 -216 -269
rect -171 -286 -87 -269
rect -42 -286 42 -269
rect 87 -286 171 -269
rect 216 -286 300 -269
rect 345 -286 429 -269
rect 474 -286 558 -269
rect 603 -286 687 -269
rect 732 -286 816 -269
rect 861 -286 945 -269
<< locali >>
rect -1043 338 -995 355
rect 995 338 1043 355
rect -1043 307 -1026 338
rect 1026 307 1043 338
rect -953 269 -945 286
rect -861 269 -853 286
rect -824 269 -816 286
rect -732 269 -724 286
rect -695 269 -687 286
rect -603 269 -595 286
rect -566 269 -558 286
rect -474 269 -466 286
rect -437 269 -429 286
rect -345 269 -337 286
rect -308 269 -300 286
rect -216 269 -208 286
rect -179 269 -171 286
rect -87 269 -79 286
rect -50 269 -42 286
rect 42 269 50 286
rect 79 269 87 286
rect 171 269 179 286
rect 208 269 216 286
rect 300 269 308 286
rect 337 269 345 286
rect 429 269 437 286
rect 466 269 474 286
rect 558 269 566 286
rect 595 269 603 286
rect 687 269 695 286
rect 724 269 732 286
rect 816 269 824 286
rect 853 269 861 286
rect 945 269 953 286
rect -976 244 -959 252
rect -976 -252 -959 -244
rect -847 244 -830 252
rect -847 -252 -830 -244
rect -718 244 -701 252
rect -718 -252 -701 -244
rect -589 244 -572 252
rect -589 -252 -572 -244
rect -460 244 -443 252
rect -460 -252 -443 -244
rect -331 244 -314 252
rect -331 -252 -314 -244
rect -202 244 -185 252
rect -202 -252 -185 -244
rect -73 244 -56 252
rect -73 -252 -56 -244
rect 56 244 73 252
rect 56 -252 73 -244
rect 185 244 202 252
rect 185 -252 202 -244
rect 314 244 331 252
rect 314 -252 331 -244
rect 443 244 460 252
rect 443 -252 460 -244
rect 572 244 589 252
rect 572 -252 589 -244
rect 701 244 718 252
rect 701 -252 718 -244
rect 830 244 847 252
rect 830 -252 847 -244
rect 959 244 976 252
rect 959 -252 976 -244
rect -953 -286 -945 -269
rect -861 -286 -853 -269
rect -824 -286 -816 -269
rect -732 -286 -724 -269
rect -695 -286 -687 -269
rect -603 -286 -595 -269
rect -566 -286 -558 -269
rect -474 -286 -466 -269
rect -437 -286 -429 -269
rect -345 -286 -337 -269
rect -308 -286 -300 -269
rect -216 -286 -208 -269
rect -179 -286 -171 -269
rect -87 -286 -79 -269
rect -50 -286 -42 -269
rect 42 -286 50 -269
rect 79 -286 87 -269
rect 171 -286 179 -269
rect 208 -286 216 -269
rect 300 -286 308 -269
rect 337 -286 345 -269
rect 429 -286 437 -269
rect 466 -286 474 -269
rect 558 -286 566 -269
rect 595 -286 603 -269
rect 687 -286 695 -269
rect 724 -286 732 -269
rect 816 -286 824 -269
rect 853 -286 861 -269
rect 945 -286 953 -269
rect -1043 -338 -1026 -307
rect 1026 -338 1043 -307
rect -1043 -355 -995 -338
rect 995 -355 1043 -338
<< viali >>
rect -945 269 -861 286
rect -816 269 -732 286
rect -687 269 -603 286
rect -558 269 -474 286
rect -429 269 -345 286
rect -300 269 -216 286
rect -171 269 -87 286
rect -42 269 42 286
rect 87 269 171 286
rect 216 269 300 286
rect 345 269 429 286
rect 474 269 558 286
rect 603 269 687 286
rect 732 269 816 286
rect 861 269 945 286
rect -976 -244 -959 244
rect -847 -244 -830 244
rect -718 -244 -701 244
rect -589 -244 -572 244
rect -460 -244 -443 244
rect -331 -244 -314 244
rect -202 -244 -185 244
rect -73 -244 -56 244
rect 56 -244 73 244
rect 185 -244 202 244
rect 314 -244 331 244
rect 443 -244 460 244
rect 572 -244 589 244
rect 701 -244 718 244
rect 830 -244 847 244
rect 959 -244 976 244
rect -945 -286 -861 -269
rect -816 -286 -732 -269
rect -687 -286 -603 -269
rect -558 -286 -474 -269
rect -429 -286 -345 -269
rect -300 -286 -216 -269
rect -171 -286 -87 -269
rect -42 -286 42 -269
rect 87 -286 171 -269
rect 216 -286 300 -269
rect 345 -286 429 -269
rect 474 -286 558 -269
rect 603 -286 687 -269
rect 732 -286 816 -269
rect 861 -286 945 -269
<< metal1 >>
rect -951 286 -855 289
rect -951 269 -945 286
rect -861 269 -855 286
rect -951 266 -855 269
rect -822 286 -726 289
rect -822 269 -816 286
rect -732 269 -726 286
rect -822 266 -726 269
rect -693 286 -597 289
rect -693 269 -687 286
rect -603 269 -597 286
rect -693 266 -597 269
rect -564 286 -468 289
rect -564 269 -558 286
rect -474 269 -468 286
rect -564 266 -468 269
rect -435 286 -339 289
rect -435 269 -429 286
rect -345 269 -339 286
rect -435 266 -339 269
rect -306 286 -210 289
rect -306 269 -300 286
rect -216 269 -210 286
rect -306 266 -210 269
rect -177 286 -81 289
rect -177 269 -171 286
rect -87 269 -81 286
rect -177 266 -81 269
rect -48 286 48 289
rect -48 269 -42 286
rect 42 269 48 286
rect -48 266 48 269
rect 81 286 177 289
rect 81 269 87 286
rect 171 269 177 286
rect 81 266 177 269
rect 210 286 306 289
rect 210 269 216 286
rect 300 269 306 286
rect 210 266 306 269
rect 339 286 435 289
rect 339 269 345 286
rect 429 269 435 286
rect 339 266 435 269
rect 468 286 564 289
rect 468 269 474 286
rect 558 269 564 286
rect 468 266 564 269
rect 597 286 693 289
rect 597 269 603 286
rect 687 269 693 286
rect 597 266 693 269
rect 726 286 822 289
rect 726 269 732 286
rect 816 269 822 286
rect 726 266 822 269
rect 855 286 951 289
rect 855 269 861 286
rect 945 269 951 286
rect 855 266 951 269
rect -979 244 -956 250
rect -979 -244 -976 244
rect -959 -244 -956 244
rect -979 -250 -956 -244
rect -850 244 -827 250
rect -850 -244 -847 244
rect -830 -244 -827 244
rect -850 -250 -827 -244
rect -721 244 -698 250
rect -721 -244 -718 244
rect -701 -244 -698 244
rect -721 -250 -698 -244
rect -592 244 -569 250
rect -592 -244 -589 244
rect -572 -244 -569 244
rect -592 -250 -569 -244
rect -463 244 -440 250
rect -463 -244 -460 244
rect -443 -244 -440 244
rect -463 -250 -440 -244
rect -334 244 -311 250
rect -334 -244 -331 244
rect -314 -244 -311 244
rect -334 -250 -311 -244
rect -205 244 -182 250
rect -205 -244 -202 244
rect -185 -244 -182 244
rect -205 -250 -182 -244
rect -76 244 -53 250
rect -76 -244 -73 244
rect -56 -244 -53 244
rect -76 -250 -53 -244
rect 53 244 76 250
rect 53 -244 56 244
rect 73 -244 76 244
rect 53 -250 76 -244
rect 182 244 205 250
rect 182 -244 185 244
rect 202 -244 205 244
rect 182 -250 205 -244
rect 311 244 334 250
rect 311 -244 314 244
rect 331 -244 334 244
rect 311 -250 334 -244
rect 440 244 463 250
rect 440 -244 443 244
rect 460 -244 463 244
rect 440 -250 463 -244
rect 569 244 592 250
rect 569 -244 572 244
rect 589 -244 592 244
rect 569 -250 592 -244
rect 698 244 721 250
rect 698 -244 701 244
rect 718 -244 721 244
rect 698 -250 721 -244
rect 827 244 850 250
rect 827 -244 830 244
rect 847 -244 850 244
rect 827 -250 850 -244
rect 956 244 979 250
rect 956 -244 959 244
rect 976 -244 979 244
rect 956 -250 979 -244
rect -951 -269 -855 -266
rect -951 -286 -945 -269
rect -861 -286 -855 -269
rect -951 -289 -855 -286
rect -822 -269 -726 -266
rect -822 -286 -816 -269
rect -732 -286 -726 -269
rect -822 -289 -726 -286
rect -693 -269 -597 -266
rect -693 -286 -687 -269
rect -603 -286 -597 -269
rect -693 -289 -597 -286
rect -564 -269 -468 -266
rect -564 -286 -558 -269
rect -474 -286 -468 -269
rect -564 -289 -468 -286
rect -435 -269 -339 -266
rect -435 -286 -429 -269
rect -345 -286 -339 -269
rect -435 -289 -339 -286
rect -306 -269 -210 -266
rect -306 -286 -300 -269
rect -216 -286 -210 -269
rect -306 -289 -210 -286
rect -177 -269 -81 -266
rect -177 -286 -171 -269
rect -87 -286 -81 -269
rect -177 -289 -81 -286
rect -48 -269 48 -266
rect -48 -286 -42 -269
rect 42 -286 48 -269
rect -48 -289 48 -286
rect 81 -269 177 -266
rect 81 -286 87 -269
rect 171 -286 177 -269
rect 81 -289 177 -286
rect 210 -269 306 -266
rect 210 -286 216 -269
rect 300 -286 306 -269
rect 210 -289 306 -286
rect 339 -269 435 -266
rect 339 -286 345 -269
rect 429 -286 435 -269
rect 339 -289 435 -286
rect 468 -269 564 -266
rect 468 -286 474 -269
rect 558 -286 564 -269
rect 468 -289 564 -286
rect 597 -269 693 -266
rect 597 -286 603 -269
rect 687 -286 693 -269
rect 597 -289 693 -286
rect 726 -269 822 -266
rect 726 -286 732 -269
rect 816 -286 822 -269
rect 726 -289 822 -286
rect 855 -269 951 -266
rect 855 -286 861 -269
rect 945 -286 951 -269
rect 855 -289 951 -286
<< properties >>
string FIXED_BBOX -1034 -346 1034 346
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 1.0 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
