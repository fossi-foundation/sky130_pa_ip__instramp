* NGSPICE file created from sky130_pa_ip__instramp.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__lsbuflv2hv_1 A LVPWR VGND VNB VPB VPWR X VPWR_uq0 VGND_uq0
+ VNB_uq0
X0 VGND a_404_1133# a_504_1221# VNB_uq0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1 a_504_1221# a_404_1133# VGND VNB_uq0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2 X a_1711_885# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
R0 VNB_uq0 VNB 0.000000
X3 X a_1711_885# VGND VNB_uq0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X4 VGND_uq0 A a_404_1133# VNB_uq0 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X5 a_1197_107# a_772_151# VGND_uq0 VNB_uq0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X6 VPWR_uq0 a_1197_107# a_504_1221# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X7 a_504_1221# a_404_1133# VGND VNB_uq0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X8 a_1197_107# a_772_151# VGND_uq0 VNB_uq0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X9 a_504_1221# a_404_1133# VGND VNB_uq0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X10 VGND a_404_1133# a_504_1221# VNB_uq0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X11 a_772_151# a_404_1133# VGND_uq0 VNB_uq0 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X12 VGND_uq0 a_772_151# a_1197_107# VNB_uq0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X13 LVPWR A a_404_1133# LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X14 VPWR a_504_1221# a_1711_885# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X15 VGND a_504_1221# a_1711_885# VNB_uq0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X16 VGND_uq0 a_772_151# a_1197_107# VNB_uq0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X17 a_772_151# a_404_1133# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X18 a_1197_107# a_772_151# VGND_uq0 VNB_uq0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X19 VPWR a_504_1221# a_1197_107# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
.ends

.subckt sky130_fd_sc_hvl__inv_1 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP a_214_n1416# a_n118_984# a_48_n1416#
+ a_n450_984# a_n580_n1546# a_n284_n1416# a_n118_n1416# a_48_984# a_380_984# a_380_n1416#
+ a_214_984# a_n284_984# a_n450_n1416#
X0 a_n118_984# a_n118_n1416# a_n580_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X1 a_380_984# a_380_n1416# a_n580_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X2 a_214_984# a_214_n1416# a_n580_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X3 a_n284_984# a_n284_n1416# a_n580_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X4 a_n450_984# a_n450_n1416# a_n580_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X5 a_48_984# a_48_n1416# a_n580_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
.ends

.subckt sky130_fd_sc_hvl__diode_2 DIODE VGND VNB VPB VPWR
X0 VNB DIODE sky130_fd_pr__diode_pw2nd_11v0 perim=3.16e+06 area=6.072e+11
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_92HZNS a_50_n100# a_n242_n322# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n242_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_TUFYNQ a_n50_n197# a_50_n100# w_n308_n397# a_n108_n100#
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n308_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt T_Gate_5V UPPER PGATE NGATE LOWER AVSS AVDD
XXM1 LOWER AVSS UPPER NGATE sky130_fd_pr__nfet_g5v0d10v5_92HZNS
XXM2 PGATE LOWER AVDD UPPER sky130_fd_pr__pfet_g5v0d10v5_TUFYNQ
.ends

.subckt Universal_R_2R_Block2 VD DVDD CMOUT R2RIN R2ROUT VIRTOUT AVSS DVSS AVDD
Xx1 VD DVDD DVSS DVSS AVDD AVDD VDbuf AVDD DVSS DVSS sky130_fd_sc_hvl__lsbuflv2hv_1
Xx2 VDbuf DVSS DVSS AVDD AVDD VDBAR sky130_fd_sc_hvl__inv_1
Xsky130_fd_pr__res_xhigh_po_0p35_Q2LWZP_0 m1_4390_n2466# m1_6792_n1970# m1_4394_n2136#
+ x13/LOWER AVSS m1_4392_n1802# m1_4394_n2136# R2ROUT R2RIN m1_4390_n2466# R2ROUT
+ m1_6792_n1970# m1_4392_n1802# sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP
Xsky130_fd_sc_hvl__diode_2_0 VD DVSS DVSS AVDD AVDD sky130_fd_sc_hvl__diode_2
Xx12 VIRTOUT VDBAR VDbuf x13/LOWER AVSS AVDD T_Gate_5V
Xx13 CMOUT VDbuf VDBAR x13/LOWER AVSS AVDD T_Gate_5V
.ends

.subckt sky130_fd_pr__res_high_po_0p69_FJD3D2 a_n199_n4646# a_n69_4084# a_n69_n4516#
X0 a_n69_4084# a_n69_n4516# a_n199_n4646# sky130_fd_pr__res_high_po_0p69 l=41
.ends

.subckt sky130_fd_pr__nfet_05v0_nvt_FEJX3A a_952_n991# a_n1352_n573# a_200_318# a_318_736#
+ a_n952_n518# a_n258_n100# a_n952_736# a_776_n100# a_n834_318# a_n776_n991# a_n258_n936#
+ a_n258_736# a_952_681# a_776_n936# a_894_736# a_n834_n518# a_n200_n573# a_318_n100#
+ a_776_318# a_200_n518# a_n1352_681# a_376_n991# a_1352_n518# a_318_n936# a_n376_n518#
+ a_894_n518# a_318_318# a_n1544_n1158# a_952_n573# a_n1352_n155# a_n952_318# a_n1410_n100#
+ a_n1410_736# a_n376_736# a_n200_681# a_n1410_n936# a_n258_n518# a_n776_n573# a_n258_318#
+ a_776_n518# a_894_318# a_952_263# a_n200_n155# a_1352_736# a_376_681# a_n1352_263#
+ a_318_n518# a_376_n573# a_n776_681# a_n952_n100# a_952_n155# a_200_736# a_n952_n936#
+ a_n1352_n991# a_n1410_318# a_n376_318# a_n200_263# a_n776_n155# a_n834_736# a_n1410_n518#
+ a_n834_n100# a_200_n100# a_1352_318# a_n200_n991# a_1352_n100# a_376_263# a_n834_n936#
+ a_n376_n100# a_776_736# a_1352_n936# a_200_n936# a_894_n100# a_376_n155# a_n376_n936#
+ a_n776_263# a_894_n936#
X0 a_1352_n518# a_952_n573# a_894_n518# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X1 a_n376_n518# a_n776_n573# a_n834_n518# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X2 a_n952_n100# a_n1352_n155# a_n1410_n100# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X3 a_n376_n100# a_n776_n155# a_n834_n100# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X4 a_200_n100# a_n200_n155# a_n258_n100# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X5 a_776_736# a_376_681# a_318_736# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X6 a_1352_736# a_952_681# a_894_736# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X7 a_n952_n518# a_n1352_n573# a_n1410_n518# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X8 a_n952_318# a_n1352_263# a_n1410_318# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X9 a_776_n936# a_376_n991# a_318_n936# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X10 a_200_n936# a_n200_n991# a_n258_n936# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X11 a_n376_318# a_n776_263# a_n834_318# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X12 a_200_318# a_n200_263# a_n258_318# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X13 a_776_n100# a_376_n155# a_318_n100# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X14 a_1352_n100# a_952_n155# a_894_n100# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X15 a_n376_n936# a_n776_n991# a_n834_n936# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X16 a_1352_n936# a_952_n991# a_894_n936# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X17 a_776_318# a_376_263# a_318_318# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X18 a_1352_318# a_952_263# a_894_318# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X19 a_n952_n936# a_n1352_n991# a_n1410_n936# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X20 a_n952_736# a_n1352_681# a_n1410_736# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X21 a_200_736# a_n200_681# a_n258_736# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X22 a_776_n518# a_376_n573# a_318_n518# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X23 a_n376_736# a_n776_681# a_n834_736# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X24 a_200_n518# a_n200_n573# a_n258_n518# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_NZU856 a_616_n1610# a_n2938_n2808# a_n2738_n500#
+ a_874_n2720# a_n1190_n1610# a_1132_1720# a_n1448_610# a_n932_610# a_n416_n1610#
+ a_1390_n1610# a_1906_n500# a_n674_n2720# a_1132_n2720# a_n2480_n500# a_n2996_1720#
+ a_n2164_n2808# a_n416_610# a_n2738_n1610# a_n2996_n2720# a_1390_610# a_2938_n1610#
+ a_n1648_n2808# a_358_n500# a_n158_1720# a_2222_n2808# a_2164_n500# a_874_610# a_1706_n2808#
+ a_n1706_n500# a_2164_n1610# a_674_n2808# a_n674_n500# a_100_n500# a_n1448_n1610#
+ a_358_610# a_616_1720# a_1648_n1610# a_n1964_1720# a_2422_1720# a_n100_n2808# a_n932_n2720#
+ a_n1190_610# a_358_n2720# a_n932_1720# a_1132_n500# a_100_n1610# a_n158_n2720# a_n2422_n2808#
+ a_1648_1720# a_n674_610# a_n1906_n2808# a_n2996_n500# a_1390_1720# a_n158_610# a_n2222_1720#
+ a_n2222_n1610# a_n2480_n2720# a_n158_n500# a_2422_n1610# a_2680_n2720# a_932_n2808#
+ a_n1132_n2808# a_n1706_n1610# a_n874_n2808# a_n1964_n2720# a_n1448_1720# a_1906_n1610#
+ a_158_n2808# a_874_n1610# a_616_n2720# a_n1190_1720# a_616_n500# a_n674_n1610# a_n1190_n2720#
+ a_n416_1720# a_2938_610# a_2422_610# a_n1964_n500# a_1132_n1610# a_1390_n2720# a_n416_n2720#
+ a_1906_610# a_2422_n500# a_2938_1720# a_n2996_n1610# a_874_1720# a_n2738_n2720#
+ a_n932_n500# a_2938_n2720# a_2480_n2808# a_2680_1720# a_1648_n500# a_1964_n2808#
+ a_n2222_n500# a_1390_n500# a_n2738_1720# a_2164_n2720# a_416_n2808# a_n358_n2808#
+ a_n2738_610# a_n1448_n2720# a_n2222_610# a_n1706_610# a_1648_n2720# a_1906_1720#
+ a_1190_n2808# a_n2480_1720# a_n1448_n500# a_n932_n1610# a_358_n1610# a_2680_610#
+ a_n2680_n2808# a_n158_n1610# a_358_1720# a_n1190_n500# a_2738_n2808# a_2164_610#
+ a_100_n2720# a_n416_n500# a_1648_610# a_2164_1720# a_1132_610# a_n1706_1720# a_2938_n500#
+ a_874_n500# a_n2480_n1610# a_100_1720# a_n674_1720# a_2680_n1610# a_n2222_n2720#
+ a_n1390_n2808# a_100_610# a_616_610# a_n1964_n1610# a_2680_n500# a_1448_n2808# a_2422_n2720#
+ a_n616_n2808# a_n3130_n2942# a_n1706_n2720# a_n2996_610# a_n2480_610# a_1906_n2720#
+ a_n1964_610#
X0 a_n2480_n2720# a_n2680_n2808# a_n2738_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X1 a_n1448_n1610# a_n1648_n2808# a_n1706_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X2 a_2938_n2720# a_2738_n2808# a_2680_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X3 a_1906_n1610# a_1706_n2808# a_1648_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X4 a_1906_n500# a_1706_n2808# a_1648_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X5 a_1648_n500# a_1448_n2808# a_1390_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X6 a_1906_1720# a_1706_n2808# a_1648_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X7 a_n1190_n2720# a_n1390_n2808# a_n1448_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X8 a_1648_1720# a_1448_n2808# a_1390_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X9 a_2938_610# a_2738_n2808# a_2680_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X10 a_n674_610# a_n874_n2808# a_n932_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X11 a_1648_n2720# a_1448_n2808# a_1390_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X12 a_n1448_610# a_n1648_n2808# a_n1706_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X13 a_n1964_610# a_n2164_n2808# a_n2222_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X14 a_874_n1610# a_674_n2808# a_616_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X15 a_2680_n1610# a_2480_n2808# a_2422_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X16 a_1132_n500# a_932_n2808# a_874_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X17 a_1132_1720# a_932_n2808# a_874_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X18 a_n1964_n1610# a_n2164_n2808# a_n2222_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X19 a_874_n500# a_674_n2808# a_616_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X20 a_1390_610# a_1190_n2808# a_1132_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X21 a_616_n1610# a_416_n2808# a_358_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X22 a_874_1720# a_674_n2808# a_616_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X23 a_2422_n1610# a_2222_n2808# a_2164_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X24 a_1390_n1610# a_1190_n2808# a_1132_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X25 a_n2738_610# a_n2938_n2808# a_n2996_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X26 a_358_n2720# a_158_n2808# a_100_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X27 a_n674_n1610# a_n874_n2808# a_n932_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X28 a_2164_610# a_1964_n2808# a_1906_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X29 a_2164_n500# a_1964_n2808# a_1906_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X30 a_2680_610# a_2480_n2808# a_2422_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X31 a_n416_n1610# a_n616_n2808# a_n674_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X32 a_616_610# a_416_n2808# a_358_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X33 a_2164_1720# a_1964_n2808# a_1906_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X34 a_n2738_n500# a_n2938_n2808# a_n2996_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X35 a_100_n2720# a_n100_n2808# a_n158_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X36 a_n2738_n2720# a_n2938_n2808# a_n2996_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X37 a_n1706_n1610# a_n1906_n2808# a_n1964_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X38 a_n2738_1720# a_n2938_n2808# a_n2996_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X39 a_n158_n2720# a_n358_n2808# a_n416_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X40 a_n2480_n500# a_n2680_n2808# a_n2738_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X41 a_n1190_610# a_n1390_n2808# a_n1448_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X42 a_1390_n500# a_1190_n2808# a_1132_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X43 a_n2480_1720# a_n2680_n2808# a_n2738_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X44 a_2164_n2720# a_1964_n2808# a_1906_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X45 a_n2222_n500# a_n2422_n2808# a_n2480_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X46 a_1390_1720# a_1190_n2808# a_1132_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X47 a_n1448_n2720# a_n1648_n2808# a_n1706_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X48 a_n2222_1720# a_n2422_n2808# a_n2480_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X49 a_n1964_n500# a_n2164_n2808# a_n2222_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X50 a_1906_n2720# a_1706_n2808# a_1648_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X51 a_n1964_1720# a_n2164_n2808# a_n2222_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X52 a_1132_n1610# a_932_n2808# a_874_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X53 a_n2480_610# a_n2680_n2808# a_n2738_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X54 a_n2222_n1610# a_n2422_n2808# a_n2480_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X55 a_100_n500# a_n100_n2808# a_n158_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X56 a_874_n2720# a_674_n2808# a_616_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X57 a_100_1720# a_n100_n2808# a_n158_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X58 a_2680_n2720# a_2480_n2808# a_2422_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X59 a_n1964_n2720# a_n2164_n2808# a_n2222_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X60 a_n932_n1610# a_n1132_n2808# a_n1190_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X61 a_358_610# a_158_n2808# a_100_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X62 a_616_n2720# a_416_n2808# a_358_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X63 a_2422_n2720# a_2222_n2808# a_2164_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X64 a_1390_n2720# a_1190_n2808# a_1132_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X65 a_2938_n500# a_2738_n2808# a_2680_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X66 a_1132_610# a_932_n2808# a_874_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X67 a_2938_1720# a_2738_n2808# a_2680_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X68 a_n416_610# a_n616_n2808# a_n674_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X69 a_n674_n2720# a_n874_n2808# a_n932_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X70 a_2422_n500# a_2222_n2808# a_2164_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X71 a_n416_n500# a_n616_n2808# a_n674_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X72 a_2422_1720# a_2222_n2808# a_2164_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X73 a_n416_n2720# a_n616_n2808# a_n674_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X74 a_n158_n500# a_n358_n2808# a_n416_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X75 a_n416_1720# a_n616_n2808# a_n674_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X76 a_n158_1720# a_n358_n2808# a_n416_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X77 a_n1706_n2720# a_n1906_n2808# a_n1964_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X78 a_n2480_n1610# a_n2680_n2808# a_n2738_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X79 a_2938_n1610# a_2738_n2808# a_2680_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X80 a_n1190_n1610# a_n1390_n2808# a_n1448_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X81 a_1906_610# a_1706_n2808# a_1648_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X82 a_1648_n1610# a_1448_n2808# a_1390_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X83 a_2422_610# a_2222_n2808# a_2164_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X84 a_1132_n2720# a_932_n2808# a_874_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X85 a_n932_610# a_n1132_n2808# a_n1190_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X86 a_874_610# a_674_n2808# a_616_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X87 a_n1706_n500# a_n1906_n2808# a_n1964_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X88 a_n158_610# a_n358_n2808# a_n416_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X89 a_n2222_n2720# a_n2422_n2808# a_n2480_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X90 a_2680_n500# a_2480_n2808# a_2422_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X91 a_n1706_1720# a_n1906_n2808# a_n1964_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X92 a_n1448_n500# a_n1648_n2808# a_n1706_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X93 a_n674_n500# a_n874_n2808# a_n932_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X94 a_n1190_n500# a_n1390_n2808# a_n1448_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X95 a_n1448_1720# a_n1648_n2808# a_n1706_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X96 a_2680_1720# a_2480_n2808# a_2422_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X97 a_n674_1720# a_n874_n2808# a_n932_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X98 a_n932_n2720# a_n1132_n2808# a_n1190_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X99 a_n1190_1720# a_n1390_n2808# a_n1448_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X100 a_100_610# a_n100_n2808# a_n158_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X101 a_n1706_610# a_n1906_n2808# a_n1964_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X102 a_358_n1610# a_158_n2808# a_100_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X103 a_n932_n500# a_n1132_n2808# a_n1190_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X104 a_n932_1720# a_n1132_n2808# a_n1190_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X105 a_n2222_610# a_n2422_n2808# a_n2480_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X106 a_616_n500# a_416_n2808# a_358_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X107 a_616_1720# a_416_n2808# a_358_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X108 a_358_n500# a_158_n2808# a_100_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X109 a_100_n1610# a_n100_n2808# a_n158_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X110 a_n2738_n1610# a_n2938_n2808# a_n2996_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X111 a_1648_610# a_1448_n2808# a_1390_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X112 a_358_1720# a_158_n2808# a_100_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X113 a_n158_n1610# a_n358_n2808# a_n416_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X114 a_2164_n1610# a_1964_n2808# a_1906_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_AJ3MPE a_72_772# a_n90_n750# a_n138_n838# a_n182_n750#
+ a_n284_n924# a_120_n750# a_28_n750#
X0 a_120_n750# a_72_772# a_28_n750# a_n284_n924# sky130_fd_pr__nfet_01v8_lvt ad=2.325 pd=15.62 as=2.325 ps=15.62 w=7.5 l=0.15
X1 a_n90_n750# a_n138_n838# a_n182_n750# a_n284_n924# sky130_fd_pr__nfet_01v8_lvt ad=2.325 pd=15.62 as=2.325 ps=15.62 w=7.5 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_UX3DP3 a_n1087_n4118# a_29_n4215# a_1029_118#
+ a_n29_n4118# a_29_21# a_n1029_21# w_n1225_n4337# a_n1087_118# a_1029_n4118# a_n1029_n4215#
+ a_n29_118#
X0 a_n29_n4118# a_n1029_n4215# a_n1087_n4118# w_n1225_n4337# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=5.8 ps=40.58 w=20 l=5
X1 a_1029_n4118# a_29_n4215# a_n29_n4118# w_n1225_n4337# sky130_fd_pr__pfet_01v8_lvt ad=5.8 pd=40.58 as=2.9 ps=20.29 w=20 l=5
X2 a_1029_118# a_29_21# a_n29_118# w_n1225_n4337# sky130_fd_pr__pfet_01v8_lvt ad=5.8 pd=40.58 as=2.9 ps=20.29 w=20 l=5
X3 a_n29_118# a_n1029_21# a_n1087_118# w_n1225_n4337# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=5.8 ps=40.58 w=20 l=5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_8UL4MK a_467_n1000# a_n803_n1000# w_n1559_n1297#
+ a_1301_n1000# a_n645_n1000# a_1143_n1000# a_189_n1000# a_n525_n1000# a_923_n1097#
+ a_1023_n1000# a_n1201_n1000# a_n367_n1000# a_n1359_n1000# a_n745_n1097# a_n89_n1000#
+ a_n247_n1000# a_645_n1097# a_865_n1000# a_n467_n1097# a_n1301_n1097# a_745_n1000#
+ a_n1081_n1000# a_367_n1097# a_89_n1097# a_587_n1000# a_309_n1000# a_31_n1000# a_n923_n1000#
+ a_1201_n1097# a_n189_n1097# a_n1023_n1097#
X0 a_n1201_n1000# a_n1301_n1097# a_n1359_n1000# w_n1559_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.5
X1 a_1301_n1000# a_1201_n1097# a_1143_n1000# w_n1559_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.5
X2 a_189_n1000# a_89_n1097# a_31_n1000# w_n1559_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.5
X3 a_n645_n1000# a_n745_n1097# a_n803_n1000# w_n1559_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.5
X4 a_745_n1000# a_645_n1097# a_587_n1000# w_n1559_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.5
X5 a_n89_n1000# a_n189_n1097# a_n247_n1000# w_n1559_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.5
X6 a_n923_n1000# a_n1023_n1097# a_n1081_n1000# w_n1559_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.5
X7 a_1023_n1000# a_923_n1097# a_865_n1000# w_n1559_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.5
X8 a_n367_n1000# a_n467_n1097# a_n525_n1000# w_n1559_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.5
X9 a_467_n1000# a_367_n1097# a_309_n1000# w_n1559_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.5
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_BHK9HY c1_n3758_n5640# c1_1466_n5640# m3_1426_n5680#
+ m3_n1186_n5680# m3_n3798_n5680# c1_n1146_n5640#
X0 c1_n3758_n5640# m3_n3798_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X1 c1_n1146_n5640# m3_n1186_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X2 c1_1466_n5640# m3_1426_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X3 c1_n3758_n5640# m3_n3798_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X4 c1_1466_n5640# m3_1426_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X5 c1_n3758_n5640# m3_n3798_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X6 c1_n1146_n5640# m3_n1186_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X7 c1_n3758_n5640# m3_n3798_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X8 c1_n1146_n5640# m3_n1186_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X9 c1_1466_n5640# m3_1426_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X10 c1_1466_n5640# m3_1426_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X11 c1_1466_n5640# m3_1426_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X12 c1_n1146_n5640# m3_n1186_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X13 c1_n3758_n5640# m3_n3798_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X14 c1_n1146_n5640# m3_n1186_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
.ends

.subckt x1_x32_OA VDD VOUT VINN VINP VBIAS w_8718_n902# w_7736_n902# VSS w_4240_n902#
XXR1 VSS m1_10706_1822# VOUT sky130_fd_pr__res_high_po_0p69_FJD3D2
Xsky130_fd_pr__nfet_05v0_nvt_FEJX3A_0 VINP VINP w_8718_n902# w_8718_n902# w_8718_n902#
+ m1_9368_n744# w_8718_n902# m1_9368_n744# w_8718_n902# VINP m1_9368_n744# m1_9368_n744#
+ VINP m1_9368_n744# m1_9368_n744# w_8718_n902# VINP w_8718_n902# m1_9368_n744# w_8718_n902#
+ VINP VINP w_8718_n902# w_8718_n902# m1_9368_n744# m1_9368_n744# w_8718_n902# w_8718_n902#
+ VINP VINP w_8718_n902# m1_9368_n744# m1_9368_n744# m1_9368_n744# VINP m1_9368_n744#
+ m1_9368_n744# VINP m1_9368_n744# m1_9368_n744# m1_9368_n744# VINP VINP w_8718_n902#
+ VINP VINP w_8718_n902# VINP VINP w_8718_n902# VINP w_8718_n902# w_8718_n902# VINP
+ m1_9368_n744# m1_9368_n744# VINP VINP w_8718_n902# m1_9368_n744# w_8718_n902# w_8718_n902#
+ w_8718_n902# VINP w_8718_n902# VINP w_8718_n902# m1_9368_n744# m1_9368_n744# w_8718_n902#
+ w_8718_n902# m1_9368_n744# VINP m1_9368_n744# VINP m1_9368_n744# sky130_fd_pr__nfet_05v0_nvt_FEJX3A
Xsky130_fd_pr__nfet_g5v0d10v5_NZU856_0 VSS VBIAS VOUT VOUT VOUT VSS VSS VSS VSS VOUT
+ VOUT VOUT VSS VSS VSS VBIAS VSS VOUT VSS VOUT w_7736_n902# VBIAS VOUT VOUT VBIAS
+ VSS VOUT VBIAS VOUT VSS VBIAS VOUT VSS VSS VOUT VSS VSS VSS w_7736_n902# VBIAS VSS
+ VOUT VOUT VSS VSS VSS VOUT VBIAS VSS VOUT VBIAS VSS VOUT VOUT VOUT VOUT VSS VOUT
+ w_7736_n902# VSS VBIAS VBIAS VOUT VBIAS VSS VSS VOUT VBIAS VOUT VSS VOUT VSS VOUT
+ VOUT VSS w_7736_n902# w_7736_n902# VSS VSS VOUT VSS VOUT w_7736_n902# w_7736_n902#
+ VSS VOUT VOUT VSS w_7736_n902# VBIAS VSS VSS VBIAS VOUT VOUT VOUT VSS VBIAS VBIAS
+ VOUT VSS VOUT VOUT VSS VOUT VBIAS VSS VSS VSS VOUT VSS VBIAS VOUT VOUT VOUT VBIAS
+ VSS VSS VSS VSS VSS VSS VOUT w_7736_n902# VOUT VSS VSS VOUT VSS VOUT VBIAS VSS VSS
+ VSS VSS VBIAS w_7736_n902# VBIAS VSS VOUT VSS VSS VOUT VSS sky130_fd_pr__nfet_g5v0d10v5_NZU856
XXM2 VINN w_8718_n902# VINP w_7736_n902# w_7736_n902# w_4240_n902# w_7736_n902# sky130_fd_pr__nfet_01v8_lvt_AJ3MPE
XXM6 m1_9368_n744# m1_4902_n766# m1_9368_n744# VDD m1_4902_n766# m1_4902_n766# VDD
+ m1_4902_n766# m1_4902_n766# m1_4902_n766# VDD sky130_fd_pr__pfet_01v8_lvt_UX3DP3
XXM8 VDD VOUT VDD VOUT VDD VDD VOUT VDD m1_9368_n744# VDD VDD VOUT VOUT m1_9368_n744#
+ VDD VOUT m1_9368_n744# VOUT m1_9368_n744# m1_9368_n744# VOUT VDD m1_9368_n744# m1_9368_n744#
+ VDD VOUT VDD VOUT m1_9368_n744# m1_9368_n744# m1_9368_n744# sky130_fd_pr__pfet_g5v0d10v5_8UL4MK
Xsky130_fd_pr__cap_mim_m3_1_BHK9HY_0 m1_9368_n744# m1_9368_n744# m1_10706_1822# m1_10706_1822#
+ m1_10706_1822# m1_9368_n744# sky130_fd_pr__cap_mim_m3_1_BHK9HY
XXM10 VINN VINN m1_4902_n766# m1_4902_n766# m1_4902_n766# w_4240_n902# m1_4902_n766#
+ w_4240_n902# m1_4902_n766# VINN w_4240_n902# w_4240_n902# VINN w_4240_n902# w_4240_n902#
+ m1_4902_n766# VINN m1_4902_n766# w_4240_n902# m1_4902_n766# VINN VINN m1_4902_n766#
+ m1_4902_n766# w_4240_n902# w_4240_n902# m1_4902_n766# w_4240_n902# VINN VINN m1_4902_n766#
+ w_4240_n902# w_4240_n902# w_4240_n902# VINN w_4240_n902# w_4240_n902# VINN w_4240_n902#
+ w_4240_n902# w_4240_n902# VINN VINN m1_4902_n766# VINN VINN m1_4902_n766# VINN VINN
+ m1_4902_n766# VINN m1_4902_n766# m1_4902_n766# VINN w_4240_n902# w_4240_n902# VINN
+ VINN m1_4902_n766# w_4240_n902# m1_4902_n766# m1_4902_n766# m1_4902_n766# VINN m1_4902_n766#
+ VINN m1_4902_n766# w_4240_n902# w_4240_n902# m1_4902_n766# m1_4902_n766# w_4240_n902#
+ VINN w_4240_n902# VINN w_4240_n902# sky130_fd_pr__nfet_05v0_nvt_FEJX3A
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_3WU84W a_n3899_n1610# a_n29_n2720# a_3067_1720#
+ a_4357_n2720# a_1261_n500# a_n287_610# a_n4673_610# a_487_n1610# a_1777_1720# a_n2609_1720#
+ a_4873_1720# a_n803_n2720# a_n3641_610# a_n5705_1720# a_n5389_n2808# a_229_n2720#
+ a_3383_n2808# a_n5189_610# a_n287_n1610# a_n3641_n2720# a_n4157_610# a_2867_n2808#
+ a_3841_n2720# a_n2351_1720# a_n1319_n500# a_5389_1720# a_3583_n500# a_n3125_610#
+ a_5447_n2808# a_n4415_n500# a_n5705_n2720# a_n2609_610# a_n4873_n2808# a_3067_n2720#
+ a_n287_n500# a_229_1720# a_n5189_n1610# a_n1061_n500# a_4099_n500# a_3583_610# a_n1577_1720#
+ a_5389_n1610# a_n4099_n2808# a_n4673_1720# a_4931_n2808# a_2093_n2808# a_2551_610#
+ a_2035_1720# a_n2351_n2720# a_4099_610# a_5131_1720# a_1577_n2808# a_2551_n2720#
+ a_803_n2808# a_n745_n2808# a_n1003_n2808# a_n4673_n1610# a_n1835_n2720# a_2809_n500#
+ a_3067_610# a_3841_1720# a_4157_n2808# a_5131_n2720# a_745_n500# a_n5189_1720# a_4873_n1610#
+ a_n4415_n2720# a_n3383_n500# a_2035_610# a_n545_1720# a_n3899_1720# a_n3583_n2808#
+ a_4615_n2720# a_1519_610# a_1003_610# a_745_n1610# a_4357_1720# a_2551_n500# a_4099_n1610#
+ a_3641_n2808# a_n5647_n2808# a_n1061_n2720# a_n545_n1610# a_1003_n1610# a_1261_n2720#
+ a_n3383_n1610# a_3067_n500# a_1777_n500# a_n3899_610# a_n3641_1720# a_3583_n1610#
+ a_n2609_n500# a_n3383_610# a_1003_1720# a_n2293_n2808# a_4873_n500# a_n2867_n1610#
+ a_n3125_n2720# a_n5705_n500# a_n2351_610# a_n2867_610# a_3325_n2720# a_n5447_n1610#
+ a_n2609_n2720# a_n1835_610# a_n1777_n2808# a_5647_n1610# a_n4157_1720# a_n4357_n2808#
+ a_2809_n2720# a_n2351_n500# a_2351_n2808# a_5389_n500# a_n2867_1720# a_n1319_610#
+ a_3325_1720# a_1835_n2808# a_n803_610# a_n4931_n1610# a_n2093_n1610# a_229_n500#
+ a_4415_n2808# a_2293_n1610# a_n3841_n2808# a_n1577_n1610# a_n1577_n500# a_n5705_610#
+ a_n4673_n500# a_2293_610# a_2035_n2720# a_n229_n2808# a_n4157_n1610# a_n29_n1610#
+ a_1777_n1610# a_n1319_n2720# a_2035_n500# a_1777_610# a_1261_610# a_n29_1720# a_5131_n500#
+ a_4357_n1610# a_1519_n2720# a_5647_1720# a_487_1720# a_n3067_n2808# a_3841_n500#
+ a_1061_n2808# a_n3899_n2720# a_n803_n1610# a_n5189_n500# a_229_n1610# a_n545_n500#
+ a_487_n2720# a_n3899_n500# a_n3641_n1610# a_2293_1720# a_n3125_1720# a_745_610#
+ a_3125_n2808# a_4357_n500# a_n1835_1720# a_3841_n1610# a_n4931_1720# a_n2551_n2808#
+ a_n287_n2720# a_5647_610# a_5131_610# a_2609_n2808# a_4615_610# a_n5131_n2808# a_n5705_n1610#
+ a_229_610# a_3067_n1610# a_n4615_n2808# a_n5447_1720# a_n3641_n500# a_n803_1720#
+ a_n5189_n2720# a_1003_n500# a_n2093_610# a_1519_1720# a_n2351_n1610# a_5389_n2720#
+ a_n1577_610# a_4615_1720# a_n1061_610# a_n2093_1720# a_2551_n1610# a_n4157_n500#
+ a_n1261_n2808# a_n1835_n1610# a_1319_n2808# a_5131_n1610# a_n2867_n500# a_n4415_n1610#
+ a_1261_1720# a_n4673_n2720# a_n545_610# a_3325_n500# a_n4931_610# a_3899_n2808#
+ a_4615_n1610# a_4873_n2720# a_287_n2808# a_n3325_n2808# a_n5447_610# a_n2809_n2808#
+ a_745_n2720# a_n1061_n1610# a_4099_n2720# a_n4415_610# a_n1319_1720# a_n29_n500#
+ a_3583_1720# a_n4415_1720# a_1261_n1610# a_5647_n500# a_n545_n2720# a_487_n500#
+ a_1003_n2720# a_n287_1720# a_n3125_n1610# a_n3383_n2720# a_4873_610# a_n1061_1720#
+ a_4099_1720# a_3325_n1610# a_3583_n2720# a_2293_n500# a_n3125_n500# a_487_610# a_n2035_n2808#
+ a_n2609_n1610# a_n2867_n2720# a_3841_610# a_5189_n2808# a_n1835_n500# a_2809_n1610#
+ a_n4931_n500# a_5389_610# a_n1519_n2808# a_n5447_n2720# a_4357_610# a_5647_n2720#
+ a_2809_1720# a_n29_610# a_3325_610# a_745_1720# a_n3383_1720# a_n5447_n500# a_2809_610#
+ a_4673_n2808# a_n5839_n2942# a_n4931_n2720# a_n2093_n2720# a_n803_n500# a_2551_1720#
+ a_2035_n1610# a_1519_n500# a_545_n2808# a_4615_n500# a_n1319_n1610# a_2293_n2720#
+ a_29_n2808# a_n487_n2808# a_n1577_n2720# a_n2093_n500# a_1519_n1610# a_n4157_n2720#
+ a_1777_n2720#
X0 a_5389_n2720# a_5189_n2808# a_5131_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X1 a_4357_n1610# a_4157_n2808# a_4099_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X2 a_n1061_1720# a_n1261_n2808# a_n1319_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X3 a_2551_n2720# a_2351_n2808# a_2293_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X4 a_n803_610# a_n1003_n2808# a_n1061_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X5 a_1003_n500# a_803_n2808# a_745_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X6 a_n1835_n2720# a_n2035_n2808# a_n2093_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X7 a_n803_n1610# a_n1003_n2808# a_n1061_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X8 a_745_610# a_545_n2808# a_487_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X9 a_1003_1720# a_803_n2808# a_745_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X10 a_5389_610# a_5189_n2808# a_5131_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X11 a_745_n500# a_545_n2808# a_487_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X12 a_n29_610# a_n229_n2808# a_n287_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X13 a_n3899_610# a_n4099_n2808# a_n4157_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X14 a_1261_n2720# a_1061_n2808# a_1003_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X15 a_745_1720# a_545_n2808# a_487_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X16 a_487_n500# a_287_n2808# a_229_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X17 a_n4931_n2720# a_n5131_n2808# a_n5189_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X18 a_487_1720# a_287_n2808# a_229_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X19 a_n4673_610# a_n4873_n2808# a_n4931_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X20 a_229_n2720# a_29_n2808# a_n29_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X21 a_n545_n2720# a_n745_n2808# a_n803_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X22 a_229_610# a_29_n2808# a_n29_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X23 a_2035_n500# a_1835_n2808# a_1777_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X24 a_4099_n500# a_3899_n2808# a_3841_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X25 a_4099_n2720# a_3899_n2808# a_3841_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X26 a_3067_n1610# a_2867_n2808# a_2809_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X27 a_2035_1720# a_1835_n2808# a_1777_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X28 a_4099_1720# a_3899_n2808# a_3841_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X29 a_n5189_610# a_n5389_n2808# a_n5447_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X30 a_1777_n500# a_1577_n2808# a_1519_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X31 a_4099_610# a_3899_n2808# a_3841_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X32 a_n2609_n500# a_n2809_n2808# a_n2867_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X33 a_3841_n500# a_3641_n2808# a_3583_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X34 a_1777_1720# a_1577_n2808# a_1519_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X35 a_n2609_1720# a_n2809_n2808# a_n2867_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X36 a_3841_1720# a_3641_n2808# a_3583_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X37 a_1519_610# a_1319_n2808# a_1261_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X38 a_3583_n500# a_3383_n2808# a_3325_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X39 a_2809_n1610# a_2609_n2808# a_2551_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X40 a_n4415_n500# a_n4615_n2808# a_n4673_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X41 a_1261_n500# a_1061_n2808# a_1003_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X42 a_1777_n1610# a_1577_n2808# a_1519_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X43 a_n5447_n1610# a_n5647_n2808# a_n5705_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X44 a_3583_1720# a_3383_n2808# a_3325_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X45 a_n3641_n2720# a_n3841_n2808# a_n3899_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X46 a_n4415_1720# a_n4615_n2808# a_n4673_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X47 a_n4157_n500# a_n4357_n2808# a_n4415_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X48 a_1261_1720# a_1061_n2808# a_1003_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X49 a_n3899_n500# a_n4099_n2808# a_n4157_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X50 a_n1835_n500# a_n2035_n2808# a_n2093_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X51 a_n4157_1720# a_n4357_n2808# a_n4415_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X52 a_4873_n1610# a_4673_n2808# a_4615_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X53 a_1519_n1610# a_1319_n2808# a_1261_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X54 a_487_610# a_287_n2808# a_229_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X55 a_n3899_1720# a_n4099_n2808# a_n4157_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X56 a_n1835_1720# a_n2035_n2808# a_n2093_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X57 a_n5189_n2720# a_n5389_n2808# a_n5447_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X58 a_n4157_n1610# a_n4357_n2808# a_n4415_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X59 a_n2351_n2720# a_n2551_n2808# a_n2609_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X60 a_1003_n2720# a_803_n2808# a_745_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X61 a_5647_n2720# a_5447_n2808# a_5389_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X62 a_4615_n1610# a_4415_n2808# a_4357_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X63 a_3583_n1610# a_3383_n2808# a_3325_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X64 a_n545_610# a_n745_n2808# a_n803_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X65 a_2809_610# a_2609_n2808# a_2551_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X66 a_n3899_n2720# a_n4099_n2808# a_n4157_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X67 a_n2867_n1610# a_n3067_n2808# a_n3125_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X68 a_n1319_610# a_n1519_n2808# a_n1577_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X69 a_n1061_n2720# a_n1261_n2808# a_n1319_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X70 a_4357_n2720# a_4157_n2808# a_4099_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X71 a_487_n1610# a_287_n2808# a_229_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X72 a_3325_610# a_3125_n2808# a_3067_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X73 a_3325_n1610# a_3125_n2808# a_3067_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X74 a_2293_n1610# a_2093_n2808# a_2035_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X75 a_n1835_610# a_n2035_n2808# a_n2093_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X76 a_n803_n2720# a_n1003_n2808# a_n1061_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X77 a_1261_610# a_1061_n2808# a_1003_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X78 a_2809_n500# a_2609_n2808# a_2551_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X79 a_n4673_n500# a_n4873_n2808# a_n4931_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X80 a_2809_1720# a_2609_n2808# a_2551_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X81 a_n2609_610# a_n2809_n2808# a_n2867_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X82 a_n287_n1610# a_n487_n2808# a_n545_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X83 a_4615_n500# a_4415_n2808# a_4357_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X84 a_n4673_1720# a_n4873_n2808# a_n4931_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X85 a_4615_610# a_4415_n2808# a_4357_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X86 a_n2351_n500# a_n2551_n2808# a_n2609_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X87 a_4357_n500# a_4157_n2808# a_4099_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X88 a_4615_1720# a_4415_n2808# a_4357_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X89 a_n3125_610# a_n3325_n2808# a_n3383_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X90 a_n2609_n1610# a_n2809_n2808# a_n2867_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X91 a_n2351_1720# a_n2551_n2808# a_n2609_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X92 a_2035_610# a_1835_n2808# a_1777_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X93 a_n2093_n500# a_n2293_n2808# a_n2351_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X94 a_4357_1720# a_4157_n2808# a_4099_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X95 a_229_n500# a_29_n2808# a_n29_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X96 a_n29_n1610# a_n229_n2808# a_n287_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X97 a_n1577_n1610# a_n1777_n2808# a_n1835_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X98 a_n2093_1720# a_n2293_n2808# a_n2351_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X99 a_n29_n500# a_n229_n2808# a_n287_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X100 a_229_1720# a_29_n2808# a_n29_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X101 a_2551_610# a_2351_n2808# a_2293_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X102 a_3067_n2720# a_2867_n2808# a_2809_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X103 a_2035_n1610# a_1835_n2808# a_1777_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X104 a_n29_1720# a_n229_n2808# a_n287_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X105 a_n1061_610# a_n1261_n2808# a_n1319_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X106 a_n1319_n1610# a_n1519_n2808# a_n1577_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X107 a_n4673_n1610# a_n4873_n2808# a_n4931_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X108 a_n287_610# a_n487_n2808# a_n545_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X109 a_2809_n2720# a_2609_n2808# a_2551_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X110 a_5131_n1610# a_4931_n2808# a_4873_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X111 a_1777_n2720# a_1577_n2808# a_1519_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X112 a_n5447_n2720# a_n5647_n2808# a_n5705_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X113 a_n4415_n1610# a_n4615_n2808# a_n4673_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X114 a_n3383_n1610# a_n3583_n2808# a_n3641_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X115 a_n4415_610# a_n4615_n2808# a_n4673_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X116 a_4873_n2720# a_4673_n2808# a_4615_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X117 a_3841_n1610# a_3641_n2808# a_3583_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X118 a_1519_n2720# a_1319_n2808# a_1261_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X119 a_n4931_610# a_n5131_n2808# a_n5189_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X120 a_3841_610# a_3641_n2808# a_3583_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X121 a_n4157_n2720# a_n4357_n2808# a_n4415_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X122 a_n3125_n1610# a_n3325_n2808# a_n3383_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X123 a_n2093_n1610# a_n2293_n2808# a_n2351_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X124 a_n2351_610# a_n2551_n2808# a_n2609_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X125 a_745_n1610# a_545_n2808# a_487_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X126 a_3067_n500# a_2867_n2808# a_2809_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X127 a_4615_n2720# a_4415_n2808# a_4357_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X128 a_5389_n1610# a_5189_n2808# a_5131_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X129 a_3583_n2720# a_3383_n2808# a_3325_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X130 a_2551_n1610# a_2351_n2808# a_2293_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X131 a_5131_n500# a_4931_n2808# a_4873_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X132 a_3067_1720# a_2867_n2808# a_2809_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X133 a_n2867_n2720# a_n3067_n2808# a_n3125_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X134 a_n1835_n1610# a_n2035_n2808# a_n2093_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X135 a_5131_1720# a_4931_n2808# a_4873_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X136 a_4873_n500# a_4673_n2808# a_4615_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X137 a_4357_610# a_4157_n2808# a_4099_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X138 a_3325_n2720# a_3125_n2808# a_3067_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X139 a_487_n2720# a_287_n2808# a_229_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X140 a_4873_1720# a_4673_n2808# a_4615_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X141 a_n1319_n500# a_n1519_n2808# a_n1577_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X142 a_2551_n500# a_2351_n2808# a_2293_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X143 a_n2867_610# a_n3067_n2808# a_n3125_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X144 a_n5447_n500# a_n5647_n2808# a_n5705_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X145 a_2293_n2720# a_2093_n2808# a_2035_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X146 a_1261_n1610# a_1061_n2808# a_1003_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X147 a_n4931_n1610# a_n5131_n2808# a_n5189_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X148 a_1777_610# a_1577_n2808# a_1519_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X149 a_n545_n500# a_n745_n2808# a_n803_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X150 a_2293_n500# a_2093_n2808# a_2035_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X151 a_n1319_1720# a_n1519_n2808# a_n1577_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X152 a_2551_1720# a_2351_n2808# a_2293_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X153 a_n5189_n500# a_n5389_n2808# a_n5447_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X154 a_n5447_1720# a_n5647_n2808# a_n5705_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X155 a_n3125_n500# a_n3325_n2808# a_n3383_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X156 a_n287_n500# a_n487_n2808# a_n545_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X157 a_n545_1720# a_n745_n2808# a_n803_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X158 a_2293_1720# a_2093_n2808# a_2035_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X159 a_2293_610# a_2093_n2808# a_2035_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X160 a_5131_610# a_4931_n2808# a_4873_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X161 a_n2867_n500# a_n3067_n2808# a_n3125_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X162 a_n803_n500# a_n1003_n2808# a_n1061_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X163 a_229_n1610# a_29_n2808# a_n29_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X164 a_n545_n1610# a_n745_n2808# a_n803_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X165 a_n5189_1720# a_n5389_n2808# a_n5447_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X166 a_n3125_1720# a_n3325_n2808# a_n3383_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X167 a_n287_1720# a_n487_n2808# a_n545_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X168 a_n3641_610# a_n3841_n2808# a_n3899_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X169 a_n4931_n500# a_n5131_n2808# a_n5189_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X170 a_n2867_1720# a_n3067_n2808# a_n3125_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X171 a_n803_1720# a_n1003_n2808# a_n1061_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X172 a_n4931_1720# a_n5131_n2808# a_n5189_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X173 a_1003_610# a_803_n2808# a_745_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X174 a_n287_n2720# a_n487_n2808# a_n545_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X175 a_5647_610# a_5447_n2808# a_5389_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X176 a_4099_n1610# a_3899_n2808# a_3841_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X177 a_n4157_610# a_n4357_n2808# a_n4415_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X178 a_3067_610# a_2867_n2808# a_2809_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X179 a_n2609_n2720# a_n2809_n2808# a_n2867_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X180 a_n1577_610# a_n1777_n2808# a_n1835_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X181 a_n29_n2720# a_n229_n2808# a_n287_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X182 a_n1577_n2720# a_n1777_n2808# a_n1835_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X183 a_3583_610# a_3383_n2808# a_3325_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X184 a_2035_n2720# a_1835_n2808# a_1777_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X185 a_n2093_610# a_n2293_n2808# a_n2351_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X186 a_n4673_n2720# a_n4873_n2808# a_n4931_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X187 a_n1319_n2720# a_n1519_n2808# a_n1577_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X188 a_n3641_n1610# a_n3841_n2808# a_n3899_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X189 a_5131_n2720# a_4931_n2808# a_4873_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X190 a_n4415_n2720# a_n4615_n2808# a_n4673_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X191 a_n5189_n1610# a_n5389_n2808# a_n5447_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X192 a_n1577_n500# a_n1777_n2808# a_n1835_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X193 a_n3383_n2720# a_n3583_n2808# a_n3641_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X194 a_n2351_n1610# a_n2551_n2808# a_n2609_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X195 a_n5447_610# a_n5647_n2808# a_n5705_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X196 a_n3641_n500# a_n3841_n2808# a_n3899_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X197 a_1003_n1610# a_803_n2808# a_745_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X198 a_1519_n500# a_1319_n2808# a_1261_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X199 a_5647_n1610# a_5447_n2808# a_5389_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X200 a_5647_n500# a_5447_n2808# a_5389_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X201 a_3841_n2720# a_3641_n2808# a_3583_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X202 a_n1577_1720# a_n1777_n2808# a_n1835_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X203 a_n3383_n500# a_n3583_n2808# a_n3641_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X204 a_n3641_1720# a_n3841_n2808# a_n3899_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X205 a_1519_1720# a_1319_n2808# a_1261_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X206 a_3325_n500# a_3125_n2808# a_3067_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X207 a_n3125_n2720# a_n3325_n2808# a_n3383_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X208 a_5389_n500# a_5189_n2808# a_5131_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X209 a_5647_1720# a_5447_n2808# a_5389_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X210 a_4873_610# a_4673_n2808# a_4615_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X211 a_n3899_n1610# a_n4099_n2808# a_n4157_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X212 a_n3383_1720# a_n3583_n2808# a_n3641_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X213 a_n1061_n500# a_n1261_n2808# a_n1319_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X214 a_n2093_n2720# a_n2293_n2808# a_n2351_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X215 a_n1061_n1610# a_n1261_n2808# a_n1319_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X216 a_3325_1720# a_3125_n2808# a_3067_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X217 a_5389_1720# a_5189_n2808# a_5131_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X218 a_n3383_610# a_n3583_n2808# a_n3641_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X219 a_745_n2720# a_545_n2808# a_487_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
.ends

.subckt Output_OA VDD VOUT VINN VINP VBIAS w_8718_n902# w_7736_n902# VSS w_4240_n902#
XXR1 VSS m1_10706_1822# VOUT sky130_fd_pr__res_high_po_0p69_FJD3D2
Xsky130_fd_pr__nfet_05v0_nvt_FEJX3A_0 VINP VINP w_8718_n902# w_8718_n902# w_8718_n902#
+ m1_9368_n744# w_8718_n902# m1_9368_n744# w_8718_n902# VINP m1_9368_n744# m1_9368_n744#
+ VINP m1_9368_n744# m1_9368_n744# w_8718_n902# VINP w_8718_n902# m1_9368_n744# w_8718_n902#
+ VINP VINP w_8718_n902# w_8718_n902# m1_9368_n744# m1_9368_n744# w_8718_n902# w_8718_n902#
+ VINP VINP w_8718_n902# m1_9368_n744# m1_9368_n744# m1_9368_n744# VINP m1_9368_n744#
+ m1_9368_n744# VINP m1_9368_n744# m1_9368_n744# m1_9368_n744# VINP VINP w_8718_n902#
+ VINP VINP w_8718_n902# VINP VINP w_8718_n902# VINP w_8718_n902# w_8718_n902# VINP
+ m1_9368_n744# m1_9368_n744# VINP VINP w_8718_n902# m1_9368_n744# w_8718_n902# w_8718_n902#
+ w_8718_n902# VINP w_8718_n902# VINP w_8718_n902# m1_9368_n744# m1_9368_n744# w_8718_n902#
+ w_8718_n902# m1_9368_n744# VINP m1_9368_n744# VINP m1_9368_n744# sky130_fd_pr__nfet_05v0_nvt_FEJX3A
Xsky130_fd_pr__nfet_g5v0d10v5_3WU84W_0 VOUT VSS VSS VOUT VOUT VOUT VSS VSS VOUT VSS
+ w_7736_n902# VOUT VSS VSS VBIAS VOUT VBIAS VSS VOUT VSS VSS VBIAS VOUT VOUT VOUT
+ w_7736_n902# VSS VSS VBIAS VOUT VSS VSS VBIAS VSS VOUT VOUT VSS VSS VSS VSS VSS
+ w_7736_n902# VBIAS VSS VBIAS VBIAS VSS VSS VOUT VSS VSS VBIAS VSS VBIAS VBIAS VBIAS
+ VSS VOUT VOUT VSS VOUT VBIAS VSS VOUT VSS w_7736_n902# VOUT VOUT VSS VSS VOUT VBIAS
+ VSS VSS VSS VOUT VOUT VSS VSS VBIAS VBIAS VSS VSS VSS VOUT VOUT VSS VOUT VOUT VSS
+ VSS VSS VOUT VSS VBIAS w_7736_n902# VOUT VSS VSS VOUT VOUT VOUT VOUT VSS VOUT VBIAS
+ VSS VSS VBIAS VOUT VOUT VBIAS w_7736_n902# VOUT VOUT VOUT VBIAS VOUT VOUT VSS VOUT
+ VBIAS VOUT VBIAS VSS VSS VSS VSS VOUT VSS VBIAS VSS VSS VOUT VOUT VSS VOUT VOUT
+ VSS VSS VOUT VSS VSS VSS VBIAS VOUT VBIAS VOUT VOUT VSS VOUT VSS VSS VOUT VSS VOUT
+ VSS VOUT VBIAS VOUT VOUT VOUT VOUT VBIAS VOUT VSS VSS VBIAS VSS VBIAS VSS VOUT VSS
+ VBIAS VOUT VSS VOUT VSS VSS VSS VSS VOUT w_7736_n902# VSS VSS VSS VSS VSS VSS VBIAS
+ VOUT VBIAS VSS VOUT VOUT VOUT VSS VSS VOUT VOUT VBIAS VSS w_7736_n902# VBIAS VBIAS
+ VOUT VBIAS VOUT VSS VSS VOUT VOUT VSS VSS VOUT VOUT VSS VSS VSS VSS VOUT VSS VOUT
+ w_7736_n902# VSS VSS VOUT VSS VOUT VSS VSS VBIAS VSS VOUT VOUT VBIAS VOUT VOUT VOUT
+ w_7736_n902# VBIAS VOUT VOUT VSS VOUT VSS VOUT VOUT VOUT VOUT VOUT VBIAS VSS VOUT
+ VSS VOUT VSS VSS VSS VBIAS VSS VOUT VOUT VBIAS VBIAS VSS VSS VSS VSS VOUT sky130_fd_pr__nfet_g5v0d10v5_3WU84W
XXM2 VINN w_8718_n902# VINP w_7736_n902# w_7736_n902# w_4240_n902# w_7736_n902# sky130_fd_pr__nfet_01v8_lvt_AJ3MPE
XXM6 m1_9368_n744# m1_4902_n766# m1_9368_n744# VDD m1_4902_n766# m1_4902_n766# VDD
+ m1_4902_n766# m1_4902_n766# m1_4902_n766# VDD sky130_fd_pr__pfet_01v8_lvt_UX3DP3
XXM8 VDD VOUT VDD VOUT VDD VDD VOUT VDD m1_9368_n744# VDD VDD VOUT VOUT m1_9368_n744#
+ VDD VOUT m1_9368_n744# VOUT m1_9368_n744# m1_9368_n744# VOUT VDD m1_9368_n744# m1_9368_n744#
+ VDD VOUT VDD VOUT m1_9368_n744# m1_9368_n744# m1_9368_n744# sky130_fd_pr__pfet_g5v0d10v5_8UL4MK
Xsky130_fd_pr__cap_mim_m3_1_BHK9HY_0 m1_9368_n744# m1_9368_n744# m1_10706_1822# m1_10706_1822#
+ m1_10706_1822# m1_9368_n744# sky130_fd_pr__cap_mim_m3_1_BHK9HY
XXM10 VINN VINN m1_4902_n766# m1_4902_n766# m1_4902_n766# w_4240_n902# m1_4902_n766#
+ w_4240_n902# m1_4902_n766# VINN w_4240_n902# w_4240_n902# VINN w_4240_n902# w_4240_n902#
+ m1_4902_n766# VINN m1_4902_n766# w_4240_n902# m1_4902_n766# VINN VINN m1_4902_n766#
+ m1_4902_n766# w_4240_n902# w_4240_n902# m1_4902_n766# w_4240_n902# VINN VINN m1_4902_n766#
+ w_4240_n902# w_4240_n902# w_4240_n902# VINN w_4240_n902# w_4240_n902# VINN w_4240_n902#
+ w_4240_n902# w_4240_n902# VINN VINN m1_4902_n766# VINN VINN m1_4902_n766# VINN VINN
+ m1_4902_n766# VINN m1_4902_n766# m1_4902_n766# VINN w_4240_n902# w_4240_n902# VINN
+ VINN m1_4902_n766# w_4240_n902# m1_4902_n766# m1_4902_n766# m1_4902_n766# VINN m1_4902_n766#
+ VINN m1_4902_n766# w_4240_n902# w_4240_n902# m1_4902_n766# m1_4902_n766# w_4240_n902#
+ VINN w_4240_n902# VINN w_4240_n902# sky130_fd_pr__nfet_05v0_nvt_FEJX3A
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_V6AMGK a_n782_n1904# a_9178_n1904# a_13494_1472#
+ a_1376_n1904# a_2704_n1904# a_5194_1472# a_11336_n1904# a_8182_1472# a_6688_n1904#
+ a_n12900_1472# a_546_n1904# a_n10908_n1904# a_n3438_1472# a_10506_1472# a_n6426_1472#
+ a_n2110_1472# a_n12070_n1904# a_n9414_1472# a_n8750_n1904# a_2206_1472# a_12996_1472#
+ a_1708_n1904# a_n10244_1472# a_4696_1472# a_n13232_1472# a_7684_1472# a_48_1472#
+ a_n2442_n1904# a_8182_n1904# a_9510_n1904# a_n11074_n1904# a_n7754_n1904# a_n5928_1472#
+ a_n1612_1472# a_n12402_n1904# a_n4600_1472# a_n8916_1472# a_1708_1472# a_10340_n1904#
+ a_5692_n1904# a_n9248_n1904# a_3202_n1904# a_n12734_1472# a_n1446_n1904# a_n13896_n1904#
+ a_2870_1472# a_7186_n1904# a_8514_n1904# a_n10078_n1904# a_n6758_n1904# a_712_1472#
+ a_13328_1472# a_n11406_n1904# a_12000_1472# a_n9248_1472# a_n284_n1904# a_4696_n1904#
+ a_n948_1472# a_5028_1472# a_8016_1472# a_n10078_1472# a_2206_n1904# a_n13066_1472#
+ a_6190_1472# a_7518_n1904# a_n1446_1472# a_n4434_1472# a_11502_1472# a_n8252_n1904#
+ a_n616_n1904# a_n7422_1472# a_3202_1472# a_7518_1472# a_13992_1472# a_6190_n1904#
+ a_n12568_1472# a_n5762_n1904# a_n10410_n1904# a_n11240_1472# a_5692_1472# a_8680_1472#
+ a_546_1472# a_9012_n1904# a_n7256_n1904# a_13660_n1904# a_n3936_1472# a_1210_n1904#
+ a_n6924_1472# a_5194_n1904# a_n9912_1472# a_2704_1472# a_6522_n1904# a_n4766_n1904#
+ a_n10742_1472# a_n13398_n1904# a_n13730_1472# a_8016_n1904# a_12664_n1904# a_n4268_1472#
+ a_11336_1472# a_n7256_1472# a_4198_n1904# a_5526_n1904# a_3036_1472# a_14158_n1904#
+ a_6024_1472# a_9012_1472# a_n11074_1472# a_n6260_n1904# a_n14062_1472# a_11668_n1904#
+ a_878_n1904# a_10838_1472# a_n3770_n1904# a_n118_n1904# a_n6758_1472# a_n2442_1472#
+ a_13826_1472# a_n9746_1472# a_n5430_1472# a_2538_1472# a_n13730_n1904# a_1210_1472#
+ a_5526_1472# a_7020_n1904# a_n5264_n1904# a_8514_1472# a_n10576_1472# a_n13564_1472#
+ a_4530_n1904# a_n2774_n1904# a_14158_1472# a_13162_n1904# a_n1944_1472# a_9842_n1904#
+ a_n4932_1472# a_n12734_n1904# a_6024_n1904# a_n7920_1472# a_n4268_n1904# a_n450_1472#
+ a_10672_n1904# a_3700_1472# a_n14228_n1904# a_3534_n1904# a_n1778_n1904# a_12166_n1904#
+ a_n2276_1472# a_8846_n1904# a_12332_1472# a_n5264_1472# a_n11738_n1904# a_5028_n1904#
+ a_n8252_1472# a_1044_1472# a_4032_1472# a_8348_1472# a_n9580_n1904# a_7020_1472#
+ a_n13398_1472# a_2538_n1904# a_n12070_1472# a_n14358_n2034# a_n3272_n1904# a_n1778_1472#
+ a_n4766_1472# a_n4600_n1904# a_11834_1472# a_n7754_1472# a_n8584_n1904# a_n948_n1904#
+ a_n284_1472# a_n13232_n1904# a_n9912_n1904# a_3534_1472# a_11170_n1904# a_6522_1472#
+ a_380_n1904# a_7850_n1904# a_9510_1472# a_n11572_1472# a_n10742_n1904# a_4032_n1904#
+ a_n2276_n1904# a_878_1472# a_n5098_1472# a_n3604_n1904# a_12166_1472# a_9344_n1904#
+ a_n7588_n1904# a_n8086_1472# a_13992_n1904# a_n12236_n1904# a_n8916_n1904# a_n2940_1472#
+ a_1542_n1904# a_10174_n1904# a_11502_n1904# a_6854_n1904# a_712_n1904# a_3036_n1904#
+ a_n2608_n1904# a_8348_n1904# a_12996_n1904# a_11668_1472# a_n3272_1472# a_10340_1472#
+ a_n7588_1472# a_n6260_1472# a_3368_1472# a_10506_n1904# a_n9082_n1904# a_5858_n1904#
+ a_2040_1472# a_6356_1472# a_9344_1472# a_n1280_n1904# a_n6592_n1904# a_n11240_n1904#
+ a_n7920_n1904# a_n118_1472# a_n4102_n1904# a_n2774_1472# a_n8086_n1904# a_n5762_1472#
+ a_12830_1472# a_n9414_n1904# a_2040_n1904# a_n8750_1472# a_n11406_1472# a_1542_1472#
+ a_5858_1472# a_n1612_n1904# a_12000_n1904# a_4530_1472# a_8846_1472# a_7352_n1904#
+ a_n5596_n1904# a_n13896_1472# a_n10244_n1904# a_n6924_n1904# a_n3106_n1904# a_n450_n1904#
+ a_10174_1472# a_4862_n1904# a_13494_n1904# a_n6094_1472# a_13162_1472# a_n8418_n1904#
+ a_1044_n1904# a_n9082_1472# a_11004_n1904# a_n10908_1472# a_9178_1472# a_n782_1472#
+ a_6356_n1904# a_214_n1904# a_n5928_n1904# a_n3106_1472# a_n7090_n1904# a_3866_n1904#
+ a_12498_n1904# a_13826_n1904# a_n5596_1472# a_n1280_1472# a_12664_1472# a_10008_n1904#
+ a_n8584_1472# a_1376_1472# a_n14228_1472# a_4364_1472# a_7352_1472# a_n2110_n1904#
+ a_n6094_n1904# a_n7422_n1904# a_n2608_1472# a_380_1472# a_5360_n1904# a_n4932_n1904#
+ a_n3770_1472# a_n1114_n1904# a_n13564_n1904# a_3866_1472# a_n12402_1472# a_n5098_n1904#
+ a_2870_n1904# a_6854_1472# a_n6426_n1904# a_9842_1472# a_12830_n1904# a_10008_1472#
+ a_4364_n1904# a_12498_1472# a_n3936_n1904# a_n616_1472# a_11170_1472# a_9676_n1904#
+ a_n7090_1472# a_n12568_n1904# a_4198_1472# a_1874_n1904# a_7186_1472# a_n11904_1472#
+ a_11834_n1904# a_n1114_1472# a_3368_n1904# a_n4102_1472# a_n8418_1472# a_13328_n1904#
+ a_48_n1904# a_10672_1472# a_n6592_1472# a_13660_1472# a_n5430_n1904# a_n9580_1472#
+ a_n12236_1472# a_6688_1472# a_10838_n1904# a_2372_1472# a_n14062_n1904# a_5360_1472#
+ a_9676_1472# a_214_1472# a_n2940_n1904# a_8680_n1904# a_n3604_1472# a_n11572_n1904#
+ a_n12900_n1904# a_n4434_n1904# a_n11738_1472# a_n13066_n1904# a_n9746_n1904# a_1874_1472#
+ a_2372_n1904# a_n10410_1472# a_4862_1472# a_3700_n1904# a_n1944_n1904# a_12332_n1904#
+ a_7850_1472# a_7684_n1904# a_n10576_n1904# a_11004_1472# a_n11904_n1904# a_n3438_n1904#
X0 a_8016_1472# a_8016_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X1 a_n616_1472# a_n616_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X2 a_3368_1472# a_3368_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X3 a_1044_1472# a_1044_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X4 a_n6924_1472# a_n6924_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X5 a_n9746_1472# a_n9746_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X6 a_n7422_1472# a_n7422_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X7 a_546_1472# a_546_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X8 a_380_1472# a_380_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X9 a_n13896_1472# a_n13896_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X10 a_n11738_1472# a_n11738_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X11 a_n11572_1472# a_n11572_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X12 a_n2940_1472# a_n2940_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X13 a_n2774_1472# a_n2774_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X14 a_n12236_1472# a_n12236_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X15 a_13826_1472# a_13826_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X16 a_11502_1472# a_11502_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X17 a_n3438_1472# a_n3438_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X18 a_13660_1472# a_13660_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X19 a_7850_1472# a_7850_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X20 a_n1114_1472# a_n1114_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X21 a_n5596_1472# a_n5596_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X22 a_n3272_1472# a_n3272_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X23 a_12000_1472# a_12000_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X24 a_8514_1472# a_8514_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X25 a_n6260_1472# a_n6260_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X26 a_n6094_1472# a_n6094_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X27 a_3866_1472# a_3866_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X28 a_1708_1472# a_1708_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X29 a_1542_1472# a_1542_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X30 a_9012_1472# a_9012_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X31 a_12498_1472# a_12498_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X32 a_10174_1472# a_10174_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X33 a_6688_1472# a_6688_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X34 a_4364_1472# a_4364_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X35 a_2206_1472# a_2206_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X36 a_2040_1472# a_2040_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X37 a_5028_1472# a_5028_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X38 a_7186_1472# a_7186_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X39 a_n12734_1472# a_n12734_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X40 a_n450_1472# a_n450_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X41 a_n3936_1472# a_n3936_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X42 a_n284_1472# a_n284_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X43 a_n1612_1472# a_n1612_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X44 a_n13232_1472# a_n13232_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X45 a_n6758_1472# a_n6758_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X46 a_n4434_1472# a_n4434_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X47 a_48_1472# a_48_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X48 a_n6592_1472# a_n6592_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X49 a_9510_1472# a_9510_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X50 a_n9580_1472# a_n9580_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X51 a_n7256_1472# a_n7256_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X52 a_10838_1472# a_10838_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X53 a_2704_1472# a_2704_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X54 a_12996_1472# a_12996_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X55 a_10672_1472# a_10672_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X56 a_4862_1472# a_4862_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X57 a_n12070_1472# a_n12070_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X58 a_13494_1472# a_13494_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X59 a_11336_1472# a_11336_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X60 a_7684_1472# a_7684_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X61 a_5526_1472# a_5526_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X62 a_5360_1472# a_5360_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X63 a_3202_1472# a_3202_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X64 a_11170_1472# a_11170_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X65 a_14158_1472# a_14158_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X66 a_8348_1472# a_8348_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X67 a_8182_1472# a_8182_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X68 a_6024_1472# a_6024_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X69 a_n782_1472# a_n782_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X70 a_n948_1472# a_n948_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X71 a_1376_1472# a_1376_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X72 a_n4932_1472# a_n4932_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X73 a_4198_1472# a_4198_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X74 a_n7920_1472# a_n7920_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X75 a_n7754_1472# a_n7754_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X76 a_878_1472# a_878_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X77 a_n8418_1472# a_n8418_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X78 a_n8252_1472# a_n8252_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X79 a_n10410_1472# a_n10410_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X80 a_n12568_1472# a_n12568_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X81 a_n10244_1472# a_n10244_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X82 a_11834_1472# a_11834_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X83 a_3700_1472# a_3700_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X84 a_n3770_1472# a_n3770_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X85 a_13992_1472# a_13992_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X86 a_n1446_1472# a_n1446_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X87 a_n13066_1472# a_n13066_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X88 a_n2110_1472# a_n2110_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X89 a_12332_1472# a_12332_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X90 a_8846_1472# a_8846_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X91 a_6522_1472# a_6522_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X92 a_n4268_1472# a_n4268_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X93 a_8680_1472# a_8680_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X94 a_1874_1472# a_1874_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X95 a_9344_1472# a_9344_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X96 a_7020_1472# a_7020_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X97 a_n7090_1472# a_n7090_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X98 a_4696_1472# a_4696_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X99 a_2538_1472# a_2538_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X100 a_2372_1472# a_2372_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X101 a_5194_1472# a_5194_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X102 a_3036_1472# a_3036_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X103 a_n8916_1472# a_n8916_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X104 a_n10908_1472# a_n10908_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X105 a_n10742_1472# a_n10742_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X106 a_n9414_1472# a_n9414_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X107 a_n1944_1472# a_n1944_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X108 a_n13730_1472# a_n13730_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X109 a_n11406_1472# a_n11406_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X110 a_214_1472# a_214_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X111 a_n13564_1472# a_n13564_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X112 a_n4766_1472# a_n4766_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X113 a_n2608_1472# a_n2608_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X114 a_12830_1472# a_12830_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X115 a_n2442_1472# a_n2442_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X116 a_n14228_1472# a_n14228_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X117 a_n14062_1472# a_n14062_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X118 a_9842_1472# a_9842_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X119 a_n7588_1472# a_n7588_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X120 a_n5430_1472# a_n5430_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X121 a_n5264_1472# a_n5264_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X122 a_n3106_1472# a_n3106_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X123 a_2870_1472# a_2870_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X124 a_n8086_1472# a_n8086_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X125 a_n10078_1472# a_n10078_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X126 a_11668_1472# a_11668_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X127 a_5858_1472# a_5858_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X128 a_3534_1472# a_3534_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X129 a_1210_1472# a_1210_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X130 a_5692_1472# a_5692_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X131 a_n1280_1472# a_n1280_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X132 a_10008_1472# a_10008_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X133 a_12166_1472# a_12166_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X134 a_6356_1472# a_6356_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X135 a_4032_1472# a_4032_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X136 a_6190_1472# a_6190_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X137 a_n9912_1472# a_n9912_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X138 a_712_1472# a_712_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X139 a_n11904_1472# a_n11904_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X140 a_9178_1472# a_9178_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X141 a_n12402_1472# a_n12402_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X142 a_n118_1472# a_n118_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X143 a_n5928_1472# a_n5928_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X144 a_n3604_1472# a_n3604_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X145 a_n5762_1472# a_n5762_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X146 a_n8750_1472# a_n8750_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X147 a_n6426_1472# a_n6426_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X148 a_n4102_1472# a_n4102_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X149 a_n8584_1472# a_n8584_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X150 a_n12900_1472# a_n12900_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X151 a_n10576_1472# a_n10576_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X152 a_n1778_1472# a_n1778_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X153 a_n9248_1472# a_n9248_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X154 a_n11240_1472# a_n11240_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X155 a_n9082_1472# a_n9082_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X156 a_n13398_1472# a_n13398_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X157 a_n11074_1472# a_n11074_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X158 a_12664_1472# a_12664_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X159 a_10506_1472# a_10506_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X160 a_10340_1472# a_10340_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X161 a_6854_1472# a_6854_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X162 a_4530_1472# a_4530_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X163 a_n4600_1472# a_n4600_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X164 a_n2276_1472# a_n2276_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X165 a_13328_1472# a_13328_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X166 a_13162_1472# a_13162_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X167 a_11004_1472# a_11004_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X168 a_9676_1472# a_9676_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X169 a_7518_1472# a_7518_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X170 a_7352_1472# a_7352_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X171 a_n5098_1472# a_n5098_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_S4N9LQ a_1708_1984# a_n1778_n2416# a_712_1984#
+ a_n948_1984# a_2538_n2416# a_n1446_1984# a_n948_n2416# a_380_n2416# a_546_1984#
+ a_n2276_n2416# a_1542_n2416# a_712_n2416# a_n2608_n2416# a_n1280_n2416# a_n2442_1984#
+ a_2538_1984# a_1210_1984# a_2040_n2416# a_n1612_n2416# a_n1944_1984# a_n450_n2416#
+ a_1044_n2416# a_n450_1984# a_214_n2416# a_n2276_1984# a_1044_1984# a_n2110_n2416#
+ a_n1778_1984# a_n284_1984# a_n1114_n2416# a_878_1984# a_1874_n2416# a_48_n2416#
+ a_2040_1984# a_n118_1984# a_n2738_n2546# a_1542_1984# a_2372_n2416# a_n1944_n2416#
+ a_n782_n2416# a_n782_1984# a_1376_n2416# a_546_n2416# a_n1280_1984# a_1376_1984#
+ a_1708_n2416# a_n2442_n2416# a_n2608_1984# a_380_1984# a_n1446_n2416# a_n616_1984#
+ a_n284_n2416# a_2206_n2416# a_n1114_1984# a_n616_n2416# a_2372_1984# a_214_1984#
+ a_1210_n2416# a_1874_1984# a_878_n2416# a_n2110_1984# a_n118_n2416# a_2206_1984#
+ a_48_1984# a_n1612_1984#
X0 a_2040_1984# a_2040_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X1 a_2206_1984# a_2206_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X2 a_n450_1984# a_n450_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X3 a_n284_1984# a_n284_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X4 a_n1612_1984# a_n1612_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X5 a_48_1984# a_48_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X6 a_n948_1984# a_n948_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X7 a_n782_1984# a_n782_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X8 a_1376_1984# a_1376_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X9 a_878_1984# a_878_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X10 a_n1446_1984# a_n1446_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X11 a_n2110_1984# a_n2110_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X12 a_1874_1984# a_1874_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X13 a_2372_1984# a_2372_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X14 a_2538_1984# a_2538_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X15 a_n1944_1984# a_n1944_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X16 a_n2608_1984# a_n2608_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X17 a_n2442_1984# a_n2442_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X18 a_214_1984# a_214_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X19 a_n1280_1984# a_n1280_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X20 a_1210_1984# a_1210_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X21 a_712_1984# a_712_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X22 a_n118_1984# a_n118_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X23 a_n2276_1984# a_n2276_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X24 a_n1778_1984# a_n1778_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X25 a_n616_1984# a_n616_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X26 a_1044_1984# a_1044_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X27 a_546_1984# a_546_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X28 a_380_1984# a_380_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X29 a_n1114_1984# a_n1114_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X30 a_1542_1984# a_1542_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X31 a_1708_1984# a_1708_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
.ends

.subckt Parallel_10B_Block2 V6 V5 V8 V9 V7 VO1 VOUT V4 V3 V2 V0 VCM w_8036_n6718#
+ VBIAS V1 w_8040_12750# w_3572_3030# w_3570_n6718# w_8038_3030# w_3574_12750# w_7054_n6718#
+ w_7056_3030# DVDD DVSS AVSS AVDD w_7058_12750#
Xx1 V8 DVDD VCM x1/R2RIN x13/R2RIN x7/VINN AVSS DVSS AVDD Universal_R_2R_Block2
Xx2 V5 DVDD VCM x6/VOUT x5/R2RIN x7/VINN AVSS DVSS AVDD Universal_R_2R_Block2
Xx3 V2 DVDD VCM x3/R2RIN x3/R2ROUT x7/VINN AVSS DVSS AVDD Universal_R_2R_Block2
Xx4 V0 DVDD VCM x8/VOUT x4/R2ROUT x7/VINN AVSS DVSS AVDD Universal_R_2R_Block2
Xx5 V6 DVDD VCM x5/R2RIN x5/R2ROUT x7/VINN AVSS DVSS AVDD Universal_R_2R_Block2
Xx6 AVDD x6/VOUT x6/VINN VCM VBIAS w_3574_12750# w_7058_12750# AVSS w_8040_12750#
+ x1_x32_OA
Xx7 AVDD VOUT x7/VINN VCM VBIAS w_3570_n6718# w_7054_n6718# AVSS w_8036_n6718# Output_OA
Xx8 AVDD x8/VOUT x8/VINN VCM VBIAS w_3572_3030# w_7056_3030# AVSS w_8038_3030# x1_x32_OA
Xx9 V4 DVDD VCM x9/R2RIN x9/R2ROUT x7/VINN AVSS DVSS AVDD Universal_R_2R_Block2
Xsky130_fd_pr__res_xhigh_po_0p35_Q2LWZP_0 m1_13604_18506# VCM m1_13272_18506# m1_12290_20904#
+ AVSS m1_12940_18506# m1_13272_18506# m1_13438_20902# x13/R2ROUT m1_13604_18506#
+ m1_13438_20902# x6/VOUT m1_12940_18506# sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP
Xsky130_fd_pr__res_xhigh_po_0p35_Q2LWZP_1 m1_10646_18508# m1_10146_20906# m1_10314_18508#
+ x9/R2ROUT AVSS m1_9982_18508# m1_10314_18508# VCM VO1 m1_10646_18508# x8/VINN m1_10146_20906#
+ m1_9982_18508# sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP
Xsky130_fd_pr__res_xhigh_po_0p35_Q2LWZP_2 m1_12122_18506# m1_11626_20906# m1_11790_18506#
+ VO1 AVSS m1_11458_18506# m1_11790_18506# x6/VINN m1_12290_20904# m1_12122_18506#
+ x6/VINN m1_11626_20906# m1_11458_18506# sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP
Xx10 V3 DVDD VCM x3/R2ROUT x9/R2RIN x7/VINN AVSS DVSS AVDD Universal_R_2R_Block2
Xx11 V1 DVDD VCM x4/R2ROUT x3/R2RIN x7/VINN AVSS DVSS AVDD Universal_R_2R_Block2
Xx12 V7 DVDD VCM x5/R2ROUT x1/R2RIN x7/VINN AVSS DVSS AVDD Universal_R_2R_Block2
Xx13 V9 DVDD VCM x13/R2RIN x13/R2ROUT x7/VINN AVSS DVSS AVDD Universal_R_2R_Block2
Xsky130_fd_pr__res_xhigh_po_0p35_V6AMGK_0 m1_13942_n11110# m1_23902_n11110# m1_28384_n7734#
+ m1_16266_n11110# m1_17594_n11110# m1_20084_n7734# m1_26226_n11110# m1_23072_n7734#
+ m1_21578_n11110# m1_1824_n7734# m1_15270_n11110# m1_3982_n11110# m1_11452_n7734#
+ m1_25396_n7734# m1_8464_n7734# m1_12780_n7734# m1_2654_n11110# m1_5476_n7734# m1_5974_n11110#
+ m1_17096_n7734# m1_27720_n7734# m1_16598_n11110# m1_4480_n7734# m1_19420_n7734#
+ m1_1492_n7734# m1_22408_n7734# x7/VINN m1_12282_n11110# m1_22906_n11110# m1_24234_n11110#
+ m1_3650_n11110# m1_6970_n11110# m1_8796_n7734# m1_13112_n7734# m1_2322_n11110# m1_10124_n7734#
+ m1_5808_n7734# m1_16432_n7734# m1_25230_n11110# m1_20582_n11110# m1_5642_n11110#
+ m1_17926_n11110# m1_2156_n7734# m1_13278_n11110# m1_994_n11110# m1_17760_n7734#
+ m1_21910_n11110# m1_23238_n11110# m1_4646_n11110# m1_7966_n11110# m1_15436_n7734#
+ m1_28052_n7734# m1_3318_n11110# m1_26724_n7734# m1_5476_n7734# m1_14606_n11110#
+ m1_19586_n11110# m1_13776_n7734# m1_19752_n7734# m1_22740_n7734# m1_4812_n7734#
+ m1_16930_n11110# m1_1824_n7734# m1_21080_n7734# m1_22242_n11110# m1_13444_n7734#
+ m1_10456_n7734# m1_26392_n7734# m1_6638_n11110# m1_14274_n11110# m1_7468_n7734#
+ m1_18092_n7734# m1_22408_n7734# m1_28716_n7734# m1_20914_n11110# m1_2156_n7734#
+ m1_8962_n11110# m1_4314_n11110# m1_3484_n7734# m1_20416_n7734# m1_23404_n7734# m1_15436_n7734#
+ m1_23902_n11110# m1_7634_n11110# m1_28550_n11110# m1_10788_n7734# m1_15934_n11110#
+ m1_7800_n7734# m1_19918_n11110# m1_4812_n7734# m1_17428_n7734# m1_21246_n11110#
+ m1_9958_n11110# m1_4148_n7734# m1_1326_n11110# m1_1160_n7734# m1_22906_n11110# m1_27554_n11110#
+ m1_10456_n7734# m1_26060_n7734# m1_7468_n7734# m1_18922_n11110# m1_20250_n11110#
+ m1_17760_n7734# m1_28882_n11110# m1_20748_n7734# m1_23736_n7734# m1_3816_n7734#
+ m1_8630_n11110# m1_828_n7734# m1_26558_n11110# m1_15602_n11110# m1_25728_n7734#
+ m1_10954_n11110# m1_14606_n11110# m1_8132_n7734# m1_12448_n7734# m1_28716_n7734#
+ m1_5144_n7734# m1_9460_n7734# m1_17428_n7734# m1_994_n11110# m1_16100_n7734# m1_20416_n7734#
+ m1_21910_n11110# m1_9626_n11110# m1_23404_n7734# m1_4148_n7734# m1_1160_n7734# m1_19254_n11110#
+ m1_11950_n11110# VOUT m1_27886_n11110# m1_12780_n7734# m1_24566_n11110# m1_9792_n7734#
+ m1_1990_n11110# m1_20914_n11110# m1_6804_n7734# m1_10622_n11110# m1_14440_n7734#
+ m1_25562_n11110# m1_18424_n7734# m1_662_n11110# m1_18258_n11110# m1_12946_n11110#
+ m1_26890_n11110# m1_12448_n7734# m1_23570_n11110# m1_27056_n7734# m1_9460_n7734#
+ m1_2986_n11110# m1_19918_n11110# m1_6472_n7734# m1_15768_n7734# m1_18756_n7734#
+ m1_23072_n7734# m1_5310_n11110# m1_21744_n7734# m1_1492_n7734# m1_17262_n11110#
+ m1_2820_n7734# AVSS m1_11618_n11110# m1_13112_n7734# m1_10124_n7734# m1_10290_n11110#
+ m1_26724_n7734# m1_7136_n7734# m1_6306_n11110# m1_13942_n11110# m1_14440_n7734#
+ m1_1658_n11110# m1_4978_n11110# m1_18424_n7734# m1_25894_n11110# m1_21412_n7734#
+ m1_15270_n11110# m1_22574_n11110# m1_24400_n7734# m1_3152_n7734# m1_3982_n11110#
+ m1_18922_n11110# m1_12614_n11110# m1_15768_n7734# m1_9792_n7734# m1_11286_n11110#
+ m1_27056_n7734# m1_24234_n11110# m1_7302_n11110# m1_6804_n7734# m1_28882_n11110#
+ m1_2654_n11110# m1_5974_n11110# m1_11784_n7734# m1_16266_n11110# m1_24898_n11110#
+ m1_26226_n11110# m1_21578_n11110# m1_15602_n11110# m1_17926_n11110# m1_12282_n11110#
+ m1_23238_n11110# m1_27886_n11110# m1_26392_n7734# m1_11452_n7734# m1_25064_n7734#
+ m1_7136_n7734# m1_8464_n7734# m1_18092_n7734# m1_25230_n11110# m1_5642_n11110# m1_20582_n11110#
+ m1_16764_n7734# m1_21080_n7734# m1_24068_n7734# m1_13610_n11110# m1_8298_n11110#
+ m1_3650_n11110# m1_6970_n11110# x7/VINN m1_10622_n11110# m1_12116_n7734# m1_6638_n11110#
+ m1_9128_n7734# m1_27720_n7734# m1_5310_n11110# m1_16930_n11110# m1_6140_n7734# m1_3484_n7734#
+ m1_16432_n7734# m1_20748_n7734# m1_13278_n11110# m1_26890_n11110# m1_19420_n7734#
+ m1_23736_n7734# m1_22242_n11110# m1_9294_n11110# m1_828_n7734# m1_4646_n11110# m1_7966_n11110#
+ m1_11618_n11110# m1_14274_n11110# m1_25064_n7734# m1_19586_n11110# m1_28218_n11110#
+ m1_8796_n7734# m1_28052_n7734# m1_6306_n11110# m1_15934_n11110# m1_5808_n7734# m1_25894_n11110#
+ m1_3816_n7734# m1_24068_n7734# m1_14108_n7734# m1_21246_n11110# m1_14938_n11110#
+ m1_8962_n11110# m1_11784_n7734# m1_7634_n11110# m1_18590_n11110# m1_27222_n11110#
+ m1_28550_n11110# m1_9128_n7734# m1_13444_n7734# m1_27388_n7734# m1_24898_n11110#
+ m1_6140_n7734# m1_16100_n7734# x6/VOUT m1_19088_n7734# m1_22076_n7734# m1_12614_n11110#
+ m1_8630_n11110# m1_7302_n11110# m1_12116_n7734# m1_15104_n7734# m1_20250_n11110#
+ m1_9958_n11110# m1_11120_n7734# m1_13610_n11110# m1_1326_n11110# m1_18756_n7734#
+ m1_2488_n7734# m1_9626_n11110# m1_17594_n11110# m1_21744_n7734# m1_8298_n11110#
+ m1_24732_n7734# m1_27554_n11110# m1_24732_n7734# m1_19254_n11110# m1_27388_n7734#
+ m1_10954_n11110# m1_14108_n7734# m1_26060_n7734# m1_24566_n11110# m1_7800_n7734#
+ m1_2322_n11110# m1_19088_n7734# m1_16598_n11110# m1_22076_n7734# m1_2820_n7734#
+ m1_26558_n11110# m1_13776_n7734# m1_18258_n11110# m1_10788_n7734# m1_6472_n7734#
+ m1_28218_n11110# m1_14938_n11110# m1_25396_n7734# m1_8132_n7734# m1_28384_n7734#
+ m1_9294_n11110# m1_5144_n7734# m1_2488_n7734# m1_21412_n7734# m1_25562_n11110# m1_17096_n7734#
+ m1_662_n11110# m1_20084_n7734# m1_24400_n7734# m1_15104_n7734# m1_11950_n11110#
+ m1_23570_n11110# m1_11120_n7734# m1_3318_n11110# m1_1990_n11110# m1_10290_n11110#
+ m1_3152_n7734# m1_1658_n11110# m1_4978_n11110# m1_16764_n7734# m1_17262_n11110#
+ m1_4480_n7734# m1_19752_n7734# m1_18590_n11110# m1_12946_n11110# m1_27222_n11110#
+ m1_22740_n7734# m1_22574_n11110# m1_4314_n11110# m1_25728_n7734# m1_2986_n11110#
+ m1_11286_n11110# sky130_fd_pr__res_xhigh_po_0p35_V6AMGK
Xsky130_fd_pr__res_xhigh_po_0p35_S4N9LQ_0 m1_14152_11224# m1_10666_6824# m1_13156_11224#
+ m1_11496_11224# x8/VINN m1_10832_11224# m1_11330_6824# m1_12658_6824# m1_12824_11224#
+ m1_10002_6824# m1_13986_6824# m1_12990_6824# x8/VOUT m1_10998_6824# m1_9836_11224#
+ m1_14816_11224# m1_13488_11224# m1_14318_6824# m1_10666_6824# m1_10500_11224# m1_11994_6824#
+ m1_13322_6824# m1_11828_11224# m1_12658_6824# m1_10168_11224# m1_13488_11224# m1_10334_6824#
+ m1_10500_11224# m1_12160_11224# m1_11330_6824# m1_13156_11224# m1_14318_6824# m1_12326_6824#
+ m1_14484_11224# m1_12160_11224# AVSS m1_13820_11224# m1_14650_6824# m1_10334_6824#
+ m1_11662_6824# m1_11496_11224# m1_13654_6824# m1_12990_6824# m1_11164_11224# m1_13820_11224#
+ m1_13986_6824# m1_10002_6824# m1_9836_11224# m1_12824_11224# m1_10998_6824# m1_11828_11224#
+ m1_11994_6824# m1_14650_6824# m1_11164_11224# m1_11662_6824# m1_14816_11224# m1_12492_11224#
+ m1_13654_6824# m1_14152_11224# m1_13322_6824# m1_10168_11224# m1_12326_6824# m1_14484_11224#
+ m1_12492_11224# m1_10832_11224# sky130_fd_pr__res_xhigh_po_0p35_S4N9LQ
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_7WHXCK a_n29_n2720# a_487_n1610# a_n287_610#
+ a_229_n2720# a_n803_n2720# a_n287_n1610# a_n287_n500# a_229_1720# a_n745_n2808#
+ a_745_n500# a_n545_1720# a_745_n1610# a_n545_n1610# a_n803_610# a_229_n500# a_n29_n1610#
+ a_n29_1720# a_n229_n2808# a_n803_n1610# a_487_1720# a_487_n2720# a_229_n1610# a_n545_n500#
+ a_745_610# a_n287_n2720# a_229_610# a_n803_1720# a_n545_610# a_287_n2808# a_745_n2720#
+ a_n545_n2720# a_n29_n500# a_487_n500# a_n287_1720# a_487_610# a_n937_n2942# a_n29_610#
+ a_745_1720# a_n803_n500# a_545_n2808# a_29_n2808# a_n487_n2808#
X0 a_n29_610# a_n229_n2808# a_n287_610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X1 a_745_610# a_545_n2808# a_487_610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X2 a_745_n500# a_545_n2808# a_487_n500# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X3 a_487_1720# a_287_n2808# a_229_1720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X4 a_745_1720# a_545_n2808# a_487_1720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X5 a_487_n500# a_287_n2808# a_229_n500# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X6 a_229_610# a_29_n2808# a_n29_610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X7 a_n545_n2720# a_n745_n2808# a_n803_n2720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X8 a_229_n2720# a_29_n2808# a_n29_n2720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X9 a_487_610# a_287_n2808# a_229_610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X10 a_n545_610# a_n745_n2808# a_n803_610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X11 a_487_n1610# a_287_n2808# a_229_n1610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X12 a_n287_n1610# a_n487_n2808# a_n545_n1610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X13 a_229_n500# a_29_n2808# a_n29_n500# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X14 a_n29_n1610# a_n229_n2808# a_n287_n1610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X15 a_229_1720# a_29_n2808# a_n29_1720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X16 a_n29_n500# a_n229_n2808# a_n287_n500# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X17 a_n29_1720# a_n229_n2808# a_n287_1720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X18 a_n287_610# a_n487_n2808# a_n545_610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X19 a_745_n1610# a_545_n2808# a_487_n1610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X20 a_487_n2720# a_287_n2808# a_229_n2720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X21 a_n545_1720# a_n745_n2808# a_n803_1720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X22 a_n545_n500# a_n745_n2808# a_n803_n500# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X23 a_n287_n500# a_n487_n2808# a_n545_n500# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X24 a_n287_1720# a_n487_n2808# a_n545_1720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X25 a_n545_n1610# a_n745_n2808# a_n803_n1610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X26 a_229_n1610# a_29_n2808# a_n29_n1610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X27 a_n287_n2720# a_n487_n2808# a_n545_n2720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X28 a_n29_n2720# a_n229_n2808# a_n287_n2720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X29 a_745_n2720# a_545_n2808# a_487_n2720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
.ends

.subckt Input_Stage_OA1 VDD VOUT VINN VINP VBIAS w_8718_n902# w_7736_n902# VSS w_4240_n902#
XXR1 VSS m1_10706_1822# VOUT sky130_fd_pr__res_high_po_0p69_FJD3D2
Xsky130_fd_pr__nfet_05v0_nvt_FEJX3A_0 VINP VINP w_8718_n902# w_8718_n902# w_8718_n902#
+ m1_9368_n744# w_8718_n902# m1_9368_n744# w_8718_n902# VINP m1_9368_n744# m1_9368_n744#
+ VINP m1_9368_n744# m1_9368_n744# w_8718_n902# VINP w_8718_n902# m1_9368_n744# w_8718_n902#
+ VINP VINP w_8718_n902# w_8718_n902# m1_9368_n744# m1_9368_n744# w_8718_n902# w_8718_n902#
+ VINP VINP w_8718_n902# m1_9368_n744# m1_9368_n744# m1_9368_n744# VINP m1_9368_n744#
+ m1_9368_n744# VINP m1_9368_n744# m1_9368_n744# m1_9368_n744# VINP VINP w_8718_n902#
+ VINP VINP w_8718_n902# VINP VINP w_8718_n902# VINP w_8718_n902# w_8718_n902# VINP
+ m1_9368_n744# m1_9368_n744# VINP VINP w_8718_n902# m1_9368_n744# w_8718_n902# w_8718_n902#
+ w_8718_n902# VINP w_8718_n902# VINP w_8718_n902# m1_9368_n744# m1_9368_n744# w_8718_n902#
+ w_8718_n902# m1_9368_n744# VINP m1_9368_n744# VINP m1_9368_n744# sky130_fd_pr__nfet_05v0_nvt_FEJX3A
XXM2 VINN w_8718_n902# VINP w_7736_n902# w_7736_n902# w_4240_n902# w_7736_n902# sky130_fd_pr__nfet_01v8_lvt_AJ3MPE
XXM6 m1_9368_n744# m1_4902_n766# m1_9368_n744# VDD m1_4902_n766# m1_4902_n766# VDD
+ m1_4902_n766# m1_4902_n766# m1_4902_n766# VDD sky130_fd_pr__pfet_01v8_lvt_UX3DP3
XXM8 VDD VOUT VDD VOUT VDD VDD VOUT VDD m1_9368_n744# VDD VDD VOUT VOUT m1_9368_n744#
+ VDD VOUT m1_9368_n744# VOUT m1_9368_n744# m1_9368_n744# VOUT VDD m1_9368_n744# m1_9368_n744#
+ VDD VOUT VDD VOUT m1_9368_n744# m1_9368_n744# m1_9368_n744# sky130_fd_pr__pfet_g5v0d10v5_8UL4MK
Xsky130_fd_pr__cap_mim_m3_1_BHK9HY_0 m1_9368_n744# m1_9368_n744# m1_10706_1822# m1_10706_1822#
+ m1_10706_1822# m1_9368_n744# sky130_fd_pr__cap_mim_m3_1_BHK9HY
Xsky130_fd_pr__nfet_g5v0d10v5_7WHXCK_0 VOUT w_7736_n902# VSS VSS VSS VSS VSS VSS VBIAS
+ VSS VOUT VSS VOUT VSS VSS VOUT VOUT VBIAS VSS w_7736_n902# w_7736_n902# VSS VOUT
+ VSS VSS VSS VSS VOUT VBIAS VSS VOUT VOUT w_7736_n902# VSS w_7736_n902# VSS VOUT
+ VSS VSS VBIAS VBIAS VBIAS sky130_fd_pr__nfet_g5v0d10v5_7WHXCK
XXM10 VINN VINN m1_4902_n766# m1_4902_n766# m1_4902_n766# w_4240_n902# m1_4902_n766#
+ w_4240_n902# m1_4902_n766# VINN w_4240_n902# w_4240_n902# VINN w_4240_n902# w_4240_n902#
+ m1_4902_n766# VINN m1_4902_n766# w_4240_n902# m1_4902_n766# VINN VINN m1_4902_n766#
+ m1_4902_n766# w_4240_n902# w_4240_n902# m1_4902_n766# w_4240_n902# VINN VINN m1_4902_n766#
+ w_4240_n902# w_4240_n902# w_4240_n902# VINN w_4240_n902# w_4240_n902# VINN w_4240_n902#
+ w_4240_n902# w_4240_n902# VINN VINN m1_4902_n766# VINN VINN m1_4902_n766# VINN VINN
+ m1_4902_n766# VINN m1_4902_n766# m1_4902_n766# VINN w_4240_n902# w_4240_n902# VINN
+ VINN m1_4902_n766# w_4240_n902# m1_4902_n766# m1_4902_n766# m1_4902_n766# VINN m1_4902_n766#
+ VINN m1_4902_n766# w_4240_n902# w_4240_n902# m1_4902_n766# m1_4902_n766# w_4240_n902#
+ VINN w_4240_n902# VINN w_4240_n902# sky130_fd_pr__nfet_05v0_nvt_FEJX3A
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_KWU84Z a_n29_n2720# a_3067_1720# a_n287_610#
+ a_1261_n500# a_487_n1610# a_1777_1720# a_n2609_1720# a_n803_n2720# a_229_n2720#
+ a_n287_n1610# a_2867_n2808# a_n2351_1720# a_n1319_n500# a_n3125_610# a_n2609_610#
+ a_n287_n500# a_3067_n2720# a_229_1720# a_n1061_n500# a_n1577_1720# a_n3259_n2942#
+ a_2093_n2808# a_2551_610# a_2035_1720# a_n2351_n2720# a_1577_n2808# a_2551_n2720#
+ a_803_n2808# a_n745_n2808# a_n1003_n2808# a_3067_610# a_2809_n500# a_n1835_n2720#
+ a_745_n500# a_2035_610# a_n545_1720# a_1519_610# a_1003_610# a_745_n1610# a_2551_n500#
+ a_n1061_n2720# a_n545_n1610# a_1003_n1610# a_1261_n2720# a_3067_n500# a_1777_n500#
+ a_n2609_n500# a_1003_1720# a_n2293_n2808# a_n2867_n1610# a_n3125_n2720# a_n2351_610#
+ a_n2867_610# a_n1835_610# a_n2609_n2720# a_n1777_n2808# a_n2351_n500# a_2809_n2720#
+ a_2351_n2808# a_n2867_1720# a_n1319_610# a_1835_n2808# a_n803_610# a_229_n500# a_n2093_n1610#
+ a_2293_n1610# a_n1577_n500# a_n1577_n1610# a_2293_610# a_2035_n2720# a_n229_n2808#
+ a_1261_610# a_1777_610# a_2035_n500# a_n29_n1610# a_1777_n1610# a_n1319_n2720# a_n29_1720#
+ a_1519_n2720# a_487_1720# a_n3067_n2808# a_1061_n2808# a_n803_n1610# a_n545_n500#
+ a_229_n1610# a_487_n2720# a_2293_1720# a_n3125_1720# a_745_610# a_n1835_1720# a_n2551_n2808#
+ a_n287_n2720# a_2609_n2808# a_229_610# a_3067_n1610# a_n803_1720# a_n2093_610# a_1003_n500#
+ a_1519_1720# a_n1577_610# a_n2351_n1610# a_n1061_610# a_n2093_1720# a_2551_n1610#
+ a_n1261_n2808# a_n1835_n1610# a_1319_n2808# a_n2867_n500# a_1261_1720# a_n545_610#
+ a_287_n2808# a_n2809_n2808# a_745_n2720# a_n1061_n1610# a_n1319_1720# a_n29_n500#
+ a_1261_n1610# a_n545_n2720# a_487_n500# a_1003_n2720# a_n287_1720# a_n3125_n1610#
+ a_n1061_1720# a_487_610# a_n3125_n500# a_2293_n500# a_n2035_n2808# a_n2609_n1610#
+ a_n2867_n2720# a_n1835_n500# a_2809_n1610# a_n1519_n2808# a_2809_1720# a_n29_610#
+ a_745_1720# a_2809_610# a_n803_n500# a_n2093_n2720# a_2551_1720# a_1519_n500# a_2035_n1610#
+ a_545_n2808# a_n1319_n1610# a_2293_n2720# a_29_n2808# a_n487_n2808# a_n2093_n500#
+ a_n1577_n2720# a_1519_n1610# a_1777_n2720#
X0 a_n1061_1720# a_n1261_n2808# a_n1319_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X1 a_2551_n2720# a_2351_n2808# a_2293_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X2 a_1003_n500# a_803_n2808# a_745_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X3 a_n803_610# a_n1003_n2808# a_n1061_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X4 a_n1835_n2720# a_n2035_n2808# a_n2093_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X5 a_n803_n1610# a_n1003_n2808# a_n1061_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X6 a_745_610# a_545_n2808# a_487_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X7 a_1003_1720# a_803_n2808# a_745_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X8 a_745_n500# a_545_n2808# a_487_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X9 a_n29_610# a_n229_n2808# a_n287_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X10 a_1261_n2720# a_1061_n2808# a_1003_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X11 a_745_1720# a_545_n2808# a_487_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X12 a_487_n500# a_287_n2808# a_229_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X13 a_487_1720# a_287_n2808# a_229_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X14 a_229_n2720# a_29_n2808# a_n29_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X15 a_n545_n2720# a_n745_n2808# a_n803_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X16 a_229_610# a_29_n2808# a_n29_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X17 a_2035_n500# a_1835_n2808# a_1777_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X18 a_3067_n1610# a_2867_n2808# a_2809_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X19 a_2035_1720# a_1835_n2808# a_1777_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X20 a_1777_n500# a_1577_n2808# a_1519_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X21 a_n2609_n500# a_n2809_n2808# a_n2867_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X22 a_1777_1720# a_1577_n2808# a_1519_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X23 a_n2609_1720# a_n2809_n2808# a_n2867_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X24 a_2809_n1610# a_2609_n2808# a_2551_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X25 a_1519_610# a_1319_n2808# a_1261_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X26 a_1777_n1610# a_1577_n2808# a_1519_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X27 a_1261_n500# a_1061_n2808# a_1003_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X28 a_1261_1720# a_1061_n2808# a_1003_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X29 a_n1835_n500# a_n2035_n2808# a_n2093_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X30 a_1519_n1610# a_1319_n2808# a_1261_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X31 a_487_610# a_287_n2808# a_229_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X32 a_n1835_1720# a_n2035_n2808# a_n2093_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X33 a_n2351_n2720# a_n2551_n2808# a_n2609_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X34 a_1003_n2720# a_803_n2808# a_745_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X35 a_2809_610# a_2609_n2808# a_2551_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X36 a_n545_610# a_n745_n2808# a_n803_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X37 a_n2867_n1610# a_n3067_n2808# a_n3125_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X38 a_n1061_n2720# a_n1261_n2808# a_n1319_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X39 a_n1319_610# a_n1519_n2808# a_n1577_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X40 a_487_n1610# a_287_n2808# a_229_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X41 a_2293_n1610# a_2093_n2808# a_2035_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X42 a_n1835_610# a_n2035_n2808# a_n2093_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X43 a_n803_n2720# a_n1003_n2808# a_n1061_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X44 a_1261_610# a_1061_n2808# a_1003_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X45 a_2809_n500# a_2609_n2808# a_2551_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X46 a_2809_1720# a_2609_n2808# a_2551_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X47 a_n287_n1610# a_n487_n2808# a_n545_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X48 a_n2609_610# a_n2809_n2808# a_n2867_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X49 a_n2351_n500# a_n2551_n2808# a_n2609_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X50 a_n2609_n1610# a_n2809_n2808# a_n2867_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X51 a_n2351_1720# a_n2551_n2808# a_n2609_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X52 a_n2093_n500# a_n2293_n2808# a_n2351_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X53 a_2035_610# a_1835_n2808# a_1777_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X54 a_n29_n1610# a_n229_n2808# a_n287_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X55 a_n1577_n1610# a_n1777_n2808# a_n1835_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X56 a_229_n500# a_29_n2808# a_n29_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X57 a_n2093_1720# a_n2293_n2808# a_n2351_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X58 a_n29_n500# a_n229_n2808# a_n287_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X59 a_229_1720# a_29_n2808# a_n29_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X60 a_3067_n2720# a_2867_n2808# a_2809_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X61 a_2035_n1610# a_1835_n2808# a_1777_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X62 a_2551_610# a_2351_n2808# a_2293_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X63 a_n29_1720# a_n229_n2808# a_n287_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X64 a_n1319_n1610# a_n1519_n2808# a_n1577_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X65 a_n1061_610# a_n1261_n2808# a_n1319_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X66 a_2809_n2720# a_2609_n2808# a_2551_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X67 a_n287_610# a_n487_n2808# a_n545_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X68 a_1777_n2720# a_1577_n2808# a_1519_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X69 a_1519_n2720# a_1319_n2808# a_1261_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X70 a_n2093_n1610# a_n2293_n2808# a_n2351_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X71 a_745_n1610# a_545_n2808# a_487_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X72 a_n2351_610# a_n2551_n2808# a_n2609_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X73 a_3067_n500# a_2867_n2808# a_2809_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X74 a_2551_n1610# a_2351_n2808# a_2293_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X75 a_3067_1720# a_2867_n2808# a_2809_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X76 a_n2867_n2720# a_n3067_n2808# a_n3125_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X77 a_n1835_n1610# a_n2035_n2808# a_n2093_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X78 a_487_n2720# a_287_n2808# a_229_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X79 a_2551_n500# a_2351_n2808# a_2293_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X80 a_n1319_n500# a_n1519_n2808# a_n1577_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X81 a_2293_n2720# a_2093_n2808# a_2035_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X82 a_1261_n1610# a_1061_n2808# a_1003_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X83 a_n2867_610# a_n3067_n2808# a_n3125_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X84 a_2293_n500# a_2093_n2808# a_2035_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X85 a_n545_n500# a_n745_n2808# a_n803_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X86 a_1777_610# a_1577_n2808# a_1519_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X87 a_n1319_1720# a_n1519_n2808# a_n1577_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X88 a_2551_1720# a_2351_n2808# a_2293_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X89 a_n287_n500# a_n487_n2808# a_n545_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X90 a_n545_1720# a_n745_n2808# a_n803_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X91 a_2293_1720# a_2093_n2808# a_2035_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X92 a_2293_610# a_2093_n2808# a_2035_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X93 a_229_n1610# a_29_n2808# a_n29_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X94 a_n545_n1610# a_n745_n2808# a_n803_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X95 a_n803_n500# a_n1003_n2808# a_n1061_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X96 a_n2867_n500# a_n3067_n2808# a_n3125_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X97 a_n287_1720# a_n487_n2808# a_n545_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X98 a_n2867_1720# a_n3067_n2808# a_n3125_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X99 a_n803_1720# a_n1003_n2808# a_n1061_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X100 a_n287_n2720# a_n487_n2808# a_n545_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X101 a_1003_610# a_803_n2808# a_745_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X102 a_n2609_n2720# a_n2809_n2808# a_n2867_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X103 a_3067_610# a_2867_n2808# a_2809_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X104 a_n29_n2720# a_n229_n2808# a_n287_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X105 a_n1577_n2720# a_n1777_n2808# a_n1835_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X106 a_n1577_610# a_n1777_n2808# a_n1835_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X107 a_2035_n2720# a_1835_n2808# a_1777_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X108 a_n2093_610# a_n2293_n2808# a_n2351_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X109 a_n1319_n2720# a_n1519_n2808# a_n1577_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X110 a_n2351_n1610# a_n2551_n2808# a_n2609_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X111 a_n1577_n500# a_n1777_n2808# a_n1835_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X112 a_1003_n1610# a_803_n2808# a_745_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X113 a_1519_n500# a_1319_n2808# a_1261_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X114 a_n1577_1720# a_n1777_n2808# a_n1835_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X115 a_1519_1720# a_1319_n2808# a_1261_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X116 a_n2093_n2720# a_n2293_n2808# a_n2351_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X117 a_n1061_n1610# a_n1261_n2808# a_n1319_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X118 a_n1061_n500# a_n1261_n2808# a_n1319_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X119 a_745_n2720# a_545_n2808# a_487_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
.ends

.subckt Input_Stage_OA2 VDD VOUT VINN VINP VBIAS w_8718_n902# w_7736_n902# VSS w_4240_n902#
XXR1 VSS m1_10706_1822# VOUT sky130_fd_pr__res_high_po_0p69_FJD3D2
Xsky130_fd_pr__nfet_05v0_nvt_FEJX3A_0 VINP VINP w_8718_n902# w_8718_n902# w_8718_n902#
+ m1_9368_n744# w_8718_n902# m1_9368_n744# w_8718_n902# VINP m1_9368_n744# m1_9368_n744#
+ VINP m1_9368_n744# m1_9368_n744# w_8718_n902# VINP w_8718_n902# m1_9368_n744# w_8718_n902#
+ VINP VINP w_8718_n902# w_8718_n902# m1_9368_n744# m1_9368_n744# w_8718_n902# w_8718_n902#
+ VINP VINP w_8718_n902# m1_9368_n744# m1_9368_n744# m1_9368_n744# VINP m1_9368_n744#
+ m1_9368_n744# VINP m1_9368_n744# m1_9368_n744# m1_9368_n744# VINP VINP w_8718_n902#
+ VINP VINP w_8718_n902# VINP VINP w_8718_n902# VINP w_8718_n902# w_8718_n902# VINP
+ m1_9368_n744# m1_9368_n744# VINP VINP w_8718_n902# m1_9368_n744# w_8718_n902# w_8718_n902#
+ w_8718_n902# VINP w_8718_n902# VINP w_8718_n902# m1_9368_n744# m1_9368_n744# w_8718_n902#
+ w_8718_n902# m1_9368_n744# VINP m1_9368_n744# VINP m1_9368_n744# sky130_fd_pr__nfet_05v0_nvt_FEJX3A
XXM2 VINN w_8718_n902# VINP w_7736_n902# w_7736_n902# w_4240_n902# w_7736_n902# sky130_fd_pr__nfet_01v8_lvt_AJ3MPE
XXM6 m1_9368_n744# m1_4902_n766# m1_9368_n744# VDD m1_4902_n766# m1_4902_n766# VDD
+ m1_4902_n766# m1_4902_n766# m1_4902_n766# VDD sky130_fd_pr__pfet_01v8_lvt_UX3DP3
XXM8 VDD VOUT VDD VOUT VDD VDD VOUT VDD m1_9368_n744# VDD VDD VOUT VOUT m1_9368_n744#
+ VDD VOUT m1_9368_n744# VOUT m1_9368_n744# m1_9368_n744# VOUT VDD m1_9368_n744# m1_9368_n744#
+ VDD VOUT VDD VOUT m1_9368_n744# m1_9368_n744# m1_9368_n744# sky130_fd_pr__pfet_g5v0d10v5_8UL4MK
Xsky130_fd_pr__cap_mim_m3_1_BHK9HY_0 m1_9368_n744# m1_9368_n744# m1_10706_1822# m1_10706_1822#
+ m1_10706_1822# m1_9368_n744# sky130_fd_pr__cap_mim_m3_1_BHK9HY
XXM10 VINN VINN m1_4902_n766# m1_4902_n766# m1_4902_n766# w_4240_n902# m1_4902_n766#
+ w_4240_n902# m1_4902_n766# VINN w_4240_n902# w_4240_n902# VINN w_4240_n902# w_4240_n902#
+ m1_4902_n766# VINN m1_4902_n766# w_4240_n902# m1_4902_n766# VINN VINN m1_4902_n766#
+ m1_4902_n766# w_4240_n902# w_4240_n902# m1_4902_n766# w_4240_n902# VINN VINN m1_4902_n766#
+ w_4240_n902# w_4240_n902# w_4240_n902# VINN w_4240_n902# w_4240_n902# VINN w_4240_n902#
+ w_4240_n902# w_4240_n902# VINN VINN m1_4902_n766# VINN VINN m1_4902_n766# VINN VINN
+ m1_4902_n766# VINN m1_4902_n766# m1_4902_n766# VINN w_4240_n902# w_4240_n902# VINN
+ VINN m1_4902_n766# w_4240_n902# m1_4902_n766# m1_4902_n766# m1_4902_n766# VINN m1_4902_n766#
+ VINN m1_4902_n766# w_4240_n902# w_4240_n902# m1_4902_n766# m1_4902_n766# w_4240_n902#
+ VINN w_4240_n902# VINN w_4240_n902# sky130_fd_pr__nfet_05v0_nvt_FEJX3A
Xsky130_fd_pr__nfet_g5v0d10v5_KWU84Z_0 VSS VSS VOUT VOUT VSS VOUT VSS VOUT VOUT VOUT
+ VBIAS VOUT VOUT VSS VSS VOUT VSS VOUT VSS VSS VSS VBIAS VSS VSS VOUT VBIAS VSS VBIAS
+ VBIAS VBIAS VSS w_7736_n902# VOUT VOUT VSS VSS VSS VSS VOUT VSS VSS VSS VSS VOUT
+ VSS VOUT VSS VSS VBIAS VOUT VSS VOUT VOUT VOUT VSS VBIAS VOUT w_7736_n902# VBIAS
+ VOUT VOUT VBIAS VOUT VOUT VSS w_7736_n902# VSS VSS w_7736_n902# VSS VBIAS VOUT VOUT
+ VSS VSS VOUT VOUT VSS VSS VSS VBIAS VBIAS VOUT VSS VOUT VSS w_7736_n902# VSS VOUT
+ VOUT VBIAS VOUT VBIAS VOUT VSS VOUT VSS VSS VSS VSS VOUT VSS VSS VSS VBIAS VOUT
+ VBIAS VOUT VOUT VSS VBIAS VBIAS VOUT VSS VOUT VSS VOUT VSS VSS VSS VOUT VSS VSS
+ VSS VSS w_7736_n902# VBIAS VSS VOUT VOUT w_7736_n902# VBIAS w_7736_n902# VSS VOUT
+ w_7736_n902# VOUT VSS VSS VSS VSS VBIAS VOUT w_7736_n902# VBIAS VBIAS VSS VSS VSS
+ VOUT sky130_fd_pr__nfet_g5v0d10v5_KWU84Z
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_TVN32V a_3368_n2141# a_n118_1709# a_48_n2141#
+ a_n2774_1709# a_1542_1709# a_n2940_n2141# a_n782_1709# a_2372_n2141# a_3700_n2141#
+ a_n1944_n2141# a_n3106_1709# a_n3438_n2141# a_n782_n2141# a_n1280_1709# a_1376_1709#
+ a_1376_n2141# a_2704_n2141# a_546_n2141# a_n2608_1709# a_380_1709# a_n3770_1709#
+ a_1708_n2141# a_3866_1709# a_n2442_n2141# a_n616_1709# a_4198_1709# a_3202_n2141#
+ a_n1446_n2141# a_n1114_1709# a_n4102_1709# a_n284_n2141# a_2206_n2141# a_2372_1709#
+ a_214_1709# a_n3604_1709# a_n616_n2141# a_1874_1709# a_1210_n2141# a_n3438_1709#
+ a_n2110_1709# a_2206_1709# a_4198_n2141# a_48_1709# a_878_n2141# a_n118_n2141# a_n1612_1709#
+ a_n3770_n2141# a_1708_1709# a_2870_1709# a_712_1709# a_n2774_n2141# a_n948_1709#
+ a_n4268_n2141# a_3534_n2141# a_n1778_n2141# a_n1446_1709# a_3202_1709# a_2538_n2141#
+ a_546_1709# a_n3272_n2141# a_n3936_1709# a_n948_n2141# a_2704_1709# a_380_n2141#
+ a_4032_n2141# a_n2276_n2141# a_n3604_n2141# a_n4268_1709# a_1542_n2141# a_3036_1709#
+ a_712_n2141# a_3036_n2141# a_n2608_n2141# a_n2442_1709# a_2538_1709# a_1210_1709#
+ a_n1280_n2141# a_n4102_n2141# a_n1944_1709# a_n450_1709# a_2040_n2141# a_3700_1709#
+ a_n1612_n2141# a_n450_n2141# a_n2276_1709# a_n3106_n2141# a_1044_1709# a_1044_n2141#
+ a_4032_1709# a_214_n2141# a_3866_n2141# a_n1778_1709# a_n284_1709# a_3534_1709#
+ a_n4398_n2271# a_n2110_n2141# a_878_1709# a_n2940_1709# a_n1114_n2141# a_2870_n2141#
+ a_n3272_1709# a_n3936_n2141# a_1874_n2141# a_2040_1709# a_3368_1709#
X0 a_n782_1709# a_n782_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X1 a_1376_1709# a_1376_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X2 a_4198_1709# a_4198_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X3 a_878_1709# a_878_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X4 a_n3770_1709# a_n3770_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X5 a_n1446_1709# a_n1446_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X6 a_3700_1709# a_3700_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X7 a_n4268_1709# a_n4268_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X8 a_n2110_1709# a_n2110_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X9 a_1874_1709# a_1874_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X10 a_2372_1709# a_2372_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X11 a_2538_1709# a_2538_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X12 a_3036_1709# a_3036_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X13 a_n1944_1709# a_n1944_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X14 a_214_1709# a_214_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X15 a_n2608_1709# a_n2608_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X16 a_n2442_1709# a_n2442_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X17 a_n3106_1709# a_n3106_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X18 a_2870_1709# a_2870_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X19 a_1210_1709# a_1210_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X20 a_3534_1709# a_3534_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X21 a_n1280_1709# a_n1280_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X22 a_4032_1709# a_4032_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X23 a_712_1709# a_712_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X24 a_n3604_1709# a_n3604_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X25 a_n118_1709# a_n118_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X26 a_n4102_1709# a_n4102_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X27 a_n1778_1709# a_n1778_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X28 a_n2276_1709# a_n2276_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X29 a_n616_1709# a_n616_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X30 a_1044_1709# a_1044_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X31 a_3368_1709# a_3368_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X32 a_380_1709# a_380_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X33 a_546_1709# a_546_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X34 a_n2940_1709# a_n2940_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X35 a_n2774_1709# a_n2774_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X36 a_n3438_1709# a_n3438_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X37 a_n3272_1709# a_n3272_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X38 a_n1114_1709# a_n1114_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X39 a_1542_1709# a_1542_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X40 a_1708_1709# a_1708_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X41 a_3866_1709# a_3866_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X42 a_2040_1709# a_2040_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X43 a_2206_1709# a_2206_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X44 a_n3936_1709# a_n3936_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X45 a_n1612_1709# a_n1612_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X46 a_n450_1709# a_n450_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X47 a_n284_1709# a_n284_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X48 a_48_1709# a_48_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X49 a_2704_1709# a_2704_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X50 a_n948_1709# a_n948_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X51 a_3202_1709# a_3202_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_QHQRGL a_1044_n2396# a_214_n2396# a_n1446_1964#
+ a_546_1964# a_n2110_n2396# a_n1114_n2396# a_n2406_n2526# a_1874_n2396# a_1210_1964#
+ a_48_n2396# a_n1944_1964# a_n450_1964# a_1044_1964# a_n1944_n2396# a_n2276_1964#
+ a_1376_n2396# a_n782_n2396# a_n1778_1964# a_546_n2396# a_n284_1964# a_1708_n2396#
+ a_878_1964# a_2040_1964# a_n1446_n2396# a_2206_n2396# a_n118_1964# a_n284_n2396#
+ a_1542_1964# a_n616_n2396# a_n782_1964# a_1210_n2396# a_1376_1964# a_n1280_1964#
+ a_380_1964# a_878_n2396# a_n118_n2396# a_n616_1964# a_n1114_1964# a_214_1964# a_n1778_n2396#
+ a_1874_1964# a_n948_n2396# a_380_n2396# a_n2276_n2396# a_2206_1964# a_1542_n2396#
+ a_712_n2396# a_n2110_1964# a_48_1964# a_1708_1964# a_n1280_n2396# a_n1612_1964#
+ a_2040_n2396# a_712_1964# a_n1612_n2396# a_n450_n2396# a_n948_1964#
X0 a_1874_1964# a_1874_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X1 a_n1944_1964# a_n1944_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X2 a_214_1964# a_214_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X3 a_1210_1964# a_1210_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X4 a_n1280_1964# a_n1280_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X5 a_712_1964# a_712_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X6 a_n118_1964# a_n118_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X7 a_n1778_1964# a_n1778_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X8 a_n2276_1964# a_n2276_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X9 a_n616_1964# a_n616_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X10 a_1044_1964# a_1044_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X11 a_380_1964# a_380_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X12 a_546_1964# a_546_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X13 a_n1114_1964# a_n1114_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X14 a_1542_1964# a_1542_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X15 a_1708_1964# a_1708_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X16 a_2040_1964# a_2040_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X17 a_2206_1964# a_2206_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X18 a_n1612_1964# a_n1612_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X19 a_n450_1964# a_n450_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X20 a_n284_1964# a_n284_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X21 a_48_1964# a_48_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X22 a_n948_1964# a_n948_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X23 a_n782_1964# a_n782_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X24 a_1376_1964# a_1376_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X25 a_878_1964# a_878_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X26 a_n1446_1964# a_n1446_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X27 a_n2110_1964# a_n2110_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
.ends

.subckt Input_Stage_v1 VINP VOUT1 VINN CM VBIAS w_18276_n26882# w_22762_n17134# w_21780_n17134#
+ w_21772_n36602# w_22754_n36602# w_18284_n17134# w_21772_n26882# w_22754_n26882#
+ w_18276_n36602# AVSS AVDD
Xx1 AVDD x1/VOUT x1/VOUT VINN VBIAS w_22754_n36602# w_21772_n36602# AVSS w_18276_n36602#
+ Input_Stage_OA1
Xx2 AVDD x2/VOUT x2/VOUT VINP VBIAS w_22754_n26882# w_21772_n26882# AVSS w_18276_n26882#
+ Input_Stage_OA1
Xx3 AVDD VOUT1 x3/VINN x3/VINP VBIAS w_22762_n17134# w_21780_n17134# AVSS w_18284_n17134#
+ Input_Stage_OA2
Xsky130_fd_pr__res_xhigh_po_0p35_TVN32V_0 m1_23074_n22690# m1_19588_n18840# m1_19754_n22690#
+ m1_16932_n18840# m1_21248_n18840# m1_16766_n22690# m1_18924_n18840# m1_22078_n22690#
+ m1_23406_n22690# m1_17762_n22690# m1_16600_n18840# m1_16434_n22690# m1_19090_n22690#
+ m1_18592_n18840# m1_21248_n18840# m1_21082_n22690# m1_22410_n22690# m1_20418_n22690#
+ m1_17264_n18840# m1_20252_n18840# m1_15936_n18840# m1_21414_n22690# m1_23572_n18840#
+ m1_17430_n22690# m1_19256_n18840# m1_23904_n18840# m1_23074_n22690# m1_18426_n22690#
+ m1_18592_n18840# x3/VINP m1_19422_n22690# m1_22078_n22690# m1_22244_n18840# m1_19920_n18840#
+ m1_16268_n18840# m1_19090_n22690# m1_21580_n18840# m1_21082_n22690# m1_16268_n18840#
+ m1_17596_n18840# m1_21912_n18840# VINP m1_19920_n18840# m1_20750_n22690# m1_19754_n22690#
+ m1_18260_n18840# m1_16102_n22690# m1_21580_n18840# m1_22576_n18840# m1_20584_n18840#
+ m1_17098_n22690# m1_18924_n18840# m1_15606_n22692# m1_23406_n22690# m1_18094_n22690#
+ m1_18260_n18840# m1_22908_n18840# m1_22410_n22690# m1_20252_n18840# m1_16434_n22690#
+ m1_15936_n18840# m1_18758_n22690# m1_22576_n18840# m1_20086_n22690# m1_23738_n22690#
+ m1_17430_n22690# m1_16102_n22690# x2/VOUT m1_21414_n22690# m1_22908_n18840# m1_20418_n22690#
+ m1_22742_n22690# m1_17098_n22690# m1_17264_n18840# m1_22244_n18840# m1_20916_n18840#
+ m1_18426_n22690# m1_15606_n22692# m1_17928_n18840# m1_19256_n18840# m1_21746_n22690#
+ m1_23572_n18840# m1_18094_n22690# m1_19422_n22690# m1_17596_n18840# m1_16766_n22690#
+ m1_20916_n18840# m1_20750_n22690# m1_23904_n18840# m1_20086_n22690# m1_23738_n22690#
+ m1_17928_n18840# m1_19588_n18840# m1_23240_n18840# AVSS m1_17762_n22690# m1_20584_n18840#
+ m1_16932_n18840# m1_18758_n22690# m1_22742_n22690# m1_16600_n18840# CM m1_21746_n22690#
+ m1_21912_n18840# m1_23240_n18840# sky130_fd_pr__res_xhigh_po_0p35_TVN32V
Xsky130_fd_pr__res_xhigh_po_0p35_TVN32V_1 m1_23104_n32408# m1_19618_n28558# m1_19784_n32408#
+ m1_16962_n28558# m1_21278_n28558# m1_16796_n32408# m1_18954_n28558# m1_22108_n32408#
+ m1_23436_n32408# m1_17792_n32408# m1_16630_n28558# m1_16464_n32408# m1_19120_n32408#
+ m1_18622_n28558# m1_21278_n28558# m1_21112_n32408# m1_22440_n32408# m1_20448_n32408#
+ m1_17294_n28558# m1_20282_n28558# m1_15966_n28558# m1_21444_n32408# m1_23602_n28558#
+ m1_17460_n32408# m1_19286_n28558# m1_23934_n28558# m1_23104_n32408# m1_18456_n32408#
+ m1_18622_n28558# x3/VINN m1_19452_n32408# m1_22108_n32408# m1_22274_n28558# m1_19950_n28558#
+ m1_16298_n28558# m1_19120_n32408# m1_21610_n28558# m1_21112_n32408# m1_16298_n28558#
+ m1_17626_n28558# m1_21942_n28558# VINN m1_19950_n28558# m1_20780_n32408# m1_19784_n32408#
+ m1_18290_n28558# m1_16132_n32408# m1_21610_n28558# m1_22606_n28558# m1_20614_n28558#
+ m1_17128_n32408# m1_18954_n28558# m1_15634_n32408# m1_23436_n32408# m1_18124_n32408#
+ m1_18290_n28558# m1_22938_n28558# m1_22440_n32408# m1_20282_n28558# m1_16464_n32408#
+ m1_15966_n28558# m1_18788_n32408# m1_22606_n28558# m1_20116_n32408# m1_23768_n32408#
+ m1_17460_n32408# m1_16132_n32408# x1/VOUT m1_21444_n32408# m1_22938_n28558# m1_20448_n32408#
+ m1_22772_n32408# m1_17128_n32408# m1_17294_n28558# m1_22274_n28558# m1_20946_n28558#
+ m1_18456_n32408# m1_15634_n32408# m1_17958_n28558# m1_19286_n28558# m1_21776_n32408#
+ m1_23602_n28558# m1_18124_n32408# m1_19452_n32408# m1_17626_n28558# m1_16796_n32408#
+ m1_20946_n28558# m1_20780_n32408# m1_23934_n28558# m1_20116_n32408# m1_23768_n32408#
+ m1_17958_n28558# m1_19618_n28558# m1_23270_n28558# AVSS m1_17792_n32408# m1_20614_n28558#
+ m1_16962_n28558# m1_18788_n32408# m1_22772_n32408# m1_16630_n28558# CM m1_21776_n32408#
+ m1_21942_n28558# m1_23270_n28558# sky130_fd_pr__res_xhigh_po_0p35_TVN32V
Xsky130_fd_pr__res_xhigh_po_0p35_QHQRGL_0 m1_18184_n12946# m1_17520_n12946# m1_15694_n8586#
+ m1_17686_n8586# m1_15196_n12946# m1_16192_n12946# AVSS m1_19180_n12946# m1_18350_n8586#
+ CM m1_15362_n8586# m1_16690_n8586# m1_18350_n8586# m1_15196_n12946# m1_15030_n8586#
+ m1_18516_n12946# m1_16524_n12946# m1_15362_n8586# m1_17852_n12946# m1_17022_n8586#
+ m1_18848_n12946# m1_18018_n8586# m1_19346_n8586# m1_15860_n12946# x3/VINP m1_17022_n8586#
+ m1_16856_n12946# m1_18682_n8586# m1_16524_n12946# m1_16358_n8586# m1_18516_n12946#
+ m1_18682_n8586# m1_16026_n8586# m1_17686_n8586# m1_18184_n12946# x3/VINN m1_16690_n8586#
+ m1_16026_n8586# m1_17354_n8586# m1_15528_n12946# m1_19014_n8586# m1_16192_n12946#
+ m1_17520_n12946# VOUT1 m1_19346_n8586# m1_18848_n12946# m1_17852_n12946# m1_15030_n8586#
+ m1_17354_n8586# m1_19014_n8586# m1_15860_n12946# m1_15694_n8586# m1_19180_n12946#
+ m1_18018_n8586# m1_15528_n12946# m1_16856_n12946# m1_16358_n8586# sky130_fd_pr__res_xhigh_po_0p35_QHQRGL
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_TZT4V2 a_100_n500# a_n292_n722# a_n158_n500#
+ a_n100_n588#
X0 a_100_n500# a_n100_n588# a_n158_n500# a_n292_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
.ends

.subckt vbias_gen_pga VBIAS IBIAS VSS
XXM4 VSS VSS VBIAS VBIAS sky130_fd_pr__nfet_g5v0d10v5_TZT4V2
R0 IBIAS VBIAS sky130_fd_pr__res_generic_m1 w=1 l=0.08
.ends

.subckt sky130_pa_ip__instramp V[9] V[8] V[7] V[6] V[5] V[4] V[3] V[2] V[1] V[0] VCM
+ IBIAS AVDD VIN DVDD VOUT AVSS DVSS
Xx1 V[6] V[5] V[8] V[9] V[7] x1/VO1 VOUT V[4] V[3] V[2] V[0] VCM w_18452_4866# x3/VBIAS
+ V[1] w_18448_24334# w_22928_14614# w_22930_4866# w_18450_14614# w_22926_24334# w_21948_4866#
+ w_21946_14614# DVDD DVSS AVSS AVDD w_21944_24334# Parallel_10B_Block2
Xx2 VIN x1/VO1 VCM VCM x3/VBIAS w_7908_14586# w_3434_24334# w_6918_24334# w_6926_4866#
+ w_3442_4866# w_7900_24334# w_6926_14586# w_3442_14586# w_7908_4866# AVSS AVDD Input_Stage_v1
Xx3 x3/VBIAS IBIAS AVSS vbias_gen_pga
.ends

