magic
tech sky130A
magscale 1 2
timestamp 1729620069
<< pwell >>
rect -30070 -6050 30070 6050
<< psubdiff >>
rect -30034 5980 -29938 6014
rect 29938 5980 30034 6014
rect -30034 5918 -30000 5980
rect 30000 5918 30034 5980
rect -30034 -5980 -30000 -5918
rect 30000 -5980 30034 -5918
rect -30034 -6014 -29938 -5980
rect 29938 -6014 30034 -5980
<< psubdiffcont >>
rect -29938 5980 29938 6014
rect -30034 -5918 -30000 5918
rect 30000 -5918 30034 5918
rect -29938 -6014 29938 -5980
<< xpolycontact >>
rect -29904 5452 -29766 5884
rect -29904 52 -29766 484
rect -29670 5452 -29532 5884
rect -29670 52 -29532 484
rect -29436 5452 -29298 5884
rect -29436 52 -29298 484
rect -29202 5452 -29064 5884
rect -29202 52 -29064 484
rect -28968 5452 -28830 5884
rect -28968 52 -28830 484
rect -28734 5452 -28596 5884
rect -28734 52 -28596 484
rect -28500 5452 -28362 5884
rect -28500 52 -28362 484
rect -28266 5452 -28128 5884
rect -28266 52 -28128 484
rect -28032 5452 -27894 5884
rect -28032 52 -27894 484
rect -27798 5452 -27660 5884
rect -27798 52 -27660 484
rect -27564 5452 -27426 5884
rect -27564 52 -27426 484
rect -27330 5452 -27192 5884
rect -27330 52 -27192 484
rect -27096 5452 -26958 5884
rect -27096 52 -26958 484
rect -26862 5452 -26724 5884
rect -26862 52 -26724 484
rect -26628 5452 -26490 5884
rect -26628 52 -26490 484
rect -26394 5452 -26256 5884
rect -26394 52 -26256 484
rect -26160 5452 -26022 5884
rect -26160 52 -26022 484
rect -25926 5452 -25788 5884
rect -25926 52 -25788 484
rect -25692 5452 -25554 5884
rect -25692 52 -25554 484
rect -25458 5452 -25320 5884
rect -25458 52 -25320 484
rect -25224 5452 -25086 5884
rect -25224 52 -25086 484
rect -24990 5452 -24852 5884
rect -24990 52 -24852 484
rect -24756 5452 -24618 5884
rect -24756 52 -24618 484
rect -24522 5452 -24384 5884
rect -24522 52 -24384 484
rect -24288 5452 -24150 5884
rect -24288 52 -24150 484
rect -24054 5452 -23916 5884
rect -24054 52 -23916 484
rect -23820 5452 -23682 5884
rect -23820 52 -23682 484
rect -23586 5452 -23448 5884
rect -23586 52 -23448 484
rect -23352 5452 -23214 5884
rect -23352 52 -23214 484
rect -23118 5452 -22980 5884
rect -23118 52 -22980 484
rect -22884 5452 -22746 5884
rect -22884 52 -22746 484
rect -22650 5452 -22512 5884
rect -22650 52 -22512 484
rect -22416 5452 -22278 5884
rect -22416 52 -22278 484
rect -22182 5452 -22044 5884
rect -22182 52 -22044 484
rect -21948 5452 -21810 5884
rect -21948 52 -21810 484
rect -21714 5452 -21576 5884
rect -21714 52 -21576 484
rect -21480 5452 -21342 5884
rect -21480 52 -21342 484
rect -21246 5452 -21108 5884
rect -21246 52 -21108 484
rect -21012 5452 -20874 5884
rect -21012 52 -20874 484
rect -20778 5452 -20640 5884
rect -20778 52 -20640 484
rect -20544 5452 -20406 5884
rect -20544 52 -20406 484
rect -20310 5452 -20172 5884
rect -20310 52 -20172 484
rect -20076 5452 -19938 5884
rect -20076 52 -19938 484
rect -19842 5452 -19704 5884
rect -19842 52 -19704 484
rect -19608 5452 -19470 5884
rect -19608 52 -19470 484
rect -19374 5452 -19236 5884
rect -19374 52 -19236 484
rect -19140 5452 -19002 5884
rect -19140 52 -19002 484
rect -18906 5452 -18768 5884
rect -18906 52 -18768 484
rect -18672 5452 -18534 5884
rect -18672 52 -18534 484
rect -18438 5452 -18300 5884
rect -18438 52 -18300 484
rect -18204 5452 -18066 5884
rect -18204 52 -18066 484
rect -17970 5452 -17832 5884
rect -17970 52 -17832 484
rect -17736 5452 -17598 5884
rect -17736 52 -17598 484
rect -17502 5452 -17364 5884
rect -17502 52 -17364 484
rect -17268 5452 -17130 5884
rect -17268 52 -17130 484
rect -17034 5452 -16896 5884
rect -17034 52 -16896 484
rect -16800 5452 -16662 5884
rect -16800 52 -16662 484
rect -16566 5452 -16428 5884
rect -16566 52 -16428 484
rect -16332 5452 -16194 5884
rect -16332 52 -16194 484
rect -16098 5452 -15960 5884
rect -16098 52 -15960 484
rect -15864 5452 -15726 5884
rect -15864 52 -15726 484
rect -15630 5452 -15492 5884
rect -15630 52 -15492 484
rect -15396 5452 -15258 5884
rect -15396 52 -15258 484
rect -15162 5452 -15024 5884
rect -15162 52 -15024 484
rect -14928 5452 -14790 5884
rect -14928 52 -14790 484
rect -14694 5452 -14556 5884
rect -14694 52 -14556 484
rect -14460 5452 -14322 5884
rect -14460 52 -14322 484
rect -14226 5452 -14088 5884
rect -14226 52 -14088 484
rect -13992 5452 -13854 5884
rect -13992 52 -13854 484
rect -13758 5452 -13620 5884
rect -13758 52 -13620 484
rect -13524 5452 -13386 5884
rect -13524 52 -13386 484
rect -13290 5452 -13152 5884
rect -13290 52 -13152 484
rect -13056 5452 -12918 5884
rect -13056 52 -12918 484
rect -12822 5452 -12684 5884
rect -12822 52 -12684 484
rect -12588 5452 -12450 5884
rect -12588 52 -12450 484
rect -12354 5452 -12216 5884
rect -12354 52 -12216 484
rect -12120 5452 -11982 5884
rect -12120 52 -11982 484
rect -11886 5452 -11748 5884
rect -11886 52 -11748 484
rect -11652 5452 -11514 5884
rect -11652 52 -11514 484
rect -11418 5452 -11280 5884
rect -11418 52 -11280 484
rect -11184 5452 -11046 5884
rect -11184 52 -11046 484
rect -10950 5452 -10812 5884
rect -10950 52 -10812 484
rect -10716 5452 -10578 5884
rect -10716 52 -10578 484
rect -10482 5452 -10344 5884
rect -10482 52 -10344 484
rect -10248 5452 -10110 5884
rect -10248 52 -10110 484
rect -10014 5452 -9876 5884
rect -10014 52 -9876 484
rect -9780 5452 -9642 5884
rect -9780 52 -9642 484
rect -9546 5452 -9408 5884
rect -9546 52 -9408 484
rect -9312 5452 -9174 5884
rect -9312 52 -9174 484
rect -9078 5452 -8940 5884
rect -9078 52 -8940 484
rect -8844 5452 -8706 5884
rect -8844 52 -8706 484
rect -8610 5452 -8472 5884
rect -8610 52 -8472 484
rect -8376 5452 -8238 5884
rect -8376 52 -8238 484
rect -8142 5452 -8004 5884
rect -8142 52 -8004 484
rect -7908 5452 -7770 5884
rect -7908 52 -7770 484
rect -7674 5452 -7536 5884
rect -7674 52 -7536 484
rect -7440 5452 -7302 5884
rect -7440 52 -7302 484
rect -7206 5452 -7068 5884
rect -7206 52 -7068 484
rect -6972 5452 -6834 5884
rect -6972 52 -6834 484
rect -6738 5452 -6600 5884
rect -6738 52 -6600 484
rect -6504 5452 -6366 5884
rect -6504 52 -6366 484
rect -6270 5452 -6132 5884
rect -6270 52 -6132 484
rect -6036 5452 -5898 5884
rect -6036 52 -5898 484
rect -5802 5452 -5664 5884
rect -5802 52 -5664 484
rect -5568 5452 -5430 5884
rect -5568 52 -5430 484
rect -5334 5452 -5196 5884
rect -5334 52 -5196 484
rect -5100 5452 -4962 5884
rect -5100 52 -4962 484
rect -4866 5452 -4728 5884
rect -4866 52 -4728 484
rect -4632 5452 -4494 5884
rect -4632 52 -4494 484
rect -4398 5452 -4260 5884
rect -4398 52 -4260 484
rect -4164 5452 -4026 5884
rect -4164 52 -4026 484
rect -3930 5452 -3792 5884
rect -3930 52 -3792 484
rect -3696 5452 -3558 5884
rect -3696 52 -3558 484
rect -3462 5452 -3324 5884
rect -3462 52 -3324 484
rect -3228 5452 -3090 5884
rect -3228 52 -3090 484
rect -2994 5452 -2856 5884
rect -2994 52 -2856 484
rect -2760 5452 -2622 5884
rect -2760 52 -2622 484
rect -2526 5452 -2388 5884
rect -2526 52 -2388 484
rect -2292 5452 -2154 5884
rect -2292 52 -2154 484
rect -2058 5452 -1920 5884
rect -2058 52 -1920 484
rect -1824 5452 -1686 5884
rect -1824 52 -1686 484
rect -1590 5452 -1452 5884
rect -1590 52 -1452 484
rect -1356 5452 -1218 5884
rect -1356 52 -1218 484
rect -1122 5452 -984 5884
rect -1122 52 -984 484
rect -888 5452 -750 5884
rect -888 52 -750 484
rect -654 5452 -516 5884
rect -654 52 -516 484
rect -420 5452 -282 5884
rect -420 52 -282 484
rect -186 5452 -48 5884
rect -186 52 -48 484
rect 48 5452 186 5884
rect 48 52 186 484
rect 282 5452 420 5884
rect 282 52 420 484
rect 516 5452 654 5884
rect 516 52 654 484
rect 750 5452 888 5884
rect 750 52 888 484
rect 984 5452 1122 5884
rect 984 52 1122 484
rect 1218 5452 1356 5884
rect 1218 52 1356 484
rect 1452 5452 1590 5884
rect 1452 52 1590 484
rect 1686 5452 1824 5884
rect 1686 52 1824 484
rect 1920 5452 2058 5884
rect 1920 52 2058 484
rect 2154 5452 2292 5884
rect 2154 52 2292 484
rect 2388 5452 2526 5884
rect 2388 52 2526 484
rect 2622 5452 2760 5884
rect 2622 52 2760 484
rect 2856 5452 2994 5884
rect 2856 52 2994 484
rect 3090 5452 3228 5884
rect 3090 52 3228 484
rect 3324 5452 3462 5884
rect 3324 52 3462 484
rect 3558 5452 3696 5884
rect 3558 52 3696 484
rect 3792 5452 3930 5884
rect 3792 52 3930 484
rect 4026 5452 4164 5884
rect 4026 52 4164 484
rect 4260 5452 4398 5884
rect 4260 52 4398 484
rect 4494 5452 4632 5884
rect 4494 52 4632 484
rect 4728 5452 4866 5884
rect 4728 52 4866 484
rect 4962 5452 5100 5884
rect 4962 52 5100 484
rect 5196 5452 5334 5884
rect 5196 52 5334 484
rect 5430 5452 5568 5884
rect 5430 52 5568 484
rect 5664 5452 5802 5884
rect 5664 52 5802 484
rect 5898 5452 6036 5884
rect 5898 52 6036 484
rect 6132 5452 6270 5884
rect 6132 52 6270 484
rect 6366 5452 6504 5884
rect 6366 52 6504 484
rect 6600 5452 6738 5884
rect 6600 52 6738 484
rect 6834 5452 6972 5884
rect 6834 52 6972 484
rect 7068 5452 7206 5884
rect 7068 52 7206 484
rect 7302 5452 7440 5884
rect 7302 52 7440 484
rect 7536 5452 7674 5884
rect 7536 52 7674 484
rect 7770 5452 7908 5884
rect 7770 52 7908 484
rect 8004 5452 8142 5884
rect 8004 52 8142 484
rect 8238 5452 8376 5884
rect 8238 52 8376 484
rect 8472 5452 8610 5884
rect 8472 52 8610 484
rect 8706 5452 8844 5884
rect 8706 52 8844 484
rect 8940 5452 9078 5884
rect 8940 52 9078 484
rect 9174 5452 9312 5884
rect 9174 52 9312 484
rect 9408 5452 9546 5884
rect 9408 52 9546 484
rect 9642 5452 9780 5884
rect 9642 52 9780 484
rect 9876 5452 10014 5884
rect 9876 52 10014 484
rect 10110 5452 10248 5884
rect 10110 52 10248 484
rect 10344 5452 10482 5884
rect 10344 52 10482 484
rect 10578 5452 10716 5884
rect 10578 52 10716 484
rect 10812 5452 10950 5884
rect 10812 52 10950 484
rect 11046 5452 11184 5884
rect 11046 52 11184 484
rect 11280 5452 11418 5884
rect 11280 52 11418 484
rect 11514 5452 11652 5884
rect 11514 52 11652 484
rect 11748 5452 11886 5884
rect 11748 52 11886 484
rect 11982 5452 12120 5884
rect 11982 52 12120 484
rect 12216 5452 12354 5884
rect 12216 52 12354 484
rect 12450 5452 12588 5884
rect 12450 52 12588 484
rect 12684 5452 12822 5884
rect 12684 52 12822 484
rect 12918 5452 13056 5884
rect 12918 52 13056 484
rect 13152 5452 13290 5884
rect 13152 52 13290 484
rect 13386 5452 13524 5884
rect 13386 52 13524 484
rect 13620 5452 13758 5884
rect 13620 52 13758 484
rect 13854 5452 13992 5884
rect 13854 52 13992 484
rect 14088 5452 14226 5884
rect 14088 52 14226 484
rect 14322 5452 14460 5884
rect 14322 52 14460 484
rect 14556 5452 14694 5884
rect 14556 52 14694 484
rect 14790 5452 14928 5884
rect 14790 52 14928 484
rect 15024 5452 15162 5884
rect 15024 52 15162 484
rect 15258 5452 15396 5884
rect 15258 52 15396 484
rect 15492 5452 15630 5884
rect 15492 52 15630 484
rect 15726 5452 15864 5884
rect 15726 52 15864 484
rect 15960 5452 16098 5884
rect 15960 52 16098 484
rect 16194 5452 16332 5884
rect 16194 52 16332 484
rect 16428 5452 16566 5884
rect 16428 52 16566 484
rect 16662 5452 16800 5884
rect 16662 52 16800 484
rect 16896 5452 17034 5884
rect 16896 52 17034 484
rect 17130 5452 17268 5884
rect 17130 52 17268 484
rect 17364 5452 17502 5884
rect 17364 52 17502 484
rect 17598 5452 17736 5884
rect 17598 52 17736 484
rect 17832 5452 17970 5884
rect 17832 52 17970 484
rect 18066 5452 18204 5884
rect 18066 52 18204 484
rect 18300 5452 18438 5884
rect 18300 52 18438 484
rect 18534 5452 18672 5884
rect 18534 52 18672 484
rect 18768 5452 18906 5884
rect 18768 52 18906 484
rect 19002 5452 19140 5884
rect 19002 52 19140 484
rect 19236 5452 19374 5884
rect 19236 52 19374 484
rect 19470 5452 19608 5884
rect 19470 52 19608 484
rect 19704 5452 19842 5884
rect 19704 52 19842 484
rect 19938 5452 20076 5884
rect 19938 52 20076 484
rect 20172 5452 20310 5884
rect 20172 52 20310 484
rect 20406 5452 20544 5884
rect 20406 52 20544 484
rect 20640 5452 20778 5884
rect 20640 52 20778 484
rect 20874 5452 21012 5884
rect 20874 52 21012 484
rect 21108 5452 21246 5884
rect 21108 52 21246 484
rect 21342 5452 21480 5884
rect 21342 52 21480 484
rect 21576 5452 21714 5884
rect 21576 52 21714 484
rect 21810 5452 21948 5884
rect 21810 52 21948 484
rect 22044 5452 22182 5884
rect 22044 52 22182 484
rect 22278 5452 22416 5884
rect 22278 52 22416 484
rect 22512 5452 22650 5884
rect 22512 52 22650 484
rect 22746 5452 22884 5884
rect 22746 52 22884 484
rect 22980 5452 23118 5884
rect 22980 52 23118 484
rect 23214 5452 23352 5884
rect 23214 52 23352 484
rect 23448 5452 23586 5884
rect 23448 52 23586 484
rect 23682 5452 23820 5884
rect 23682 52 23820 484
rect 23916 5452 24054 5884
rect 23916 52 24054 484
rect 24150 5452 24288 5884
rect 24150 52 24288 484
rect 24384 5452 24522 5884
rect 24384 52 24522 484
rect 24618 5452 24756 5884
rect 24618 52 24756 484
rect 24852 5452 24990 5884
rect 24852 52 24990 484
rect 25086 5452 25224 5884
rect 25086 52 25224 484
rect 25320 5452 25458 5884
rect 25320 52 25458 484
rect 25554 5452 25692 5884
rect 25554 52 25692 484
rect 25788 5452 25926 5884
rect 25788 52 25926 484
rect 26022 5452 26160 5884
rect 26022 52 26160 484
rect 26256 5452 26394 5884
rect 26256 52 26394 484
rect 26490 5452 26628 5884
rect 26490 52 26628 484
rect 26724 5452 26862 5884
rect 26724 52 26862 484
rect 26958 5452 27096 5884
rect 26958 52 27096 484
rect 27192 5452 27330 5884
rect 27192 52 27330 484
rect 27426 5452 27564 5884
rect 27426 52 27564 484
rect 27660 5452 27798 5884
rect 27660 52 27798 484
rect 27894 5452 28032 5884
rect 27894 52 28032 484
rect 28128 5452 28266 5884
rect 28128 52 28266 484
rect 28362 5452 28500 5884
rect 28362 52 28500 484
rect 28596 5452 28734 5884
rect 28596 52 28734 484
rect 28830 5452 28968 5884
rect 28830 52 28968 484
rect 29064 5452 29202 5884
rect 29064 52 29202 484
rect 29298 5452 29436 5884
rect 29298 52 29436 484
rect 29532 5452 29670 5884
rect 29532 52 29670 484
rect 29766 5452 29904 5884
rect 29766 52 29904 484
rect -29904 -484 -29766 -52
rect -29904 -5884 -29766 -5452
rect -29670 -484 -29532 -52
rect -29670 -5884 -29532 -5452
rect -29436 -484 -29298 -52
rect -29436 -5884 -29298 -5452
rect -29202 -484 -29064 -52
rect -29202 -5884 -29064 -5452
rect -28968 -484 -28830 -52
rect -28968 -5884 -28830 -5452
rect -28734 -484 -28596 -52
rect -28734 -5884 -28596 -5452
rect -28500 -484 -28362 -52
rect -28500 -5884 -28362 -5452
rect -28266 -484 -28128 -52
rect -28266 -5884 -28128 -5452
rect -28032 -484 -27894 -52
rect -28032 -5884 -27894 -5452
rect -27798 -484 -27660 -52
rect -27798 -5884 -27660 -5452
rect -27564 -484 -27426 -52
rect -27564 -5884 -27426 -5452
rect -27330 -484 -27192 -52
rect -27330 -5884 -27192 -5452
rect -27096 -484 -26958 -52
rect -27096 -5884 -26958 -5452
rect -26862 -484 -26724 -52
rect -26862 -5884 -26724 -5452
rect -26628 -484 -26490 -52
rect -26628 -5884 -26490 -5452
rect -26394 -484 -26256 -52
rect -26394 -5884 -26256 -5452
rect -26160 -484 -26022 -52
rect -26160 -5884 -26022 -5452
rect -25926 -484 -25788 -52
rect -25926 -5884 -25788 -5452
rect -25692 -484 -25554 -52
rect -25692 -5884 -25554 -5452
rect -25458 -484 -25320 -52
rect -25458 -5884 -25320 -5452
rect -25224 -484 -25086 -52
rect -25224 -5884 -25086 -5452
rect -24990 -484 -24852 -52
rect -24990 -5884 -24852 -5452
rect -24756 -484 -24618 -52
rect -24756 -5884 -24618 -5452
rect -24522 -484 -24384 -52
rect -24522 -5884 -24384 -5452
rect -24288 -484 -24150 -52
rect -24288 -5884 -24150 -5452
rect -24054 -484 -23916 -52
rect -24054 -5884 -23916 -5452
rect -23820 -484 -23682 -52
rect -23820 -5884 -23682 -5452
rect -23586 -484 -23448 -52
rect -23586 -5884 -23448 -5452
rect -23352 -484 -23214 -52
rect -23352 -5884 -23214 -5452
rect -23118 -484 -22980 -52
rect -23118 -5884 -22980 -5452
rect -22884 -484 -22746 -52
rect -22884 -5884 -22746 -5452
rect -22650 -484 -22512 -52
rect -22650 -5884 -22512 -5452
rect -22416 -484 -22278 -52
rect -22416 -5884 -22278 -5452
rect -22182 -484 -22044 -52
rect -22182 -5884 -22044 -5452
rect -21948 -484 -21810 -52
rect -21948 -5884 -21810 -5452
rect -21714 -484 -21576 -52
rect -21714 -5884 -21576 -5452
rect -21480 -484 -21342 -52
rect -21480 -5884 -21342 -5452
rect -21246 -484 -21108 -52
rect -21246 -5884 -21108 -5452
rect -21012 -484 -20874 -52
rect -21012 -5884 -20874 -5452
rect -20778 -484 -20640 -52
rect -20778 -5884 -20640 -5452
rect -20544 -484 -20406 -52
rect -20544 -5884 -20406 -5452
rect -20310 -484 -20172 -52
rect -20310 -5884 -20172 -5452
rect -20076 -484 -19938 -52
rect -20076 -5884 -19938 -5452
rect -19842 -484 -19704 -52
rect -19842 -5884 -19704 -5452
rect -19608 -484 -19470 -52
rect -19608 -5884 -19470 -5452
rect -19374 -484 -19236 -52
rect -19374 -5884 -19236 -5452
rect -19140 -484 -19002 -52
rect -19140 -5884 -19002 -5452
rect -18906 -484 -18768 -52
rect -18906 -5884 -18768 -5452
rect -18672 -484 -18534 -52
rect -18672 -5884 -18534 -5452
rect -18438 -484 -18300 -52
rect -18438 -5884 -18300 -5452
rect -18204 -484 -18066 -52
rect -18204 -5884 -18066 -5452
rect -17970 -484 -17832 -52
rect -17970 -5884 -17832 -5452
rect -17736 -484 -17598 -52
rect -17736 -5884 -17598 -5452
rect -17502 -484 -17364 -52
rect -17502 -5884 -17364 -5452
rect -17268 -484 -17130 -52
rect -17268 -5884 -17130 -5452
rect -17034 -484 -16896 -52
rect -17034 -5884 -16896 -5452
rect -16800 -484 -16662 -52
rect -16800 -5884 -16662 -5452
rect -16566 -484 -16428 -52
rect -16566 -5884 -16428 -5452
rect -16332 -484 -16194 -52
rect -16332 -5884 -16194 -5452
rect -16098 -484 -15960 -52
rect -16098 -5884 -15960 -5452
rect -15864 -484 -15726 -52
rect -15864 -5884 -15726 -5452
rect -15630 -484 -15492 -52
rect -15630 -5884 -15492 -5452
rect -15396 -484 -15258 -52
rect -15396 -5884 -15258 -5452
rect -15162 -484 -15024 -52
rect -15162 -5884 -15024 -5452
rect -14928 -484 -14790 -52
rect -14928 -5884 -14790 -5452
rect -14694 -484 -14556 -52
rect -14694 -5884 -14556 -5452
rect -14460 -484 -14322 -52
rect -14460 -5884 -14322 -5452
rect -14226 -484 -14088 -52
rect -14226 -5884 -14088 -5452
rect -13992 -484 -13854 -52
rect -13992 -5884 -13854 -5452
rect -13758 -484 -13620 -52
rect -13758 -5884 -13620 -5452
rect -13524 -484 -13386 -52
rect -13524 -5884 -13386 -5452
rect -13290 -484 -13152 -52
rect -13290 -5884 -13152 -5452
rect -13056 -484 -12918 -52
rect -13056 -5884 -12918 -5452
rect -12822 -484 -12684 -52
rect -12822 -5884 -12684 -5452
rect -12588 -484 -12450 -52
rect -12588 -5884 -12450 -5452
rect -12354 -484 -12216 -52
rect -12354 -5884 -12216 -5452
rect -12120 -484 -11982 -52
rect -12120 -5884 -11982 -5452
rect -11886 -484 -11748 -52
rect -11886 -5884 -11748 -5452
rect -11652 -484 -11514 -52
rect -11652 -5884 -11514 -5452
rect -11418 -484 -11280 -52
rect -11418 -5884 -11280 -5452
rect -11184 -484 -11046 -52
rect -11184 -5884 -11046 -5452
rect -10950 -484 -10812 -52
rect -10950 -5884 -10812 -5452
rect -10716 -484 -10578 -52
rect -10716 -5884 -10578 -5452
rect -10482 -484 -10344 -52
rect -10482 -5884 -10344 -5452
rect -10248 -484 -10110 -52
rect -10248 -5884 -10110 -5452
rect -10014 -484 -9876 -52
rect -10014 -5884 -9876 -5452
rect -9780 -484 -9642 -52
rect -9780 -5884 -9642 -5452
rect -9546 -484 -9408 -52
rect -9546 -5884 -9408 -5452
rect -9312 -484 -9174 -52
rect -9312 -5884 -9174 -5452
rect -9078 -484 -8940 -52
rect -9078 -5884 -8940 -5452
rect -8844 -484 -8706 -52
rect -8844 -5884 -8706 -5452
rect -8610 -484 -8472 -52
rect -8610 -5884 -8472 -5452
rect -8376 -484 -8238 -52
rect -8376 -5884 -8238 -5452
rect -8142 -484 -8004 -52
rect -8142 -5884 -8004 -5452
rect -7908 -484 -7770 -52
rect -7908 -5884 -7770 -5452
rect -7674 -484 -7536 -52
rect -7674 -5884 -7536 -5452
rect -7440 -484 -7302 -52
rect -7440 -5884 -7302 -5452
rect -7206 -484 -7068 -52
rect -7206 -5884 -7068 -5452
rect -6972 -484 -6834 -52
rect -6972 -5884 -6834 -5452
rect -6738 -484 -6600 -52
rect -6738 -5884 -6600 -5452
rect -6504 -484 -6366 -52
rect -6504 -5884 -6366 -5452
rect -6270 -484 -6132 -52
rect -6270 -5884 -6132 -5452
rect -6036 -484 -5898 -52
rect -6036 -5884 -5898 -5452
rect -5802 -484 -5664 -52
rect -5802 -5884 -5664 -5452
rect -5568 -484 -5430 -52
rect -5568 -5884 -5430 -5452
rect -5334 -484 -5196 -52
rect -5334 -5884 -5196 -5452
rect -5100 -484 -4962 -52
rect -5100 -5884 -4962 -5452
rect -4866 -484 -4728 -52
rect -4866 -5884 -4728 -5452
rect -4632 -484 -4494 -52
rect -4632 -5884 -4494 -5452
rect -4398 -484 -4260 -52
rect -4398 -5884 -4260 -5452
rect -4164 -484 -4026 -52
rect -4164 -5884 -4026 -5452
rect -3930 -484 -3792 -52
rect -3930 -5884 -3792 -5452
rect -3696 -484 -3558 -52
rect -3696 -5884 -3558 -5452
rect -3462 -484 -3324 -52
rect -3462 -5884 -3324 -5452
rect -3228 -484 -3090 -52
rect -3228 -5884 -3090 -5452
rect -2994 -484 -2856 -52
rect -2994 -5884 -2856 -5452
rect -2760 -484 -2622 -52
rect -2760 -5884 -2622 -5452
rect -2526 -484 -2388 -52
rect -2526 -5884 -2388 -5452
rect -2292 -484 -2154 -52
rect -2292 -5884 -2154 -5452
rect -2058 -484 -1920 -52
rect -2058 -5884 -1920 -5452
rect -1824 -484 -1686 -52
rect -1824 -5884 -1686 -5452
rect -1590 -484 -1452 -52
rect -1590 -5884 -1452 -5452
rect -1356 -484 -1218 -52
rect -1356 -5884 -1218 -5452
rect -1122 -484 -984 -52
rect -1122 -5884 -984 -5452
rect -888 -484 -750 -52
rect -888 -5884 -750 -5452
rect -654 -484 -516 -52
rect -654 -5884 -516 -5452
rect -420 -484 -282 -52
rect -420 -5884 -282 -5452
rect -186 -484 -48 -52
rect -186 -5884 -48 -5452
rect 48 -484 186 -52
rect 48 -5884 186 -5452
rect 282 -484 420 -52
rect 282 -5884 420 -5452
rect 516 -484 654 -52
rect 516 -5884 654 -5452
rect 750 -484 888 -52
rect 750 -5884 888 -5452
rect 984 -484 1122 -52
rect 984 -5884 1122 -5452
rect 1218 -484 1356 -52
rect 1218 -5884 1356 -5452
rect 1452 -484 1590 -52
rect 1452 -5884 1590 -5452
rect 1686 -484 1824 -52
rect 1686 -5884 1824 -5452
rect 1920 -484 2058 -52
rect 1920 -5884 2058 -5452
rect 2154 -484 2292 -52
rect 2154 -5884 2292 -5452
rect 2388 -484 2526 -52
rect 2388 -5884 2526 -5452
rect 2622 -484 2760 -52
rect 2622 -5884 2760 -5452
rect 2856 -484 2994 -52
rect 2856 -5884 2994 -5452
rect 3090 -484 3228 -52
rect 3090 -5884 3228 -5452
rect 3324 -484 3462 -52
rect 3324 -5884 3462 -5452
rect 3558 -484 3696 -52
rect 3558 -5884 3696 -5452
rect 3792 -484 3930 -52
rect 3792 -5884 3930 -5452
rect 4026 -484 4164 -52
rect 4026 -5884 4164 -5452
rect 4260 -484 4398 -52
rect 4260 -5884 4398 -5452
rect 4494 -484 4632 -52
rect 4494 -5884 4632 -5452
rect 4728 -484 4866 -52
rect 4728 -5884 4866 -5452
rect 4962 -484 5100 -52
rect 4962 -5884 5100 -5452
rect 5196 -484 5334 -52
rect 5196 -5884 5334 -5452
rect 5430 -484 5568 -52
rect 5430 -5884 5568 -5452
rect 5664 -484 5802 -52
rect 5664 -5884 5802 -5452
rect 5898 -484 6036 -52
rect 5898 -5884 6036 -5452
rect 6132 -484 6270 -52
rect 6132 -5884 6270 -5452
rect 6366 -484 6504 -52
rect 6366 -5884 6504 -5452
rect 6600 -484 6738 -52
rect 6600 -5884 6738 -5452
rect 6834 -484 6972 -52
rect 6834 -5884 6972 -5452
rect 7068 -484 7206 -52
rect 7068 -5884 7206 -5452
rect 7302 -484 7440 -52
rect 7302 -5884 7440 -5452
rect 7536 -484 7674 -52
rect 7536 -5884 7674 -5452
rect 7770 -484 7908 -52
rect 7770 -5884 7908 -5452
rect 8004 -484 8142 -52
rect 8004 -5884 8142 -5452
rect 8238 -484 8376 -52
rect 8238 -5884 8376 -5452
rect 8472 -484 8610 -52
rect 8472 -5884 8610 -5452
rect 8706 -484 8844 -52
rect 8706 -5884 8844 -5452
rect 8940 -484 9078 -52
rect 8940 -5884 9078 -5452
rect 9174 -484 9312 -52
rect 9174 -5884 9312 -5452
rect 9408 -484 9546 -52
rect 9408 -5884 9546 -5452
rect 9642 -484 9780 -52
rect 9642 -5884 9780 -5452
rect 9876 -484 10014 -52
rect 9876 -5884 10014 -5452
rect 10110 -484 10248 -52
rect 10110 -5884 10248 -5452
rect 10344 -484 10482 -52
rect 10344 -5884 10482 -5452
rect 10578 -484 10716 -52
rect 10578 -5884 10716 -5452
rect 10812 -484 10950 -52
rect 10812 -5884 10950 -5452
rect 11046 -484 11184 -52
rect 11046 -5884 11184 -5452
rect 11280 -484 11418 -52
rect 11280 -5884 11418 -5452
rect 11514 -484 11652 -52
rect 11514 -5884 11652 -5452
rect 11748 -484 11886 -52
rect 11748 -5884 11886 -5452
rect 11982 -484 12120 -52
rect 11982 -5884 12120 -5452
rect 12216 -484 12354 -52
rect 12216 -5884 12354 -5452
rect 12450 -484 12588 -52
rect 12450 -5884 12588 -5452
rect 12684 -484 12822 -52
rect 12684 -5884 12822 -5452
rect 12918 -484 13056 -52
rect 12918 -5884 13056 -5452
rect 13152 -484 13290 -52
rect 13152 -5884 13290 -5452
rect 13386 -484 13524 -52
rect 13386 -5884 13524 -5452
rect 13620 -484 13758 -52
rect 13620 -5884 13758 -5452
rect 13854 -484 13992 -52
rect 13854 -5884 13992 -5452
rect 14088 -484 14226 -52
rect 14088 -5884 14226 -5452
rect 14322 -484 14460 -52
rect 14322 -5884 14460 -5452
rect 14556 -484 14694 -52
rect 14556 -5884 14694 -5452
rect 14790 -484 14928 -52
rect 14790 -5884 14928 -5452
rect 15024 -484 15162 -52
rect 15024 -5884 15162 -5452
rect 15258 -484 15396 -52
rect 15258 -5884 15396 -5452
rect 15492 -484 15630 -52
rect 15492 -5884 15630 -5452
rect 15726 -484 15864 -52
rect 15726 -5884 15864 -5452
rect 15960 -484 16098 -52
rect 15960 -5884 16098 -5452
rect 16194 -484 16332 -52
rect 16194 -5884 16332 -5452
rect 16428 -484 16566 -52
rect 16428 -5884 16566 -5452
rect 16662 -484 16800 -52
rect 16662 -5884 16800 -5452
rect 16896 -484 17034 -52
rect 16896 -5884 17034 -5452
rect 17130 -484 17268 -52
rect 17130 -5884 17268 -5452
rect 17364 -484 17502 -52
rect 17364 -5884 17502 -5452
rect 17598 -484 17736 -52
rect 17598 -5884 17736 -5452
rect 17832 -484 17970 -52
rect 17832 -5884 17970 -5452
rect 18066 -484 18204 -52
rect 18066 -5884 18204 -5452
rect 18300 -484 18438 -52
rect 18300 -5884 18438 -5452
rect 18534 -484 18672 -52
rect 18534 -5884 18672 -5452
rect 18768 -484 18906 -52
rect 18768 -5884 18906 -5452
rect 19002 -484 19140 -52
rect 19002 -5884 19140 -5452
rect 19236 -484 19374 -52
rect 19236 -5884 19374 -5452
rect 19470 -484 19608 -52
rect 19470 -5884 19608 -5452
rect 19704 -484 19842 -52
rect 19704 -5884 19842 -5452
rect 19938 -484 20076 -52
rect 19938 -5884 20076 -5452
rect 20172 -484 20310 -52
rect 20172 -5884 20310 -5452
rect 20406 -484 20544 -52
rect 20406 -5884 20544 -5452
rect 20640 -484 20778 -52
rect 20640 -5884 20778 -5452
rect 20874 -484 21012 -52
rect 20874 -5884 21012 -5452
rect 21108 -484 21246 -52
rect 21108 -5884 21246 -5452
rect 21342 -484 21480 -52
rect 21342 -5884 21480 -5452
rect 21576 -484 21714 -52
rect 21576 -5884 21714 -5452
rect 21810 -484 21948 -52
rect 21810 -5884 21948 -5452
rect 22044 -484 22182 -52
rect 22044 -5884 22182 -5452
rect 22278 -484 22416 -52
rect 22278 -5884 22416 -5452
rect 22512 -484 22650 -52
rect 22512 -5884 22650 -5452
rect 22746 -484 22884 -52
rect 22746 -5884 22884 -5452
rect 22980 -484 23118 -52
rect 22980 -5884 23118 -5452
rect 23214 -484 23352 -52
rect 23214 -5884 23352 -5452
rect 23448 -484 23586 -52
rect 23448 -5884 23586 -5452
rect 23682 -484 23820 -52
rect 23682 -5884 23820 -5452
rect 23916 -484 24054 -52
rect 23916 -5884 24054 -5452
rect 24150 -484 24288 -52
rect 24150 -5884 24288 -5452
rect 24384 -484 24522 -52
rect 24384 -5884 24522 -5452
rect 24618 -484 24756 -52
rect 24618 -5884 24756 -5452
rect 24852 -484 24990 -52
rect 24852 -5884 24990 -5452
rect 25086 -484 25224 -52
rect 25086 -5884 25224 -5452
rect 25320 -484 25458 -52
rect 25320 -5884 25458 -5452
rect 25554 -484 25692 -52
rect 25554 -5884 25692 -5452
rect 25788 -484 25926 -52
rect 25788 -5884 25926 -5452
rect 26022 -484 26160 -52
rect 26022 -5884 26160 -5452
rect 26256 -484 26394 -52
rect 26256 -5884 26394 -5452
rect 26490 -484 26628 -52
rect 26490 -5884 26628 -5452
rect 26724 -484 26862 -52
rect 26724 -5884 26862 -5452
rect 26958 -484 27096 -52
rect 26958 -5884 27096 -5452
rect 27192 -484 27330 -52
rect 27192 -5884 27330 -5452
rect 27426 -484 27564 -52
rect 27426 -5884 27564 -5452
rect 27660 -484 27798 -52
rect 27660 -5884 27798 -5452
rect 27894 -484 28032 -52
rect 27894 -5884 28032 -5452
rect 28128 -484 28266 -52
rect 28128 -5884 28266 -5452
rect 28362 -484 28500 -52
rect 28362 -5884 28500 -5452
rect 28596 -484 28734 -52
rect 28596 -5884 28734 -5452
rect 28830 -484 28968 -52
rect 28830 -5884 28968 -5452
rect 29064 -484 29202 -52
rect 29064 -5884 29202 -5452
rect 29298 -484 29436 -52
rect 29298 -5884 29436 -5452
rect 29532 -484 29670 -52
rect 29532 -5884 29670 -5452
rect 29766 -484 29904 -52
rect 29766 -5884 29904 -5452
<< ppolyres >>
rect -29904 484 -29766 5452
rect -29670 484 -29532 5452
rect -29436 484 -29298 5452
rect -29202 484 -29064 5452
rect -28968 484 -28830 5452
rect -28734 484 -28596 5452
rect -28500 484 -28362 5452
rect -28266 484 -28128 5452
rect -28032 484 -27894 5452
rect -27798 484 -27660 5452
rect -27564 484 -27426 5452
rect -27330 484 -27192 5452
rect -27096 484 -26958 5452
rect -26862 484 -26724 5452
rect -26628 484 -26490 5452
rect -26394 484 -26256 5452
rect -26160 484 -26022 5452
rect -25926 484 -25788 5452
rect -25692 484 -25554 5452
rect -25458 484 -25320 5452
rect -25224 484 -25086 5452
rect -24990 484 -24852 5452
rect -24756 484 -24618 5452
rect -24522 484 -24384 5452
rect -24288 484 -24150 5452
rect -24054 484 -23916 5452
rect -23820 484 -23682 5452
rect -23586 484 -23448 5452
rect -23352 484 -23214 5452
rect -23118 484 -22980 5452
rect -22884 484 -22746 5452
rect -22650 484 -22512 5452
rect -22416 484 -22278 5452
rect -22182 484 -22044 5452
rect -21948 484 -21810 5452
rect -21714 484 -21576 5452
rect -21480 484 -21342 5452
rect -21246 484 -21108 5452
rect -21012 484 -20874 5452
rect -20778 484 -20640 5452
rect -20544 484 -20406 5452
rect -20310 484 -20172 5452
rect -20076 484 -19938 5452
rect -19842 484 -19704 5452
rect -19608 484 -19470 5452
rect -19374 484 -19236 5452
rect -19140 484 -19002 5452
rect -18906 484 -18768 5452
rect -18672 484 -18534 5452
rect -18438 484 -18300 5452
rect -18204 484 -18066 5452
rect -17970 484 -17832 5452
rect -17736 484 -17598 5452
rect -17502 484 -17364 5452
rect -17268 484 -17130 5452
rect -17034 484 -16896 5452
rect -16800 484 -16662 5452
rect -16566 484 -16428 5452
rect -16332 484 -16194 5452
rect -16098 484 -15960 5452
rect -15864 484 -15726 5452
rect -15630 484 -15492 5452
rect -15396 484 -15258 5452
rect -15162 484 -15024 5452
rect -14928 484 -14790 5452
rect -14694 484 -14556 5452
rect -14460 484 -14322 5452
rect -14226 484 -14088 5452
rect -13992 484 -13854 5452
rect -13758 484 -13620 5452
rect -13524 484 -13386 5452
rect -13290 484 -13152 5452
rect -13056 484 -12918 5452
rect -12822 484 -12684 5452
rect -12588 484 -12450 5452
rect -12354 484 -12216 5452
rect -12120 484 -11982 5452
rect -11886 484 -11748 5452
rect -11652 484 -11514 5452
rect -11418 484 -11280 5452
rect -11184 484 -11046 5452
rect -10950 484 -10812 5452
rect -10716 484 -10578 5452
rect -10482 484 -10344 5452
rect -10248 484 -10110 5452
rect -10014 484 -9876 5452
rect -9780 484 -9642 5452
rect -9546 484 -9408 5452
rect -9312 484 -9174 5452
rect -9078 484 -8940 5452
rect -8844 484 -8706 5452
rect -8610 484 -8472 5452
rect -8376 484 -8238 5452
rect -8142 484 -8004 5452
rect -7908 484 -7770 5452
rect -7674 484 -7536 5452
rect -7440 484 -7302 5452
rect -7206 484 -7068 5452
rect -6972 484 -6834 5452
rect -6738 484 -6600 5452
rect -6504 484 -6366 5452
rect -6270 484 -6132 5452
rect -6036 484 -5898 5452
rect -5802 484 -5664 5452
rect -5568 484 -5430 5452
rect -5334 484 -5196 5452
rect -5100 484 -4962 5452
rect -4866 484 -4728 5452
rect -4632 484 -4494 5452
rect -4398 484 -4260 5452
rect -4164 484 -4026 5452
rect -3930 484 -3792 5452
rect -3696 484 -3558 5452
rect -3462 484 -3324 5452
rect -3228 484 -3090 5452
rect -2994 484 -2856 5452
rect -2760 484 -2622 5452
rect -2526 484 -2388 5452
rect -2292 484 -2154 5452
rect -2058 484 -1920 5452
rect -1824 484 -1686 5452
rect -1590 484 -1452 5452
rect -1356 484 -1218 5452
rect -1122 484 -984 5452
rect -888 484 -750 5452
rect -654 484 -516 5452
rect -420 484 -282 5452
rect -186 484 -48 5452
rect 48 484 186 5452
rect 282 484 420 5452
rect 516 484 654 5452
rect 750 484 888 5452
rect 984 484 1122 5452
rect 1218 484 1356 5452
rect 1452 484 1590 5452
rect 1686 484 1824 5452
rect 1920 484 2058 5452
rect 2154 484 2292 5452
rect 2388 484 2526 5452
rect 2622 484 2760 5452
rect 2856 484 2994 5452
rect 3090 484 3228 5452
rect 3324 484 3462 5452
rect 3558 484 3696 5452
rect 3792 484 3930 5452
rect 4026 484 4164 5452
rect 4260 484 4398 5452
rect 4494 484 4632 5452
rect 4728 484 4866 5452
rect 4962 484 5100 5452
rect 5196 484 5334 5452
rect 5430 484 5568 5452
rect 5664 484 5802 5452
rect 5898 484 6036 5452
rect 6132 484 6270 5452
rect 6366 484 6504 5452
rect 6600 484 6738 5452
rect 6834 484 6972 5452
rect 7068 484 7206 5452
rect 7302 484 7440 5452
rect 7536 484 7674 5452
rect 7770 484 7908 5452
rect 8004 484 8142 5452
rect 8238 484 8376 5452
rect 8472 484 8610 5452
rect 8706 484 8844 5452
rect 8940 484 9078 5452
rect 9174 484 9312 5452
rect 9408 484 9546 5452
rect 9642 484 9780 5452
rect 9876 484 10014 5452
rect 10110 484 10248 5452
rect 10344 484 10482 5452
rect 10578 484 10716 5452
rect 10812 484 10950 5452
rect 11046 484 11184 5452
rect 11280 484 11418 5452
rect 11514 484 11652 5452
rect 11748 484 11886 5452
rect 11982 484 12120 5452
rect 12216 484 12354 5452
rect 12450 484 12588 5452
rect 12684 484 12822 5452
rect 12918 484 13056 5452
rect 13152 484 13290 5452
rect 13386 484 13524 5452
rect 13620 484 13758 5452
rect 13854 484 13992 5452
rect 14088 484 14226 5452
rect 14322 484 14460 5452
rect 14556 484 14694 5452
rect 14790 484 14928 5452
rect 15024 484 15162 5452
rect 15258 484 15396 5452
rect 15492 484 15630 5452
rect 15726 484 15864 5452
rect 15960 484 16098 5452
rect 16194 484 16332 5452
rect 16428 484 16566 5452
rect 16662 484 16800 5452
rect 16896 484 17034 5452
rect 17130 484 17268 5452
rect 17364 484 17502 5452
rect 17598 484 17736 5452
rect 17832 484 17970 5452
rect 18066 484 18204 5452
rect 18300 484 18438 5452
rect 18534 484 18672 5452
rect 18768 484 18906 5452
rect 19002 484 19140 5452
rect 19236 484 19374 5452
rect 19470 484 19608 5452
rect 19704 484 19842 5452
rect 19938 484 20076 5452
rect 20172 484 20310 5452
rect 20406 484 20544 5452
rect 20640 484 20778 5452
rect 20874 484 21012 5452
rect 21108 484 21246 5452
rect 21342 484 21480 5452
rect 21576 484 21714 5452
rect 21810 484 21948 5452
rect 22044 484 22182 5452
rect 22278 484 22416 5452
rect 22512 484 22650 5452
rect 22746 484 22884 5452
rect 22980 484 23118 5452
rect 23214 484 23352 5452
rect 23448 484 23586 5452
rect 23682 484 23820 5452
rect 23916 484 24054 5452
rect 24150 484 24288 5452
rect 24384 484 24522 5452
rect 24618 484 24756 5452
rect 24852 484 24990 5452
rect 25086 484 25224 5452
rect 25320 484 25458 5452
rect 25554 484 25692 5452
rect 25788 484 25926 5452
rect 26022 484 26160 5452
rect 26256 484 26394 5452
rect 26490 484 26628 5452
rect 26724 484 26862 5452
rect 26958 484 27096 5452
rect 27192 484 27330 5452
rect 27426 484 27564 5452
rect 27660 484 27798 5452
rect 27894 484 28032 5452
rect 28128 484 28266 5452
rect 28362 484 28500 5452
rect 28596 484 28734 5452
rect 28830 484 28968 5452
rect 29064 484 29202 5452
rect 29298 484 29436 5452
rect 29532 484 29670 5452
rect 29766 484 29904 5452
rect -29904 -5452 -29766 -484
rect -29670 -5452 -29532 -484
rect -29436 -5452 -29298 -484
rect -29202 -5452 -29064 -484
rect -28968 -5452 -28830 -484
rect -28734 -5452 -28596 -484
rect -28500 -5452 -28362 -484
rect -28266 -5452 -28128 -484
rect -28032 -5452 -27894 -484
rect -27798 -5452 -27660 -484
rect -27564 -5452 -27426 -484
rect -27330 -5452 -27192 -484
rect -27096 -5452 -26958 -484
rect -26862 -5452 -26724 -484
rect -26628 -5452 -26490 -484
rect -26394 -5452 -26256 -484
rect -26160 -5452 -26022 -484
rect -25926 -5452 -25788 -484
rect -25692 -5452 -25554 -484
rect -25458 -5452 -25320 -484
rect -25224 -5452 -25086 -484
rect -24990 -5452 -24852 -484
rect -24756 -5452 -24618 -484
rect -24522 -5452 -24384 -484
rect -24288 -5452 -24150 -484
rect -24054 -5452 -23916 -484
rect -23820 -5452 -23682 -484
rect -23586 -5452 -23448 -484
rect -23352 -5452 -23214 -484
rect -23118 -5452 -22980 -484
rect -22884 -5452 -22746 -484
rect -22650 -5452 -22512 -484
rect -22416 -5452 -22278 -484
rect -22182 -5452 -22044 -484
rect -21948 -5452 -21810 -484
rect -21714 -5452 -21576 -484
rect -21480 -5452 -21342 -484
rect -21246 -5452 -21108 -484
rect -21012 -5452 -20874 -484
rect -20778 -5452 -20640 -484
rect -20544 -5452 -20406 -484
rect -20310 -5452 -20172 -484
rect -20076 -5452 -19938 -484
rect -19842 -5452 -19704 -484
rect -19608 -5452 -19470 -484
rect -19374 -5452 -19236 -484
rect -19140 -5452 -19002 -484
rect -18906 -5452 -18768 -484
rect -18672 -5452 -18534 -484
rect -18438 -5452 -18300 -484
rect -18204 -5452 -18066 -484
rect -17970 -5452 -17832 -484
rect -17736 -5452 -17598 -484
rect -17502 -5452 -17364 -484
rect -17268 -5452 -17130 -484
rect -17034 -5452 -16896 -484
rect -16800 -5452 -16662 -484
rect -16566 -5452 -16428 -484
rect -16332 -5452 -16194 -484
rect -16098 -5452 -15960 -484
rect -15864 -5452 -15726 -484
rect -15630 -5452 -15492 -484
rect -15396 -5452 -15258 -484
rect -15162 -5452 -15024 -484
rect -14928 -5452 -14790 -484
rect -14694 -5452 -14556 -484
rect -14460 -5452 -14322 -484
rect -14226 -5452 -14088 -484
rect -13992 -5452 -13854 -484
rect -13758 -5452 -13620 -484
rect -13524 -5452 -13386 -484
rect -13290 -5452 -13152 -484
rect -13056 -5452 -12918 -484
rect -12822 -5452 -12684 -484
rect -12588 -5452 -12450 -484
rect -12354 -5452 -12216 -484
rect -12120 -5452 -11982 -484
rect -11886 -5452 -11748 -484
rect -11652 -5452 -11514 -484
rect -11418 -5452 -11280 -484
rect -11184 -5452 -11046 -484
rect -10950 -5452 -10812 -484
rect -10716 -5452 -10578 -484
rect -10482 -5452 -10344 -484
rect -10248 -5452 -10110 -484
rect -10014 -5452 -9876 -484
rect -9780 -5452 -9642 -484
rect -9546 -5452 -9408 -484
rect -9312 -5452 -9174 -484
rect -9078 -5452 -8940 -484
rect -8844 -5452 -8706 -484
rect -8610 -5452 -8472 -484
rect -8376 -5452 -8238 -484
rect -8142 -5452 -8004 -484
rect -7908 -5452 -7770 -484
rect -7674 -5452 -7536 -484
rect -7440 -5452 -7302 -484
rect -7206 -5452 -7068 -484
rect -6972 -5452 -6834 -484
rect -6738 -5452 -6600 -484
rect -6504 -5452 -6366 -484
rect -6270 -5452 -6132 -484
rect -6036 -5452 -5898 -484
rect -5802 -5452 -5664 -484
rect -5568 -5452 -5430 -484
rect -5334 -5452 -5196 -484
rect -5100 -5452 -4962 -484
rect -4866 -5452 -4728 -484
rect -4632 -5452 -4494 -484
rect -4398 -5452 -4260 -484
rect -4164 -5452 -4026 -484
rect -3930 -5452 -3792 -484
rect -3696 -5452 -3558 -484
rect -3462 -5452 -3324 -484
rect -3228 -5452 -3090 -484
rect -2994 -5452 -2856 -484
rect -2760 -5452 -2622 -484
rect -2526 -5452 -2388 -484
rect -2292 -5452 -2154 -484
rect -2058 -5452 -1920 -484
rect -1824 -5452 -1686 -484
rect -1590 -5452 -1452 -484
rect -1356 -5452 -1218 -484
rect -1122 -5452 -984 -484
rect -888 -5452 -750 -484
rect -654 -5452 -516 -484
rect -420 -5452 -282 -484
rect -186 -5452 -48 -484
rect 48 -5452 186 -484
rect 282 -5452 420 -484
rect 516 -5452 654 -484
rect 750 -5452 888 -484
rect 984 -5452 1122 -484
rect 1218 -5452 1356 -484
rect 1452 -5452 1590 -484
rect 1686 -5452 1824 -484
rect 1920 -5452 2058 -484
rect 2154 -5452 2292 -484
rect 2388 -5452 2526 -484
rect 2622 -5452 2760 -484
rect 2856 -5452 2994 -484
rect 3090 -5452 3228 -484
rect 3324 -5452 3462 -484
rect 3558 -5452 3696 -484
rect 3792 -5452 3930 -484
rect 4026 -5452 4164 -484
rect 4260 -5452 4398 -484
rect 4494 -5452 4632 -484
rect 4728 -5452 4866 -484
rect 4962 -5452 5100 -484
rect 5196 -5452 5334 -484
rect 5430 -5452 5568 -484
rect 5664 -5452 5802 -484
rect 5898 -5452 6036 -484
rect 6132 -5452 6270 -484
rect 6366 -5452 6504 -484
rect 6600 -5452 6738 -484
rect 6834 -5452 6972 -484
rect 7068 -5452 7206 -484
rect 7302 -5452 7440 -484
rect 7536 -5452 7674 -484
rect 7770 -5452 7908 -484
rect 8004 -5452 8142 -484
rect 8238 -5452 8376 -484
rect 8472 -5452 8610 -484
rect 8706 -5452 8844 -484
rect 8940 -5452 9078 -484
rect 9174 -5452 9312 -484
rect 9408 -5452 9546 -484
rect 9642 -5452 9780 -484
rect 9876 -5452 10014 -484
rect 10110 -5452 10248 -484
rect 10344 -5452 10482 -484
rect 10578 -5452 10716 -484
rect 10812 -5452 10950 -484
rect 11046 -5452 11184 -484
rect 11280 -5452 11418 -484
rect 11514 -5452 11652 -484
rect 11748 -5452 11886 -484
rect 11982 -5452 12120 -484
rect 12216 -5452 12354 -484
rect 12450 -5452 12588 -484
rect 12684 -5452 12822 -484
rect 12918 -5452 13056 -484
rect 13152 -5452 13290 -484
rect 13386 -5452 13524 -484
rect 13620 -5452 13758 -484
rect 13854 -5452 13992 -484
rect 14088 -5452 14226 -484
rect 14322 -5452 14460 -484
rect 14556 -5452 14694 -484
rect 14790 -5452 14928 -484
rect 15024 -5452 15162 -484
rect 15258 -5452 15396 -484
rect 15492 -5452 15630 -484
rect 15726 -5452 15864 -484
rect 15960 -5452 16098 -484
rect 16194 -5452 16332 -484
rect 16428 -5452 16566 -484
rect 16662 -5452 16800 -484
rect 16896 -5452 17034 -484
rect 17130 -5452 17268 -484
rect 17364 -5452 17502 -484
rect 17598 -5452 17736 -484
rect 17832 -5452 17970 -484
rect 18066 -5452 18204 -484
rect 18300 -5452 18438 -484
rect 18534 -5452 18672 -484
rect 18768 -5452 18906 -484
rect 19002 -5452 19140 -484
rect 19236 -5452 19374 -484
rect 19470 -5452 19608 -484
rect 19704 -5452 19842 -484
rect 19938 -5452 20076 -484
rect 20172 -5452 20310 -484
rect 20406 -5452 20544 -484
rect 20640 -5452 20778 -484
rect 20874 -5452 21012 -484
rect 21108 -5452 21246 -484
rect 21342 -5452 21480 -484
rect 21576 -5452 21714 -484
rect 21810 -5452 21948 -484
rect 22044 -5452 22182 -484
rect 22278 -5452 22416 -484
rect 22512 -5452 22650 -484
rect 22746 -5452 22884 -484
rect 22980 -5452 23118 -484
rect 23214 -5452 23352 -484
rect 23448 -5452 23586 -484
rect 23682 -5452 23820 -484
rect 23916 -5452 24054 -484
rect 24150 -5452 24288 -484
rect 24384 -5452 24522 -484
rect 24618 -5452 24756 -484
rect 24852 -5452 24990 -484
rect 25086 -5452 25224 -484
rect 25320 -5452 25458 -484
rect 25554 -5452 25692 -484
rect 25788 -5452 25926 -484
rect 26022 -5452 26160 -484
rect 26256 -5452 26394 -484
rect 26490 -5452 26628 -484
rect 26724 -5452 26862 -484
rect 26958 -5452 27096 -484
rect 27192 -5452 27330 -484
rect 27426 -5452 27564 -484
rect 27660 -5452 27798 -484
rect 27894 -5452 28032 -484
rect 28128 -5452 28266 -484
rect 28362 -5452 28500 -484
rect 28596 -5452 28734 -484
rect 28830 -5452 28968 -484
rect 29064 -5452 29202 -484
rect 29298 -5452 29436 -484
rect 29532 -5452 29670 -484
rect 29766 -5452 29904 -484
<< locali >>
rect -30034 5980 -29938 6014
rect 29938 5980 30034 6014
rect -30034 5918 -30000 5980
rect 30000 5918 30034 5980
rect -30034 -5980 -30000 -5918
rect 30000 -5980 30034 -5918
rect -30034 -6014 -29938 -5980
rect 29938 -6014 30034 -5980
<< viali >>
rect -29888 5469 -29782 5866
rect -29654 5469 -29548 5866
rect -29420 5469 -29314 5866
rect -29186 5469 -29080 5866
rect -28952 5469 -28846 5866
rect -28718 5469 -28612 5866
rect -28484 5469 -28378 5866
rect -28250 5469 -28144 5866
rect -28016 5469 -27910 5866
rect -27782 5469 -27676 5866
rect -27548 5469 -27442 5866
rect -27314 5469 -27208 5866
rect -27080 5469 -26974 5866
rect -26846 5469 -26740 5866
rect -26612 5469 -26506 5866
rect -26378 5469 -26272 5866
rect -26144 5469 -26038 5866
rect -25910 5469 -25804 5866
rect -25676 5469 -25570 5866
rect -25442 5469 -25336 5866
rect -25208 5469 -25102 5866
rect -24974 5469 -24868 5866
rect -24740 5469 -24634 5866
rect -24506 5469 -24400 5866
rect -24272 5469 -24166 5866
rect -24038 5469 -23932 5866
rect -23804 5469 -23698 5866
rect -23570 5469 -23464 5866
rect -23336 5469 -23230 5866
rect -23102 5469 -22996 5866
rect -22868 5469 -22762 5866
rect -22634 5469 -22528 5866
rect -22400 5469 -22294 5866
rect -22166 5469 -22060 5866
rect -21932 5469 -21826 5866
rect -21698 5469 -21592 5866
rect -21464 5469 -21358 5866
rect -21230 5469 -21124 5866
rect -20996 5469 -20890 5866
rect -20762 5469 -20656 5866
rect -20528 5469 -20422 5866
rect -20294 5469 -20188 5866
rect -20060 5469 -19954 5866
rect -19826 5469 -19720 5866
rect -19592 5469 -19486 5866
rect -19358 5469 -19252 5866
rect -19124 5469 -19018 5866
rect -18890 5469 -18784 5866
rect -18656 5469 -18550 5866
rect -18422 5469 -18316 5866
rect -18188 5469 -18082 5866
rect -17954 5469 -17848 5866
rect -17720 5469 -17614 5866
rect -17486 5469 -17380 5866
rect -17252 5469 -17146 5866
rect -17018 5469 -16912 5866
rect -16784 5469 -16678 5866
rect -16550 5469 -16444 5866
rect -16316 5469 -16210 5866
rect -16082 5469 -15976 5866
rect -15848 5469 -15742 5866
rect -15614 5469 -15508 5866
rect -15380 5469 -15274 5866
rect -15146 5469 -15040 5866
rect -14912 5469 -14806 5866
rect -14678 5469 -14572 5866
rect -14444 5469 -14338 5866
rect -14210 5469 -14104 5866
rect -13976 5469 -13870 5866
rect -13742 5469 -13636 5866
rect -13508 5469 -13402 5866
rect -13274 5469 -13168 5866
rect -13040 5469 -12934 5866
rect -12806 5469 -12700 5866
rect -12572 5469 -12466 5866
rect -12338 5469 -12232 5866
rect -12104 5469 -11998 5866
rect -11870 5469 -11764 5866
rect -11636 5469 -11530 5866
rect -11402 5469 -11296 5866
rect -11168 5469 -11062 5866
rect -10934 5469 -10828 5866
rect -10700 5469 -10594 5866
rect -10466 5469 -10360 5866
rect -10232 5469 -10126 5866
rect -9998 5469 -9892 5866
rect -9764 5469 -9658 5866
rect -9530 5469 -9424 5866
rect -9296 5469 -9190 5866
rect -9062 5469 -8956 5866
rect -8828 5469 -8722 5866
rect -8594 5469 -8488 5866
rect -8360 5469 -8254 5866
rect -8126 5469 -8020 5866
rect -7892 5469 -7786 5866
rect -7658 5469 -7552 5866
rect -7424 5469 -7318 5866
rect -7190 5469 -7084 5866
rect -6956 5469 -6850 5866
rect -6722 5469 -6616 5866
rect -6488 5469 -6382 5866
rect -6254 5469 -6148 5866
rect -6020 5469 -5914 5866
rect -5786 5469 -5680 5866
rect -5552 5469 -5446 5866
rect -5318 5469 -5212 5866
rect -5084 5469 -4978 5866
rect -4850 5469 -4744 5866
rect -4616 5469 -4510 5866
rect -4382 5469 -4276 5866
rect -4148 5469 -4042 5866
rect -3914 5469 -3808 5866
rect -3680 5469 -3574 5866
rect -3446 5469 -3340 5866
rect -3212 5469 -3106 5866
rect -2978 5469 -2872 5866
rect -2744 5469 -2638 5866
rect -2510 5469 -2404 5866
rect -2276 5469 -2170 5866
rect -2042 5469 -1936 5866
rect -1808 5469 -1702 5866
rect -1574 5469 -1468 5866
rect -1340 5469 -1234 5866
rect -1106 5469 -1000 5866
rect -872 5469 -766 5866
rect -638 5469 -532 5866
rect -404 5469 -298 5866
rect -170 5469 -64 5866
rect 64 5469 170 5866
rect 298 5469 404 5866
rect 532 5469 638 5866
rect 766 5469 872 5866
rect 1000 5469 1106 5866
rect 1234 5469 1340 5866
rect 1468 5469 1574 5866
rect 1702 5469 1808 5866
rect 1936 5469 2042 5866
rect 2170 5469 2276 5866
rect 2404 5469 2510 5866
rect 2638 5469 2744 5866
rect 2872 5469 2978 5866
rect 3106 5469 3212 5866
rect 3340 5469 3446 5866
rect 3574 5469 3680 5866
rect 3808 5469 3914 5866
rect 4042 5469 4148 5866
rect 4276 5469 4382 5866
rect 4510 5469 4616 5866
rect 4744 5469 4850 5866
rect 4978 5469 5084 5866
rect 5212 5469 5318 5866
rect 5446 5469 5552 5866
rect 5680 5469 5786 5866
rect 5914 5469 6020 5866
rect 6148 5469 6254 5866
rect 6382 5469 6488 5866
rect 6616 5469 6722 5866
rect 6850 5469 6956 5866
rect 7084 5469 7190 5866
rect 7318 5469 7424 5866
rect 7552 5469 7658 5866
rect 7786 5469 7892 5866
rect 8020 5469 8126 5866
rect 8254 5469 8360 5866
rect 8488 5469 8594 5866
rect 8722 5469 8828 5866
rect 8956 5469 9062 5866
rect 9190 5469 9296 5866
rect 9424 5469 9530 5866
rect 9658 5469 9764 5866
rect 9892 5469 9998 5866
rect 10126 5469 10232 5866
rect 10360 5469 10466 5866
rect 10594 5469 10700 5866
rect 10828 5469 10934 5866
rect 11062 5469 11168 5866
rect 11296 5469 11402 5866
rect 11530 5469 11636 5866
rect 11764 5469 11870 5866
rect 11998 5469 12104 5866
rect 12232 5469 12338 5866
rect 12466 5469 12572 5866
rect 12700 5469 12806 5866
rect 12934 5469 13040 5866
rect 13168 5469 13274 5866
rect 13402 5469 13508 5866
rect 13636 5469 13742 5866
rect 13870 5469 13976 5866
rect 14104 5469 14210 5866
rect 14338 5469 14444 5866
rect 14572 5469 14678 5866
rect 14806 5469 14912 5866
rect 15040 5469 15146 5866
rect 15274 5469 15380 5866
rect 15508 5469 15614 5866
rect 15742 5469 15848 5866
rect 15976 5469 16082 5866
rect 16210 5469 16316 5866
rect 16444 5469 16550 5866
rect 16678 5469 16784 5866
rect 16912 5469 17018 5866
rect 17146 5469 17252 5866
rect 17380 5469 17486 5866
rect 17614 5469 17720 5866
rect 17848 5469 17954 5866
rect 18082 5469 18188 5866
rect 18316 5469 18422 5866
rect 18550 5469 18656 5866
rect 18784 5469 18890 5866
rect 19018 5469 19124 5866
rect 19252 5469 19358 5866
rect 19486 5469 19592 5866
rect 19720 5469 19826 5866
rect 19954 5469 20060 5866
rect 20188 5469 20294 5866
rect 20422 5469 20528 5866
rect 20656 5469 20762 5866
rect 20890 5469 20996 5866
rect 21124 5469 21230 5866
rect 21358 5469 21464 5866
rect 21592 5469 21698 5866
rect 21826 5469 21932 5866
rect 22060 5469 22166 5866
rect 22294 5469 22400 5866
rect 22528 5469 22634 5866
rect 22762 5469 22868 5866
rect 22996 5469 23102 5866
rect 23230 5469 23336 5866
rect 23464 5469 23570 5866
rect 23698 5469 23804 5866
rect 23932 5469 24038 5866
rect 24166 5469 24272 5866
rect 24400 5469 24506 5866
rect 24634 5469 24740 5866
rect 24868 5469 24974 5866
rect 25102 5469 25208 5866
rect 25336 5469 25442 5866
rect 25570 5469 25676 5866
rect 25804 5469 25910 5866
rect 26038 5469 26144 5866
rect 26272 5469 26378 5866
rect 26506 5469 26612 5866
rect 26740 5469 26846 5866
rect 26974 5469 27080 5866
rect 27208 5469 27314 5866
rect 27442 5469 27548 5866
rect 27676 5469 27782 5866
rect 27910 5469 28016 5866
rect 28144 5469 28250 5866
rect 28378 5469 28484 5866
rect 28612 5469 28718 5866
rect 28846 5469 28952 5866
rect 29080 5469 29186 5866
rect 29314 5469 29420 5866
rect 29548 5469 29654 5866
rect 29782 5469 29888 5866
rect -29888 70 -29782 467
rect -29654 70 -29548 467
rect -29420 70 -29314 467
rect -29186 70 -29080 467
rect -28952 70 -28846 467
rect -28718 70 -28612 467
rect -28484 70 -28378 467
rect -28250 70 -28144 467
rect -28016 70 -27910 467
rect -27782 70 -27676 467
rect -27548 70 -27442 467
rect -27314 70 -27208 467
rect -27080 70 -26974 467
rect -26846 70 -26740 467
rect -26612 70 -26506 467
rect -26378 70 -26272 467
rect -26144 70 -26038 467
rect -25910 70 -25804 467
rect -25676 70 -25570 467
rect -25442 70 -25336 467
rect -25208 70 -25102 467
rect -24974 70 -24868 467
rect -24740 70 -24634 467
rect -24506 70 -24400 467
rect -24272 70 -24166 467
rect -24038 70 -23932 467
rect -23804 70 -23698 467
rect -23570 70 -23464 467
rect -23336 70 -23230 467
rect -23102 70 -22996 467
rect -22868 70 -22762 467
rect -22634 70 -22528 467
rect -22400 70 -22294 467
rect -22166 70 -22060 467
rect -21932 70 -21826 467
rect -21698 70 -21592 467
rect -21464 70 -21358 467
rect -21230 70 -21124 467
rect -20996 70 -20890 467
rect -20762 70 -20656 467
rect -20528 70 -20422 467
rect -20294 70 -20188 467
rect -20060 70 -19954 467
rect -19826 70 -19720 467
rect -19592 70 -19486 467
rect -19358 70 -19252 467
rect -19124 70 -19018 467
rect -18890 70 -18784 467
rect -18656 70 -18550 467
rect -18422 70 -18316 467
rect -18188 70 -18082 467
rect -17954 70 -17848 467
rect -17720 70 -17614 467
rect -17486 70 -17380 467
rect -17252 70 -17146 467
rect -17018 70 -16912 467
rect -16784 70 -16678 467
rect -16550 70 -16444 467
rect -16316 70 -16210 467
rect -16082 70 -15976 467
rect -15848 70 -15742 467
rect -15614 70 -15508 467
rect -15380 70 -15274 467
rect -15146 70 -15040 467
rect -14912 70 -14806 467
rect -14678 70 -14572 467
rect -14444 70 -14338 467
rect -14210 70 -14104 467
rect -13976 70 -13870 467
rect -13742 70 -13636 467
rect -13508 70 -13402 467
rect -13274 70 -13168 467
rect -13040 70 -12934 467
rect -12806 70 -12700 467
rect -12572 70 -12466 467
rect -12338 70 -12232 467
rect -12104 70 -11998 467
rect -11870 70 -11764 467
rect -11636 70 -11530 467
rect -11402 70 -11296 467
rect -11168 70 -11062 467
rect -10934 70 -10828 467
rect -10700 70 -10594 467
rect -10466 70 -10360 467
rect -10232 70 -10126 467
rect -9998 70 -9892 467
rect -9764 70 -9658 467
rect -9530 70 -9424 467
rect -9296 70 -9190 467
rect -9062 70 -8956 467
rect -8828 70 -8722 467
rect -8594 70 -8488 467
rect -8360 70 -8254 467
rect -8126 70 -8020 467
rect -7892 70 -7786 467
rect -7658 70 -7552 467
rect -7424 70 -7318 467
rect -7190 70 -7084 467
rect -6956 70 -6850 467
rect -6722 70 -6616 467
rect -6488 70 -6382 467
rect -6254 70 -6148 467
rect -6020 70 -5914 467
rect -5786 70 -5680 467
rect -5552 70 -5446 467
rect -5318 70 -5212 467
rect -5084 70 -4978 467
rect -4850 70 -4744 467
rect -4616 70 -4510 467
rect -4382 70 -4276 467
rect -4148 70 -4042 467
rect -3914 70 -3808 467
rect -3680 70 -3574 467
rect -3446 70 -3340 467
rect -3212 70 -3106 467
rect -2978 70 -2872 467
rect -2744 70 -2638 467
rect -2510 70 -2404 467
rect -2276 70 -2170 467
rect -2042 70 -1936 467
rect -1808 70 -1702 467
rect -1574 70 -1468 467
rect -1340 70 -1234 467
rect -1106 70 -1000 467
rect -872 70 -766 467
rect -638 70 -532 467
rect -404 70 -298 467
rect -170 70 -64 467
rect 64 70 170 467
rect 298 70 404 467
rect 532 70 638 467
rect 766 70 872 467
rect 1000 70 1106 467
rect 1234 70 1340 467
rect 1468 70 1574 467
rect 1702 70 1808 467
rect 1936 70 2042 467
rect 2170 70 2276 467
rect 2404 70 2510 467
rect 2638 70 2744 467
rect 2872 70 2978 467
rect 3106 70 3212 467
rect 3340 70 3446 467
rect 3574 70 3680 467
rect 3808 70 3914 467
rect 4042 70 4148 467
rect 4276 70 4382 467
rect 4510 70 4616 467
rect 4744 70 4850 467
rect 4978 70 5084 467
rect 5212 70 5318 467
rect 5446 70 5552 467
rect 5680 70 5786 467
rect 5914 70 6020 467
rect 6148 70 6254 467
rect 6382 70 6488 467
rect 6616 70 6722 467
rect 6850 70 6956 467
rect 7084 70 7190 467
rect 7318 70 7424 467
rect 7552 70 7658 467
rect 7786 70 7892 467
rect 8020 70 8126 467
rect 8254 70 8360 467
rect 8488 70 8594 467
rect 8722 70 8828 467
rect 8956 70 9062 467
rect 9190 70 9296 467
rect 9424 70 9530 467
rect 9658 70 9764 467
rect 9892 70 9998 467
rect 10126 70 10232 467
rect 10360 70 10466 467
rect 10594 70 10700 467
rect 10828 70 10934 467
rect 11062 70 11168 467
rect 11296 70 11402 467
rect 11530 70 11636 467
rect 11764 70 11870 467
rect 11998 70 12104 467
rect 12232 70 12338 467
rect 12466 70 12572 467
rect 12700 70 12806 467
rect 12934 70 13040 467
rect 13168 70 13274 467
rect 13402 70 13508 467
rect 13636 70 13742 467
rect 13870 70 13976 467
rect 14104 70 14210 467
rect 14338 70 14444 467
rect 14572 70 14678 467
rect 14806 70 14912 467
rect 15040 70 15146 467
rect 15274 70 15380 467
rect 15508 70 15614 467
rect 15742 70 15848 467
rect 15976 70 16082 467
rect 16210 70 16316 467
rect 16444 70 16550 467
rect 16678 70 16784 467
rect 16912 70 17018 467
rect 17146 70 17252 467
rect 17380 70 17486 467
rect 17614 70 17720 467
rect 17848 70 17954 467
rect 18082 70 18188 467
rect 18316 70 18422 467
rect 18550 70 18656 467
rect 18784 70 18890 467
rect 19018 70 19124 467
rect 19252 70 19358 467
rect 19486 70 19592 467
rect 19720 70 19826 467
rect 19954 70 20060 467
rect 20188 70 20294 467
rect 20422 70 20528 467
rect 20656 70 20762 467
rect 20890 70 20996 467
rect 21124 70 21230 467
rect 21358 70 21464 467
rect 21592 70 21698 467
rect 21826 70 21932 467
rect 22060 70 22166 467
rect 22294 70 22400 467
rect 22528 70 22634 467
rect 22762 70 22868 467
rect 22996 70 23102 467
rect 23230 70 23336 467
rect 23464 70 23570 467
rect 23698 70 23804 467
rect 23932 70 24038 467
rect 24166 70 24272 467
rect 24400 70 24506 467
rect 24634 70 24740 467
rect 24868 70 24974 467
rect 25102 70 25208 467
rect 25336 70 25442 467
rect 25570 70 25676 467
rect 25804 70 25910 467
rect 26038 70 26144 467
rect 26272 70 26378 467
rect 26506 70 26612 467
rect 26740 70 26846 467
rect 26974 70 27080 467
rect 27208 70 27314 467
rect 27442 70 27548 467
rect 27676 70 27782 467
rect 27910 70 28016 467
rect 28144 70 28250 467
rect 28378 70 28484 467
rect 28612 70 28718 467
rect 28846 70 28952 467
rect 29080 70 29186 467
rect 29314 70 29420 467
rect 29548 70 29654 467
rect 29782 70 29888 467
rect -29888 -467 -29782 -70
rect -29654 -467 -29548 -70
rect -29420 -467 -29314 -70
rect -29186 -467 -29080 -70
rect -28952 -467 -28846 -70
rect -28718 -467 -28612 -70
rect -28484 -467 -28378 -70
rect -28250 -467 -28144 -70
rect -28016 -467 -27910 -70
rect -27782 -467 -27676 -70
rect -27548 -467 -27442 -70
rect -27314 -467 -27208 -70
rect -27080 -467 -26974 -70
rect -26846 -467 -26740 -70
rect -26612 -467 -26506 -70
rect -26378 -467 -26272 -70
rect -26144 -467 -26038 -70
rect -25910 -467 -25804 -70
rect -25676 -467 -25570 -70
rect -25442 -467 -25336 -70
rect -25208 -467 -25102 -70
rect -24974 -467 -24868 -70
rect -24740 -467 -24634 -70
rect -24506 -467 -24400 -70
rect -24272 -467 -24166 -70
rect -24038 -467 -23932 -70
rect -23804 -467 -23698 -70
rect -23570 -467 -23464 -70
rect -23336 -467 -23230 -70
rect -23102 -467 -22996 -70
rect -22868 -467 -22762 -70
rect -22634 -467 -22528 -70
rect -22400 -467 -22294 -70
rect -22166 -467 -22060 -70
rect -21932 -467 -21826 -70
rect -21698 -467 -21592 -70
rect -21464 -467 -21358 -70
rect -21230 -467 -21124 -70
rect -20996 -467 -20890 -70
rect -20762 -467 -20656 -70
rect -20528 -467 -20422 -70
rect -20294 -467 -20188 -70
rect -20060 -467 -19954 -70
rect -19826 -467 -19720 -70
rect -19592 -467 -19486 -70
rect -19358 -467 -19252 -70
rect -19124 -467 -19018 -70
rect -18890 -467 -18784 -70
rect -18656 -467 -18550 -70
rect -18422 -467 -18316 -70
rect -18188 -467 -18082 -70
rect -17954 -467 -17848 -70
rect -17720 -467 -17614 -70
rect -17486 -467 -17380 -70
rect -17252 -467 -17146 -70
rect -17018 -467 -16912 -70
rect -16784 -467 -16678 -70
rect -16550 -467 -16444 -70
rect -16316 -467 -16210 -70
rect -16082 -467 -15976 -70
rect -15848 -467 -15742 -70
rect -15614 -467 -15508 -70
rect -15380 -467 -15274 -70
rect -15146 -467 -15040 -70
rect -14912 -467 -14806 -70
rect -14678 -467 -14572 -70
rect -14444 -467 -14338 -70
rect -14210 -467 -14104 -70
rect -13976 -467 -13870 -70
rect -13742 -467 -13636 -70
rect -13508 -467 -13402 -70
rect -13274 -467 -13168 -70
rect -13040 -467 -12934 -70
rect -12806 -467 -12700 -70
rect -12572 -467 -12466 -70
rect -12338 -467 -12232 -70
rect -12104 -467 -11998 -70
rect -11870 -467 -11764 -70
rect -11636 -467 -11530 -70
rect -11402 -467 -11296 -70
rect -11168 -467 -11062 -70
rect -10934 -467 -10828 -70
rect -10700 -467 -10594 -70
rect -10466 -467 -10360 -70
rect -10232 -467 -10126 -70
rect -9998 -467 -9892 -70
rect -9764 -467 -9658 -70
rect -9530 -467 -9424 -70
rect -9296 -467 -9190 -70
rect -9062 -467 -8956 -70
rect -8828 -467 -8722 -70
rect -8594 -467 -8488 -70
rect -8360 -467 -8254 -70
rect -8126 -467 -8020 -70
rect -7892 -467 -7786 -70
rect -7658 -467 -7552 -70
rect -7424 -467 -7318 -70
rect -7190 -467 -7084 -70
rect -6956 -467 -6850 -70
rect -6722 -467 -6616 -70
rect -6488 -467 -6382 -70
rect -6254 -467 -6148 -70
rect -6020 -467 -5914 -70
rect -5786 -467 -5680 -70
rect -5552 -467 -5446 -70
rect -5318 -467 -5212 -70
rect -5084 -467 -4978 -70
rect -4850 -467 -4744 -70
rect -4616 -467 -4510 -70
rect -4382 -467 -4276 -70
rect -4148 -467 -4042 -70
rect -3914 -467 -3808 -70
rect -3680 -467 -3574 -70
rect -3446 -467 -3340 -70
rect -3212 -467 -3106 -70
rect -2978 -467 -2872 -70
rect -2744 -467 -2638 -70
rect -2510 -467 -2404 -70
rect -2276 -467 -2170 -70
rect -2042 -467 -1936 -70
rect -1808 -467 -1702 -70
rect -1574 -467 -1468 -70
rect -1340 -467 -1234 -70
rect -1106 -467 -1000 -70
rect -872 -467 -766 -70
rect -638 -467 -532 -70
rect -404 -467 -298 -70
rect -170 -467 -64 -70
rect 64 -467 170 -70
rect 298 -467 404 -70
rect 532 -467 638 -70
rect 766 -467 872 -70
rect 1000 -467 1106 -70
rect 1234 -467 1340 -70
rect 1468 -467 1574 -70
rect 1702 -467 1808 -70
rect 1936 -467 2042 -70
rect 2170 -467 2276 -70
rect 2404 -467 2510 -70
rect 2638 -467 2744 -70
rect 2872 -467 2978 -70
rect 3106 -467 3212 -70
rect 3340 -467 3446 -70
rect 3574 -467 3680 -70
rect 3808 -467 3914 -70
rect 4042 -467 4148 -70
rect 4276 -467 4382 -70
rect 4510 -467 4616 -70
rect 4744 -467 4850 -70
rect 4978 -467 5084 -70
rect 5212 -467 5318 -70
rect 5446 -467 5552 -70
rect 5680 -467 5786 -70
rect 5914 -467 6020 -70
rect 6148 -467 6254 -70
rect 6382 -467 6488 -70
rect 6616 -467 6722 -70
rect 6850 -467 6956 -70
rect 7084 -467 7190 -70
rect 7318 -467 7424 -70
rect 7552 -467 7658 -70
rect 7786 -467 7892 -70
rect 8020 -467 8126 -70
rect 8254 -467 8360 -70
rect 8488 -467 8594 -70
rect 8722 -467 8828 -70
rect 8956 -467 9062 -70
rect 9190 -467 9296 -70
rect 9424 -467 9530 -70
rect 9658 -467 9764 -70
rect 9892 -467 9998 -70
rect 10126 -467 10232 -70
rect 10360 -467 10466 -70
rect 10594 -467 10700 -70
rect 10828 -467 10934 -70
rect 11062 -467 11168 -70
rect 11296 -467 11402 -70
rect 11530 -467 11636 -70
rect 11764 -467 11870 -70
rect 11998 -467 12104 -70
rect 12232 -467 12338 -70
rect 12466 -467 12572 -70
rect 12700 -467 12806 -70
rect 12934 -467 13040 -70
rect 13168 -467 13274 -70
rect 13402 -467 13508 -70
rect 13636 -467 13742 -70
rect 13870 -467 13976 -70
rect 14104 -467 14210 -70
rect 14338 -467 14444 -70
rect 14572 -467 14678 -70
rect 14806 -467 14912 -70
rect 15040 -467 15146 -70
rect 15274 -467 15380 -70
rect 15508 -467 15614 -70
rect 15742 -467 15848 -70
rect 15976 -467 16082 -70
rect 16210 -467 16316 -70
rect 16444 -467 16550 -70
rect 16678 -467 16784 -70
rect 16912 -467 17018 -70
rect 17146 -467 17252 -70
rect 17380 -467 17486 -70
rect 17614 -467 17720 -70
rect 17848 -467 17954 -70
rect 18082 -467 18188 -70
rect 18316 -467 18422 -70
rect 18550 -467 18656 -70
rect 18784 -467 18890 -70
rect 19018 -467 19124 -70
rect 19252 -467 19358 -70
rect 19486 -467 19592 -70
rect 19720 -467 19826 -70
rect 19954 -467 20060 -70
rect 20188 -467 20294 -70
rect 20422 -467 20528 -70
rect 20656 -467 20762 -70
rect 20890 -467 20996 -70
rect 21124 -467 21230 -70
rect 21358 -467 21464 -70
rect 21592 -467 21698 -70
rect 21826 -467 21932 -70
rect 22060 -467 22166 -70
rect 22294 -467 22400 -70
rect 22528 -467 22634 -70
rect 22762 -467 22868 -70
rect 22996 -467 23102 -70
rect 23230 -467 23336 -70
rect 23464 -467 23570 -70
rect 23698 -467 23804 -70
rect 23932 -467 24038 -70
rect 24166 -467 24272 -70
rect 24400 -467 24506 -70
rect 24634 -467 24740 -70
rect 24868 -467 24974 -70
rect 25102 -467 25208 -70
rect 25336 -467 25442 -70
rect 25570 -467 25676 -70
rect 25804 -467 25910 -70
rect 26038 -467 26144 -70
rect 26272 -467 26378 -70
rect 26506 -467 26612 -70
rect 26740 -467 26846 -70
rect 26974 -467 27080 -70
rect 27208 -467 27314 -70
rect 27442 -467 27548 -70
rect 27676 -467 27782 -70
rect 27910 -467 28016 -70
rect 28144 -467 28250 -70
rect 28378 -467 28484 -70
rect 28612 -467 28718 -70
rect 28846 -467 28952 -70
rect 29080 -467 29186 -70
rect 29314 -467 29420 -70
rect 29548 -467 29654 -70
rect 29782 -467 29888 -70
rect -29888 -5866 -29782 -5469
rect -29654 -5866 -29548 -5469
rect -29420 -5866 -29314 -5469
rect -29186 -5866 -29080 -5469
rect -28952 -5866 -28846 -5469
rect -28718 -5866 -28612 -5469
rect -28484 -5866 -28378 -5469
rect -28250 -5866 -28144 -5469
rect -28016 -5866 -27910 -5469
rect -27782 -5866 -27676 -5469
rect -27548 -5866 -27442 -5469
rect -27314 -5866 -27208 -5469
rect -27080 -5866 -26974 -5469
rect -26846 -5866 -26740 -5469
rect -26612 -5866 -26506 -5469
rect -26378 -5866 -26272 -5469
rect -26144 -5866 -26038 -5469
rect -25910 -5866 -25804 -5469
rect -25676 -5866 -25570 -5469
rect -25442 -5866 -25336 -5469
rect -25208 -5866 -25102 -5469
rect -24974 -5866 -24868 -5469
rect -24740 -5866 -24634 -5469
rect -24506 -5866 -24400 -5469
rect -24272 -5866 -24166 -5469
rect -24038 -5866 -23932 -5469
rect -23804 -5866 -23698 -5469
rect -23570 -5866 -23464 -5469
rect -23336 -5866 -23230 -5469
rect -23102 -5866 -22996 -5469
rect -22868 -5866 -22762 -5469
rect -22634 -5866 -22528 -5469
rect -22400 -5866 -22294 -5469
rect -22166 -5866 -22060 -5469
rect -21932 -5866 -21826 -5469
rect -21698 -5866 -21592 -5469
rect -21464 -5866 -21358 -5469
rect -21230 -5866 -21124 -5469
rect -20996 -5866 -20890 -5469
rect -20762 -5866 -20656 -5469
rect -20528 -5866 -20422 -5469
rect -20294 -5866 -20188 -5469
rect -20060 -5866 -19954 -5469
rect -19826 -5866 -19720 -5469
rect -19592 -5866 -19486 -5469
rect -19358 -5866 -19252 -5469
rect -19124 -5866 -19018 -5469
rect -18890 -5866 -18784 -5469
rect -18656 -5866 -18550 -5469
rect -18422 -5866 -18316 -5469
rect -18188 -5866 -18082 -5469
rect -17954 -5866 -17848 -5469
rect -17720 -5866 -17614 -5469
rect -17486 -5866 -17380 -5469
rect -17252 -5866 -17146 -5469
rect -17018 -5866 -16912 -5469
rect -16784 -5866 -16678 -5469
rect -16550 -5866 -16444 -5469
rect -16316 -5866 -16210 -5469
rect -16082 -5866 -15976 -5469
rect -15848 -5866 -15742 -5469
rect -15614 -5866 -15508 -5469
rect -15380 -5866 -15274 -5469
rect -15146 -5866 -15040 -5469
rect -14912 -5866 -14806 -5469
rect -14678 -5866 -14572 -5469
rect -14444 -5866 -14338 -5469
rect -14210 -5866 -14104 -5469
rect -13976 -5866 -13870 -5469
rect -13742 -5866 -13636 -5469
rect -13508 -5866 -13402 -5469
rect -13274 -5866 -13168 -5469
rect -13040 -5866 -12934 -5469
rect -12806 -5866 -12700 -5469
rect -12572 -5866 -12466 -5469
rect -12338 -5866 -12232 -5469
rect -12104 -5866 -11998 -5469
rect -11870 -5866 -11764 -5469
rect -11636 -5866 -11530 -5469
rect -11402 -5866 -11296 -5469
rect -11168 -5866 -11062 -5469
rect -10934 -5866 -10828 -5469
rect -10700 -5866 -10594 -5469
rect -10466 -5866 -10360 -5469
rect -10232 -5866 -10126 -5469
rect -9998 -5866 -9892 -5469
rect -9764 -5866 -9658 -5469
rect -9530 -5866 -9424 -5469
rect -9296 -5866 -9190 -5469
rect -9062 -5866 -8956 -5469
rect -8828 -5866 -8722 -5469
rect -8594 -5866 -8488 -5469
rect -8360 -5866 -8254 -5469
rect -8126 -5866 -8020 -5469
rect -7892 -5866 -7786 -5469
rect -7658 -5866 -7552 -5469
rect -7424 -5866 -7318 -5469
rect -7190 -5866 -7084 -5469
rect -6956 -5866 -6850 -5469
rect -6722 -5866 -6616 -5469
rect -6488 -5866 -6382 -5469
rect -6254 -5866 -6148 -5469
rect -6020 -5866 -5914 -5469
rect -5786 -5866 -5680 -5469
rect -5552 -5866 -5446 -5469
rect -5318 -5866 -5212 -5469
rect -5084 -5866 -4978 -5469
rect -4850 -5866 -4744 -5469
rect -4616 -5866 -4510 -5469
rect -4382 -5866 -4276 -5469
rect -4148 -5866 -4042 -5469
rect -3914 -5866 -3808 -5469
rect -3680 -5866 -3574 -5469
rect -3446 -5866 -3340 -5469
rect -3212 -5866 -3106 -5469
rect -2978 -5866 -2872 -5469
rect -2744 -5866 -2638 -5469
rect -2510 -5866 -2404 -5469
rect -2276 -5866 -2170 -5469
rect -2042 -5866 -1936 -5469
rect -1808 -5866 -1702 -5469
rect -1574 -5866 -1468 -5469
rect -1340 -5866 -1234 -5469
rect -1106 -5866 -1000 -5469
rect -872 -5866 -766 -5469
rect -638 -5866 -532 -5469
rect -404 -5866 -298 -5469
rect -170 -5866 -64 -5469
rect 64 -5866 170 -5469
rect 298 -5866 404 -5469
rect 532 -5866 638 -5469
rect 766 -5866 872 -5469
rect 1000 -5866 1106 -5469
rect 1234 -5866 1340 -5469
rect 1468 -5866 1574 -5469
rect 1702 -5866 1808 -5469
rect 1936 -5866 2042 -5469
rect 2170 -5866 2276 -5469
rect 2404 -5866 2510 -5469
rect 2638 -5866 2744 -5469
rect 2872 -5866 2978 -5469
rect 3106 -5866 3212 -5469
rect 3340 -5866 3446 -5469
rect 3574 -5866 3680 -5469
rect 3808 -5866 3914 -5469
rect 4042 -5866 4148 -5469
rect 4276 -5866 4382 -5469
rect 4510 -5866 4616 -5469
rect 4744 -5866 4850 -5469
rect 4978 -5866 5084 -5469
rect 5212 -5866 5318 -5469
rect 5446 -5866 5552 -5469
rect 5680 -5866 5786 -5469
rect 5914 -5866 6020 -5469
rect 6148 -5866 6254 -5469
rect 6382 -5866 6488 -5469
rect 6616 -5866 6722 -5469
rect 6850 -5866 6956 -5469
rect 7084 -5866 7190 -5469
rect 7318 -5866 7424 -5469
rect 7552 -5866 7658 -5469
rect 7786 -5866 7892 -5469
rect 8020 -5866 8126 -5469
rect 8254 -5866 8360 -5469
rect 8488 -5866 8594 -5469
rect 8722 -5866 8828 -5469
rect 8956 -5866 9062 -5469
rect 9190 -5866 9296 -5469
rect 9424 -5866 9530 -5469
rect 9658 -5866 9764 -5469
rect 9892 -5866 9998 -5469
rect 10126 -5866 10232 -5469
rect 10360 -5866 10466 -5469
rect 10594 -5866 10700 -5469
rect 10828 -5866 10934 -5469
rect 11062 -5866 11168 -5469
rect 11296 -5866 11402 -5469
rect 11530 -5866 11636 -5469
rect 11764 -5866 11870 -5469
rect 11998 -5866 12104 -5469
rect 12232 -5866 12338 -5469
rect 12466 -5866 12572 -5469
rect 12700 -5866 12806 -5469
rect 12934 -5866 13040 -5469
rect 13168 -5866 13274 -5469
rect 13402 -5866 13508 -5469
rect 13636 -5866 13742 -5469
rect 13870 -5866 13976 -5469
rect 14104 -5866 14210 -5469
rect 14338 -5866 14444 -5469
rect 14572 -5866 14678 -5469
rect 14806 -5866 14912 -5469
rect 15040 -5866 15146 -5469
rect 15274 -5866 15380 -5469
rect 15508 -5866 15614 -5469
rect 15742 -5866 15848 -5469
rect 15976 -5866 16082 -5469
rect 16210 -5866 16316 -5469
rect 16444 -5866 16550 -5469
rect 16678 -5866 16784 -5469
rect 16912 -5866 17018 -5469
rect 17146 -5866 17252 -5469
rect 17380 -5866 17486 -5469
rect 17614 -5866 17720 -5469
rect 17848 -5866 17954 -5469
rect 18082 -5866 18188 -5469
rect 18316 -5866 18422 -5469
rect 18550 -5866 18656 -5469
rect 18784 -5866 18890 -5469
rect 19018 -5866 19124 -5469
rect 19252 -5866 19358 -5469
rect 19486 -5866 19592 -5469
rect 19720 -5866 19826 -5469
rect 19954 -5866 20060 -5469
rect 20188 -5866 20294 -5469
rect 20422 -5866 20528 -5469
rect 20656 -5866 20762 -5469
rect 20890 -5866 20996 -5469
rect 21124 -5866 21230 -5469
rect 21358 -5866 21464 -5469
rect 21592 -5866 21698 -5469
rect 21826 -5866 21932 -5469
rect 22060 -5866 22166 -5469
rect 22294 -5866 22400 -5469
rect 22528 -5866 22634 -5469
rect 22762 -5866 22868 -5469
rect 22996 -5866 23102 -5469
rect 23230 -5866 23336 -5469
rect 23464 -5866 23570 -5469
rect 23698 -5866 23804 -5469
rect 23932 -5866 24038 -5469
rect 24166 -5866 24272 -5469
rect 24400 -5866 24506 -5469
rect 24634 -5866 24740 -5469
rect 24868 -5866 24974 -5469
rect 25102 -5866 25208 -5469
rect 25336 -5866 25442 -5469
rect 25570 -5866 25676 -5469
rect 25804 -5866 25910 -5469
rect 26038 -5866 26144 -5469
rect 26272 -5866 26378 -5469
rect 26506 -5866 26612 -5469
rect 26740 -5866 26846 -5469
rect 26974 -5866 27080 -5469
rect 27208 -5866 27314 -5469
rect 27442 -5866 27548 -5469
rect 27676 -5866 27782 -5469
rect 27910 -5866 28016 -5469
rect 28144 -5866 28250 -5469
rect 28378 -5866 28484 -5469
rect 28612 -5866 28718 -5469
rect 28846 -5866 28952 -5469
rect 29080 -5866 29186 -5469
rect 29314 -5866 29420 -5469
rect 29548 -5866 29654 -5469
rect 29782 -5866 29888 -5469
<< metal1 >>
rect -29894 5866 -29776 5878
rect -29894 5469 -29888 5866
rect -29782 5469 -29776 5866
rect -29894 5457 -29776 5469
rect -29660 5866 -29542 5878
rect -29660 5469 -29654 5866
rect -29548 5469 -29542 5866
rect -29660 5457 -29542 5469
rect -29426 5866 -29308 5878
rect -29426 5469 -29420 5866
rect -29314 5469 -29308 5866
rect -29426 5457 -29308 5469
rect -29192 5866 -29074 5878
rect -29192 5469 -29186 5866
rect -29080 5469 -29074 5866
rect -29192 5457 -29074 5469
rect -28958 5866 -28840 5878
rect -28958 5469 -28952 5866
rect -28846 5469 -28840 5866
rect -28958 5457 -28840 5469
rect -28724 5866 -28606 5878
rect -28724 5469 -28718 5866
rect -28612 5469 -28606 5866
rect -28724 5457 -28606 5469
rect -28490 5866 -28372 5878
rect -28490 5469 -28484 5866
rect -28378 5469 -28372 5866
rect -28490 5457 -28372 5469
rect -28256 5866 -28138 5878
rect -28256 5469 -28250 5866
rect -28144 5469 -28138 5866
rect -28256 5457 -28138 5469
rect -28022 5866 -27904 5878
rect -28022 5469 -28016 5866
rect -27910 5469 -27904 5866
rect -28022 5457 -27904 5469
rect -27788 5866 -27670 5878
rect -27788 5469 -27782 5866
rect -27676 5469 -27670 5866
rect -27788 5457 -27670 5469
rect -27554 5866 -27436 5878
rect -27554 5469 -27548 5866
rect -27442 5469 -27436 5866
rect -27554 5457 -27436 5469
rect -27320 5866 -27202 5878
rect -27320 5469 -27314 5866
rect -27208 5469 -27202 5866
rect -27320 5457 -27202 5469
rect -27086 5866 -26968 5878
rect -27086 5469 -27080 5866
rect -26974 5469 -26968 5866
rect -27086 5457 -26968 5469
rect -26852 5866 -26734 5878
rect -26852 5469 -26846 5866
rect -26740 5469 -26734 5866
rect -26852 5457 -26734 5469
rect -26618 5866 -26500 5878
rect -26618 5469 -26612 5866
rect -26506 5469 -26500 5866
rect -26618 5457 -26500 5469
rect -26384 5866 -26266 5878
rect -26384 5469 -26378 5866
rect -26272 5469 -26266 5866
rect -26384 5457 -26266 5469
rect -26150 5866 -26032 5878
rect -26150 5469 -26144 5866
rect -26038 5469 -26032 5866
rect -26150 5457 -26032 5469
rect -25916 5866 -25798 5878
rect -25916 5469 -25910 5866
rect -25804 5469 -25798 5866
rect -25916 5457 -25798 5469
rect -25682 5866 -25564 5878
rect -25682 5469 -25676 5866
rect -25570 5469 -25564 5866
rect -25682 5457 -25564 5469
rect -25448 5866 -25330 5878
rect -25448 5469 -25442 5866
rect -25336 5469 -25330 5866
rect -25448 5457 -25330 5469
rect -25214 5866 -25096 5878
rect -25214 5469 -25208 5866
rect -25102 5469 -25096 5866
rect -25214 5457 -25096 5469
rect -24980 5866 -24862 5878
rect -24980 5469 -24974 5866
rect -24868 5469 -24862 5866
rect -24980 5457 -24862 5469
rect -24746 5866 -24628 5878
rect -24746 5469 -24740 5866
rect -24634 5469 -24628 5866
rect -24746 5457 -24628 5469
rect -24512 5866 -24394 5878
rect -24512 5469 -24506 5866
rect -24400 5469 -24394 5866
rect -24512 5457 -24394 5469
rect -24278 5866 -24160 5878
rect -24278 5469 -24272 5866
rect -24166 5469 -24160 5866
rect -24278 5457 -24160 5469
rect -24044 5866 -23926 5878
rect -24044 5469 -24038 5866
rect -23932 5469 -23926 5866
rect -24044 5457 -23926 5469
rect -23810 5866 -23692 5878
rect -23810 5469 -23804 5866
rect -23698 5469 -23692 5866
rect -23810 5457 -23692 5469
rect -23576 5866 -23458 5878
rect -23576 5469 -23570 5866
rect -23464 5469 -23458 5866
rect -23576 5457 -23458 5469
rect -23342 5866 -23224 5878
rect -23342 5469 -23336 5866
rect -23230 5469 -23224 5866
rect -23342 5457 -23224 5469
rect -23108 5866 -22990 5878
rect -23108 5469 -23102 5866
rect -22996 5469 -22990 5866
rect -23108 5457 -22990 5469
rect -22874 5866 -22756 5878
rect -22874 5469 -22868 5866
rect -22762 5469 -22756 5866
rect -22874 5457 -22756 5469
rect -22640 5866 -22522 5878
rect -22640 5469 -22634 5866
rect -22528 5469 -22522 5866
rect -22640 5457 -22522 5469
rect -22406 5866 -22288 5878
rect -22406 5469 -22400 5866
rect -22294 5469 -22288 5866
rect -22406 5457 -22288 5469
rect -22172 5866 -22054 5878
rect -22172 5469 -22166 5866
rect -22060 5469 -22054 5866
rect -22172 5457 -22054 5469
rect -21938 5866 -21820 5878
rect -21938 5469 -21932 5866
rect -21826 5469 -21820 5866
rect -21938 5457 -21820 5469
rect -21704 5866 -21586 5878
rect -21704 5469 -21698 5866
rect -21592 5469 -21586 5866
rect -21704 5457 -21586 5469
rect -21470 5866 -21352 5878
rect -21470 5469 -21464 5866
rect -21358 5469 -21352 5866
rect -21470 5457 -21352 5469
rect -21236 5866 -21118 5878
rect -21236 5469 -21230 5866
rect -21124 5469 -21118 5866
rect -21236 5457 -21118 5469
rect -21002 5866 -20884 5878
rect -21002 5469 -20996 5866
rect -20890 5469 -20884 5866
rect -21002 5457 -20884 5469
rect -20768 5866 -20650 5878
rect -20768 5469 -20762 5866
rect -20656 5469 -20650 5866
rect -20768 5457 -20650 5469
rect -20534 5866 -20416 5878
rect -20534 5469 -20528 5866
rect -20422 5469 -20416 5866
rect -20534 5457 -20416 5469
rect -20300 5866 -20182 5878
rect -20300 5469 -20294 5866
rect -20188 5469 -20182 5866
rect -20300 5457 -20182 5469
rect -20066 5866 -19948 5878
rect -20066 5469 -20060 5866
rect -19954 5469 -19948 5866
rect -20066 5457 -19948 5469
rect -19832 5866 -19714 5878
rect -19832 5469 -19826 5866
rect -19720 5469 -19714 5866
rect -19832 5457 -19714 5469
rect -19598 5866 -19480 5878
rect -19598 5469 -19592 5866
rect -19486 5469 -19480 5866
rect -19598 5457 -19480 5469
rect -19364 5866 -19246 5878
rect -19364 5469 -19358 5866
rect -19252 5469 -19246 5866
rect -19364 5457 -19246 5469
rect -19130 5866 -19012 5878
rect -19130 5469 -19124 5866
rect -19018 5469 -19012 5866
rect -19130 5457 -19012 5469
rect -18896 5866 -18778 5878
rect -18896 5469 -18890 5866
rect -18784 5469 -18778 5866
rect -18896 5457 -18778 5469
rect -18662 5866 -18544 5878
rect -18662 5469 -18656 5866
rect -18550 5469 -18544 5866
rect -18662 5457 -18544 5469
rect -18428 5866 -18310 5878
rect -18428 5469 -18422 5866
rect -18316 5469 -18310 5866
rect -18428 5457 -18310 5469
rect -18194 5866 -18076 5878
rect -18194 5469 -18188 5866
rect -18082 5469 -18076 5866
rect -18194 5457 -18076 5469
rect -17960 5866 -17842 5878
rect -17960 5469 -17954 5866
rect -17848 5469 -17842 5866
rect -17960 5457 -17842 5469
rect -17726 5866 -17608 5878
rect -17726 5469 -17720 5866
rect -17614 5469 -17608 5866
rect -17726 5457 -17608 5469
rect -17492 5866 -17374 5878
rect -17492 5469 -17486 5866
rect -17380 5469 -17374 5866
rect -17492 5457 -17374 5469
rect -17258 5866 -17140 5878
rect -17258 5469 -17252 5866
rect -17146 5469 -17140 5866
rect -17258 5457 -17140 5469
rect -17024 5866 -16906 5878
rect -17024 5469 -17018 5866
rect -16912 5469 -16906 5866
rect -17024 5457 -16906 5469
rect -16790 5866 -16672 5878
rect -16790 5469 -16784 5866
rect -16678 5469 -16672 5866
rect -16790 5457 -16672 5469
rect -16556 5866 -16438 5878
rect -16556 5469 -16550 5866
rect -16444 5469 -16438 5866
rect -16556 5457 -16438 5469
rect -16322 5866 -16204 5878
rect -16322 5469 -16316 5866
rect -16210 5469 -16204 5866
rect -16322 5457 -16204 5469
rect -16088 5866 -15970 5878
rect -16088 5469 -16082 5866
rect -15976 5469 -15970 5866
rect -16088 5457 -15970 5469
rect -15854 5866 -15736 5878
rect -15854 5469 -15848 5866
rect -15742 5469 -15736 5866
rect -15854 5457 -15736 5469
rect -15620 5866 -15502 5878
rect -15620 5469 -15614 5866
rect -15508 5469 -15502 5866
rect -15620 5457 -15502 5469
rect -15386 5866 -15268 5878
rect -15386 5469 -15380 5866
rect -15274 5469 -15268 5866
rect -15386 5457 -15268 5469
rect -15152 5866 -15034 5878
rect -15152 5469 -15146 5866
rect -15040 5469 -15034 5866
rect -15152 5457 -15034 5469
rect -14918 5866 -14800 5878
rect -14918 5469 -14912 5866
rect -14806 5469 -14800 5866
rect -14918 5457 -14800 5469
rect -14684 5866 -14566 5878
rect -14684 5469 -14678 5866
rect -14572 5469 -14566 5866
rect -14684 5457 -14566 5469
rect -14450 5866 -14332 5878
rect -14450 5469 -14444 5866
rect -14338 5469 -14332 5866
rect -14450 5457 -14332 5469
rect -14216 5866 -14098 5878
rect -14216 5469 -14210 5866
rect -14104 5469 -14098 5866
rect -14216 5457 -14098 5469
rect -13982 5866 -13864 5878
rect -13982 5469 -13976 5866
rect -13870 5469 -13864 5866
rect -13982 5457 -13864 5469
rect -13748 5866 -13630 5878
rect -13748 5469 -13742 5866
rect -13636 5469 -13630 5866
rect -13748 5457 -13630 5469
rect -13514 5866 -13396 5878
rect -13514 5469 -13508 5866
rect -13402 5469 -13396 5866
rect -13514 5457 -13396 5469
rect -13280 5866 -13162 5878
rect -13280 5469 -13274 5866
rect -13168 5469 -13162 5866
rect -13280 5457 -13162 5469
rect -13046 5866 -12928 5878
rect -13046 5469 -13040 5866
rect -12934 5469 -12928 5866
rect -13046 5457 -12928 5469
rect -12812 5866 -12694 5878
rect -12812 5469 -12806 5866
rect -12700 5469 -12694 5866
rect -12812 5457 -12694 5469
rect -12578 5866 -12460 5878
rect -12578 5469 -12572 5866
rect -12466 5469 -12460 5866
rect -12578 5457 -12460 5469
rect -12344 5866 -12226 5878
rect -12344 5469 -12338 5866
rect -12232 5469 -12226 5866
rect -12344 5457 -12226 5469
rect -12110 5866 -11992 5878
rect -12110 5469 -12104 5866
rect -11998 5469 -11992 5866
rect -12110 5457 -11992 5469
rect -11876 5866 -11758 5878
rect -11876 5469 -11870 5866
rect -11764 5469 -11758 5866
rect -11876 5457 -11758 5469
rect -11642 5866 -11524 5878
rect -11642 5469 -11636 5866
rect -11530 5469 -11524 5866
rect -11642 5457 -11524 5469
rect -11408 5866 -11290 5878
rect -11408 5469 -11402 5866
rect -11296 5469 -11290 5866
rect -11408 5457 -11290 5469
rect -11174 5866 -11056 5878
rect -11174 5469 -11168 5866
rect -11062 5469 -11056 5866
rect -11174 5457 -11056 5469
rect -10940 5866 -10822 5878
rect -10940 5469 -10934 5866
rect -10828 5469 -10822 5866
rect -10940 5457 -10822 5469
rect -10706 5866 -10588 5878
rect -10706 5469 -10700 5866
rect -10594 5469 -10588 5866
rect -10706 5457 -10588 5469
rect -10472 5866 -10354 5878
rect -10472 5469 -10466 5866
rect -10360 5469 -10354 5866
rect -10472 5457 -10354 5469
rect -10238 5866 -10120 5878
rect -10238 5469 -10232 5866
rect -10126 5469 -10120 5866
rect -10238 5457 -10120 5469
rect -10004 5866 -9886 5878
rect -10004 5469 -9998 5866
rect -9892 5469 -9886 5866
rect -10004 5457 -9886 5469
rect -9770 5866 -9652 5878
rect -9770 5469 -9764 5866
rect -9658 5469 -9652 5866
rect -9770 5457 -9652 5469
rect -9536 5866 -9418 5878
rect -9536 5469 -9530 5866
rect -9424 5469 -9418 5866
rect -9536 5457 -9418 5469
rect -9302 5866 -9184 5878
rect -9302 5469 -9296 5866
rect -9190 5469 -9184 5866
rect -9302 5457 -9184 5469
rect -9068 5866 -8950 5878
rect -9068 5469 -9062 5866
rect -8956 5469 -8950 5866
rect -9068 5457 -8950 5469
rect -8834 5866 -8716 5878
rect -8834 5469 -8828 5866
rect -8722 5469 -8716 5866
rect -8834 5457 -8716 5469
rect -8600 5866 -8482 5878
rect -8600 5469 -8594 5866
rect -8488 5469 -8482 5866
rect -8600 5457 -8482 5469
rect -8366 5866 -8248 5878
rect -8366 5469 -8360 5866
rect -8254 5469 -8248 5866
rect -8366 5457 -8248 5469
rect -8132 5866 -8014 5878
rect -8132 5469 -8126 5866
rect -8020 5469 -8014 5866
rect -8132 5457 -8014 5469
rect -7898 5866 -7780 5878
rect -7898 5469 -7892 5866
rect -7786 5469 -7780 5866
rect -7898 5457 -7780 5469
rect -7664 5866 -7546 5878
rect -7664 5469 -7658 5866
rect -7552 5469 -7546 5866
rect -7664 5457 -7546 5469
rect -7430 5866 -7312 5878
rect -7430 5469 -7424 5866
rect -7318 5469 -7312 5866
rect -7430 5457 -7312 5469
rect -7196 5866 -7078 5878
rect -7196 5469 -7190 5866
rect -7084 5469 -7078 5866
rect -7196 5457 -7078 5469
rect -6962 5866 -6844 5878
rect -6962 5469 -6956 5866
rect -6850 5469 -6844 5866
rect -6962 5457 -6844 5469
rect -6728 5866 -6610 5878
rect -6728 5469 -6722 5866
rect -6616 5469 -6610 5866
rect -6728 5457 -6610 5469
rect -6494 5866 -6376 5878
rect -6494 5469 -6488 5866
rect -6382 5469 -6376 5866
rect -6494 5457 -6376 5469
rect -6260 5866 -6142 5878
rect -6260 5469 -6254 5866
rect -6148 5469 -6142 5866
rect -6260 5457 -6142 5469
rect -6026 5866 -5908 5878
rect -6026 5469 -6020 5866
rect -5914 5469 -5908 5866
rect -6026 5457 -5908 5469
rect -5792 5866 -5674 5878
rect -5792 5469 -5786 5866
rect -5680 5469 -5674 5866
rect -5792 5457 -5674 5469
rect -5558 5866 -5440 5878
rect -5558 5469 -5552 5866
rect -5446 5469 -5440 5866
rect -5558 5457 -5440 5469
rect -5324 5866 -5206 5878
rect -5324 5469 -5318 5866
rect -5212 5469 -5206 5866
rect -5324 5457 -5206 5469
rect -5090 5866 -4972 5878
rect -5090 5469 -5084 5866
rect -4978 5469 -4972 5866
rect -5090 5457 -4972 5469
rect -4856 5866 -4738 5878
rect -4856 5469 -4850 5866
rect -4744 5469 -4738 5866
rect -4856 5457 -4738 5469
rect -4622 5866 -4504 5878
rect -4622 5469 -4616 5866
rect -4510 5469 -4504 5866
rect -4622 5457 -4504 5469
rect -4388 5866 -4270 5878
rect -4388 5469 -4382 5866
rect -4276 5469 -4270 5866
rect -4388 5457 -4270 5469
rect -4154 5866 -4036 5878
rect -4154 5469 -4148 5866
rect -4042 5469 -4036 5866
rect -4154 5457 -4036 5469
rect -3920 5866 -3802 5878
rect -3920 5469 -3914 5866
rect -3808 5469 -3802 5866
rect -3920 5457 -3802 5469
rect -3686 5866 -3568 5878
rect -3686 5469 -3680 5866
rect -3574 5469 -3568 5866
rect -3686 5457 -3568 5469
rect -3452 5866 -3334 5878
rect -3452 5469 -3446 5866
rect -3340 5469 -3334 5866
rect -3452 5457 -3334 5469
rect -3218 5866 -3100 5878
rect -3218 5469 -3212 5866
rect -3106 5469 -3100 5866
rect -3218 5457 -3100 5469
rect -2984 5866 -2866 5878
rect -2984 5469 -2978 5866
rect -2872 5469 -2866 5866
rect -2984 5457 -2866 5469
rect -2750 5866 -2632 5878
rect -2750 5469 -2744 5866
rect -2638 5469 -2632 5866
rect -2750 5457 -2632 5469
rect -2516 5866 -2398 5878
rect -2516 5469 -2510 5866
rect -2404 5469 -2398 5866
rect -2516 5457 -2398 5469
rect -2282 5866 -2164 5878
rect -2282 5469 -2276 5866
rect -2170 5469 -2164 5866
rect -2282 5457 -2164 5469
rect -2048 5866 -1930 5878
rect -2048 5469 -2042 5866
rect -1936 5469 -1930 5866
rect -2048 5457 -1930 5469
rect -1814 5866 -1696 5878
rect -1814 5469 -1808 5866
rect -1702 5469 -1696 5866
rect -1814 5457 -1696 5469
rect -1580 5866 -1462 5878
rect -1580 5469 -1574 5866
rect -1468 5469 -1462 5866
rect -1580 5457 -1462 5469
rect -1346 5866 -1228 5878
rect -1346 5469 -1340 5866
rect -1234 5469 -1228 5866
rect -1346 5457 -1228 5469
rect -1112 5866 -994 5878
rect -1112 5469 -1106 5866
rect -1000 5469 -994 5866
rect -1112 5457 -994 5469
rect -878 5866 -760 5878
rect -878 5469 -872 5866
rect -766 5469 -760 5866
rect -878 5457 -760 5469
rect -644 5866 -526 5878
rect -644 5469 -638 5866
rect -532 5469 -526 5866
rect -644 5457 -526 5469
rect -410 5866 -292 5878
rect -410 5469 -404 5866
rect -298 5469 -292 5866
rect -410 5457 -292 5469
rect -176 5866 -58 5878
rect -176 5469 -170 5866
rect -64 5469 -58 5866
rect -176 5457 -58 5469
rect 58 5866 176 5878
rect 58 5469 64 5866
rect 170 5469 176 5866
rect 58 5457 176 5469
rect 292 5866 410 5878
rect 292 5469 298 5866
rect 404 5469 410 5866
rect 292 5457 410 5469
rect 526 5866 644 5878
rect 526 5469 532 5866
rect 638 5469 644 5866
rect 526 5457 644 5469
rect 760 5866 878 5878
rect 760 5469 766 5866
rect 872 5469 878 5866
rect 760 5457 878 5469
rect 994 5866 1112 5878
rect 994 5469 1000 5866
rect 1106 5469 1112 5866
rect 994 5457 1112 5469
rect 1228 5866 1346 5878
rect 1228 5469 1234 5866
rect 1340 5469 1346 5866
rect 1228 5457 1346 5469
rect 1462 5866 1580 5878
rect 1462 5469 1468 5866
rect 1574 5469 1580 5866
rect 1462 5457 1580 5469
rect 1696 5866 1814 5878
rect 1696 5469 1702 5866
rect 1808 5469 1814 5866
rect 1696 5457 1814 5469
rect 1930 5866 2048 5878
rect 1930 5469 1936 5866
rect 2042 5469 2048 5866
rect 1930 5457 2048 5469
rect 2164 5866 2282 5878
rect 2164 5469 2170 5866
rect 2276 5469 2282 5866
rect 2164 5457 2282 5469
rect 2398 5866 2516 5878
rect 2398 5469 2404 5866
rect 2510 5469 2516 5866
rect 2398 5457 2516 5469
rect 2632 5866 2750 5878
rect 2632 5469 2638 5866
rect 2744 5469 2750 5866
rect 2632 5457 2750 5469
rect 2866 5866 2984 5878
rect 2866 5469 2872 5866
rect 2978 5469 2984 5866
rect 2866 5457 2984 5469
rect 3100 5866 3218 5878
rect 3100 5469 3106 5866
rect 3212 5469 3218 5866
rect 3100 5457 3218 5469
rect 3334 5866 3452 5878
rect 3334 5469 3340 5866
rect 3446 5469 3452 5866
rect 3334 5457 3452 5469
rect 3568 5866 3686 5878
rect 3568 5469 3574 5866
rect 3680 5469 3686 5866
rect 3568 5457 3686 5469
rect 3802 5866 3920 5878
rect 3802 5469 3808 5866
rect 3914 5469 3920 5866
rect 3802 5457 3920 5469
rect 4036 5866 4154 5878
rect 4036 5469 4042 5866
rect 4148 5469 4154 5866
rect 4036 5457 4154 5469
rect 4270 5866 4388 5878
rect 4270 5469 4276 5866
rect 4382 5469 4388 5866
rect 4270 5457 4388 5469
rect 4504 5866 4622 5878
rect 4504 5469 4510 5866
rect 4616 5469 4622 5866
rect 4504 5457 4622 5469
rect 4738 5866 4856 5878
rect 4738 5469 4744 5866
rect 4850 5469 4856 5866
rect 4738 5457 4856 5469
rect 4972 5866 5090 5878
rect 4972 5469 4978 5866
rect 5084 5469 5090 5866
rect 4972 5457 5090 5469
rect 5206 5866 5324 5878
rect 5206 5469 5212 5866
rect 5318 5469 5324 5866
rect 5206 5457 5324 5469
rect 5440 5866 5558 5878
rect 5440 5469 5446 5866
rect 5552 5469 5558 5866
rect 5440 5457 5558 5469
rect 5674 5866 5792 5878
rect 5674 5469 5680 5866
rect 5786 5469 5792 5866
rect 5674 5457 5792 5469
rect 5908 5866 6026 5878
rect 5908 5469 5914 5866
rect 6020 5469 6026 5866
rect 5908 5457 6026 5469
rect 6142 5866 6260 5878
rect 6142 5469 6148 5866
rect 6254 5469 6260 5866
rect 6142 5457 6260 5469
rect 6376 5866 6494 5878
rect 6376 5469 6382 5866
rect 6488 5469 6494 5866
rect 6376 5457 6494 5469
rect 6610 5866 6728 5878
rect 6610 5469 6616 5866
rect 6722 5469 6728 5866
rect 6610 5457 6728 5469
rect 6844 5866 6962 5878
rect 6844 5469 6850 5866
rect 6956 5469 6962 5866
rect 6844 5457 6962 5469
rect 7078 5866 7196 5878
rect 7078 5469 7084 5866
rect 7190 5469 7196 5866
rect 7078 5457 7196 5469
rect 7312 5866 7430 5878
rect 7312 5469 7318 5866
rect 7424 5469 7430 5866
rect 7312 5457 7430 5469
rect 7546 5866 7664 5878
rect 7546 5469 7552 5866
rect 7658 5469 7664 5866
rect 7546 5457 7664 5469
rect 7780 5866 7898 5878
rect 7780 5469 7786 5866
rect 7892 5469 7898 5866
rect 7780 5457 7898 5469
rect 8014 5866 8132 5878
rect 8014 5469 8020 5866
rect 8126 5469 8132 5866
rect 8014 5457 8132 5469
rect 8248 5866 8366 5878
rect 8248 5469 8254 5866
rect 8360 5469 8366 5866
rect 8248 5457 8366 5469
rect 8482 5866 8600 5878
rect 8482 5469 8488 5866
rect 8594 5469 8600 5866
rect 8482 5457 8600 5469
rect 8716 5866 8834 5878
rect 8716 5469 8722 5866
rect 8828 5469 8834 5866
rect 8716 5457 8834 5469
rect 8950 5866 9068 5878
rect 8950 5469 8956 5866
rect 9062 5469 9068 5866
rect 8950 5457 9068 5469
rect 9184 5866 9302 5878
rect 9184 5469 9190 5866
rect 9296 5469 9302 5866
rect 9184 5457 9302 5469
rect 9418 5866 9536 5878
rect 9418 5469 9424 5866
rect 9530 5469 9536 5866
rect 9418 5457 9536 5469
rect 9652 5866 9770 5878
rect 9652 5469 9658 5866
rect 9764 5469 9770 5866
rect 9652 5457 9770 5469
rect 9886 5866 10004 5878
rect 9886 5469 9892 5866
rect 9998 5469 10004 5866
rect 9886 5457 10004 5469
rect 10120 5866 10238 5878
rect 10120 5469 10126 5866
rect 10232 5469 10238 5866
rect 10120 5457 10238 5469
rect 10354 5866 10472 5878
rect 10354 5469 10360 5866
rect 10466 5469 10472 5866
rect 10354 5457 10472 5469
rect 10588 5866 10706 5878
rect 10588 5469 10594 5866
rect 10700 5469 10706 5866
rect 10588 5457 10706 5469
rect 10822 5866 10940 5878
rect 10822 5469 10828 5866
rect 10934 5469 10940 5866
rect 10822 5457 10940 5469
rect 11056 5866 11174 5878
rect 11056 5469 11062 5866
rect 11168 5469 11174 5866
rect 11056 5457 11174 5469
rect 11290 5866 11408 5878
rect 11290 5469 11296 5866
rect 11402 5469 11408 5866
rect 11290 5457 11408 5469
rect 11524 5866 11642 5878
rect 11524 5469 11530 5866
rect 11636 5469 11642 5866
rect 11524 5457 11642 5469
rect 11758 5866 11876 5878
rect 11758 5469 11764 5866
rect 11870 5469 11876 5866
rect 11758 5457 11876 5469
rect 11992 5866 12110 5878
rect 11992 5469 11998 5866
rect 12104 5469 12110 5866
rect 11992 5457 12110 5469
rect 12226 5866 12344 5878
rect 12226 5469 12232 5866
rect 12338 5469 12344 5866
rect 12226 5457 12344 5469
rect 12460 5866 12578 5878
rect 12460 5469 12466 5866
rect 12572 5469 12578 5866
rect 12460 5457 12578 5469
rect 12694 5866 12812 5878
rect 12694 5469 12700 5866
rect 12806 5469 12812 5866
rect 12694 5457 12812 5469
rect 12928 5866 13046 5878
rect 12928 5469 12934 5866
rect 13040 5469 13046 5866
rect 12928 5457 13046 5469
rect 13162 5866 13280 5878
rect 13162 5469 13168 5866
rect 13274 5469 13280 5866
rect 13162 5457 13280 5469
rect 13396 5866 13514 5878
rect 13396 5469 13402 5866
rect 13508 5469 13514 5866
rect 13396 5457 13514 5469
rect 13630 5866 13748 5878
rect 13630 5469 13636 5866
rect 13742 5469 13748 5866
rect 13630 5457 13748 5469
rect 13864 5866 13982 5878
rect 13864 5469 13870 5866
rect 13976 5469 13982 5866
rect 13864 5457 13982 5469
rect 14098 5866 14216 5878
rect 14098 5469 14104 5866
rect 14210 5469 14216 5866
rect 14098 5457 14216 5469
rect 14332 5866 14450 5878
rect 14332 5469 14338 5866
rect 14444 5469 14450 5866
rect 14332 5457 14450 5469
rect 14566 5866 14684 5878
rect 14566 5469 14572 5866
rect 14678 5469 14684 5866
rect 14566 5457 14684 5469
rect 14800 5866 14918 5878
rect 14800 5469 14806 5866
rect 14912 5469 14918 5866
rect 14800 5457 14918 5469
rect 15034 5866 15152 5878
rect 15034 5469 15040 5866
rect 15146 5469 15152 5866
rect 15034 5457 15152 5469
rect 15268 5866 15386 5878
rect 15268 5469 15274 5866
rect 15380 5469 15386 5866
rect 15268 5457 15386 5469
rect 15502 5866 15620 5878
rect 15502 5469 15508 5866
rect 15614 5469 15620 5866
rect 15502 5457 15620 5469
rect 15736 5866 15854 5878
rect 15736 5469 15742 5866
rect 15848 5469 15854 5866
rect 15736 5457 15854 5469
rect 15970 5866 16088 5878
rect 15970 5469 15976 5866
rect 16082 5469 16088 5866
rect 15970 5457 16088 5469
rect 16204 5866 16322 5878
rect 16204 5469 16210 5866
rect 16316 5469 16322 5866
rect 16204 5457 16322 5469
rect 16438 5866 16556 5878
rect 16438 5469 16444 5866
rect 16550 5469 16556 5866
rect 16438 5457 16556 5469
rect 16672 5866 16790 5878
rect 16672 5469 16678 5866
rect 16784 5469 16790 5866
rect 16672 5457 16790 5469
rect 16906 5866 17024 5878
rect 16906 5469 16912 5866
rect 17018 5469 17024 5866
rect 16906 5457 17024 5469
rect 17140 5866 17258 5878
rect 17140 5469 17146 5866
rect 17252 5469 17258 5866
rect 17140 5457 17258 5469
rect 17374 5866 17492 5878
rect 17374 5469 17380 5866
rect 17486 5469 17492 5866
rect 17374 5457 17492 5469
rect 17608 5866 17726 5878
rect 17608 5469 17614 5866
rect 17720 5469 17726 5866
rect 17608 5457 17726 5469
rect 17842 5866 17960 5878
rect 17842 5469 17848 5866
rect 17954 5469 17960 5866
rect 17842 5457 17960 5469
rect 18076 5866 18194 5878
rect 18076 5469 18082 5866
rect 18188 5469 18194 5866
rect 18076 5457 18194 5469
rect 18310 5866 18428 5878
rect 18310 5469 18316 5866
rect 18422 5469 18428 5866
rect 18310 5457 18428 5469
rect 18544 5866 18662 5878
rect 18544 5469 18550 5866
rect 18656 5469 18662 5866
rect 18544 5457 18662 5469
rect 18778 5866 18896 5878
rect 18778 5469 18784 5866
rect 18890 5469 18896 5866
rect 18778 5457 18896 5469
rect 19012 5866 19130 5878
rect 19012 5469 19018 5866
rect 19124 5469 19130 5866
rect 19012 5457 19130 5469
rect 19246 5866 19364 5878
rect 19246 5469 19252 5866
rect 19358 5469 19364 5866
rect 19246 5457 19364 5469
rect 19480 5866 19598 5878
rect 19480 5469 19486 5866
rect 19592 5469 19598 5866
rect 19480 5457 19598 5469
rect 19714 5866 19832 5878
rect 19714 5469 19720 5866
rect 19826 5469 19832 5866
rect 19714 5457 19832 5469
rect 19948 5866 20066 5878
rect 19948 5469 19954 5866
rect 20060 5469 20066 5866
rect 19948 5457 20066 5469
rect 20182 5866 20300 5878
rect 20182 5469 20188 5866
rect 20294 5469 20300 5866
rect 20182 5457 20300 5469
rect 20416 5866 20534 5878
rect 20416 5469 20422 5866
rect 20528 5469 20534 5866
rect 20416 5457 20534 5469
rect 20650 5866 20768 5878
rect 20650 5469 20656 5866
rect 20762 5469 20768 5866
rect 20650 5457 20768 5469
rect 20884 5866 21002 5878
rect 20884 5469 20890 5866
rect 20996 5469 21002 5866
rect 20884 5457 21002 5469
rect 21118 5866 21236 5878
rect 21118 5469 21124 5866
rect 21230 5469 21236 5866
rect 21118 5457 21236 5469
rect 21352 5866 21470 5878
rect 21352 5469 21358 5866
rect 21464 5469 21470 5866
rect 21352 5457 21470 5469
rect 21586 5866 21704 5878
rect 21586 5469 21592 5866
rect 21698 5469 21704 5866
rect 21586 5457 21704 5469
rect 21820 5866 21938 5878
rect 21820 5469 21826 5866
rect 21932 5469 21938 5866
rect 21820 5457 21938 5469
rect 22054 5866 22172 5878
rect 22054 5469 22060 5866
rect 22166 5469 22172 5866
rect 22054 5457 22172 5469
rect 22288 5866 22406 5878
rect 22288 5469 22294 5866
rect 22400 5469 22406 5866
rect 22288 5457 22406 5469
rect 22522 5866 22640 5878
rect 22522 5469 22528 5866
rect 22634 5469 22640 5866
rect 22522 5457 22640 5469
rect 22756 5866 22874 5878
rect 22756 5469 22762 5866
rect 22868 5469 22874 5866
rect 22756 5457 22874 5469
rect 22990 5866 23108 5878
rect 22990 5469 22996 5866
rect 23102 5469 23108 5866
rect 22990 5457 23108 5469
rect 23224 5866 23342 5878
rect 23224 5469 23230 5866
rect 23336 5469 23342 5866
rect 23224 5457 23342 5469
rect 23458 5866 23576 5878
rect 23458 5469 23464 5866
rect 23570 5469 23576 5866
rect 23458 5457 23576 5469
rect 23692 5866 23810 5878
rect 23692 5469 23698 5866
rect 23804 5469 23810 5866
rect 23692 5457 23810 5469
rect 23926 5866 24044 5878
rect 23926 5469 23932 5866
rect 24038 5469 24044 5866
rect 23926 5457 24044 5469
rect 24160 5866 24278 5878
rect 24160 5469 24166 5866
rect 24272 5469 24278 5866
rect 24160 5457 24278 5469
rect 24394 5866 24512 5878
rect 24394 5469 24400 5866
rect 24506 5469 24512 5866
rect 24394 5457 24512 5469
rect 24628 5866 24746 5878
rect 24628 5469 24634 5866
rect 24740 5469 24746 5866
rect 24628 5457 24746 5469
rect 24862 5866 24980 5878
rect 24862 5469 24868 5866
rect 24974 5469 24980 5866
rect 24862 5457 24980 5469
rect 25096 5866 25214 5878
rect 25096 5469 25102 5866
rect 25208 5469 25214 5866
rect 25096 5457 25214 5469
rect 25330 5866 25448 5878
rect 25330 5469 25336 5866
rect 25442 5469 25448 5866
rect 25330 5457 25448 5469
rect 25564 5866 25682 5878
rect 25564 5469 25570 5866
rect 25676 5469 25682 5866
rect 25564 5457 25682 5469
rect 25798 5866 25916 5878
rect 25798 5469 25804 5866
rect 25910 5469 25916 5866
rect 25798 5457 25916 5469
rect 26032 5866 26150 5878
rect 26032 5469 26038 5866
rect 26144 5469 26150 5866
rect 26032 5457 26150 5469
rect 26266 5866 26384 5878
rect 26266 5469 26272 5866
rect 26378 5469 26384 5866
rect 26266 5457 26384 5469
rect 26500 5866 26618 5878
rect 26500 5469 26506 5866
rect 26612 5469 26618 5866
rect 26500 5457 26618 5469
rect 26734 5866 26852 5878
rect 26734 5469 26740 5866
rect 26846 5469 26852 5866
rect 26734 5457 26852 5469
rect 26968 5866 27086 5878
rect 26968 5469 26974 5866
rect 27080 5469 27086 5866
rect 26968 5457 27086 5469
rect 27202 5866 27320 5878
rect 27202 5469 27208 5866
rect 27314 5469 27320 5866
rect 27202 5457 27320 5469
rect 27436 5866 27554 5878
rect 27436 5469 27442 5866
rect 27548 5469 27554 5866
rect 27436 5457 27554 5469
rect 27670 5866 27788 5878
rect 27670 5469 27676 5866
rect 27782 5469 27788 5866
rect 27670 5457 27788 5469
rect 27904 5866 28022 5878
rect 27904 5469 27910 5866
rect 28016 5469 28022 5866
rect 27904 5457 28022 5469
rect 28138 5866 28256 5878
rect 28138 5469 28144 5866
rect 28250 5469 28256 5866
rect 28138 5457 28256 5469
rect 28372 5866 28490 5878
rect 28372 5469 28378 5866
rect 28484 5469 28490 5866
rect 28372 5457 28490 5469
rect 28606 5866 28724 5878
rect 28606 5469 28612 5866
rect 28718 5469 28724 5866
rect 28606 5457 28724 5469
rect 28840 5866 28958 5878
rect 28840 5469 28846 5866
rect 28952 5469 28958 5866
rect 28840 5457 28958 5469
rect 29074 5866 29192 5878
rect 29074 5469 29080 5866
rect 29186 5469 29192 5866
rect 29074 5457 29192 5469
rect 29308 5866 29426 5878
rect 29308 5469 29314 5866
rect 29420 5469 29426 5866
rect 29308 5457 29426 5469
rect 29542 5866 29660 5878
rect 29542 5469 29548 5866
rect 29654 5469 29660 5866
rect 29542 5457 29660 5469
rect 29776 5866 29894 5878
rect 29776 5469 29782 5866
rect 29888 5469 29894 5866
rect 29776 5457 29894 5469
rect -29894 467 -29776 479
rect -29894 70 -29888 467
rect -29782 70 -29776 467
rect -29894 58 -29776 70
rect -29660 467 -29542 479
rect -29660 70 -29654 467
rect -29548 70 -29542 467
rect -29660 58 -29542 70
rect -29426 467 -29308 479
rect -29426 70 -29420 467
rect -29314 70 -29308 467
rect -29426 58 -29308 70
rect -29192 467 -29074 479
rect -29192 70 -29186 467
rect -29080 70 -29074 467
rect -29192 58 -29074 70
rect -28958 467 -28840 479
rect -28958 70 -28952 467
rect -28846 70 -28840 467
rect -28958 58 -28840 70
rect -28724 467 -28606 479
rect -28724 70 -28718 467
rect -28612 70 -28606 467
rect -28724 58 -28606 70
rect -28490 467 -28372 479
rect -28490 70 -28484 467
rect -28378 70 -28372 467
rect -28490 58 -28372 70
rect -28256 467 -28138 479
rect -28256 70 -28250 467
rect -28144 70 -28138 467
rect -28256 58 -28138 70
rect -28022 467 -27904 479
rect -28022 70 -28016 467
rect -27910 70 -27904 467
rect -28022 58 -27904 70
rect -27788 467 -27670 479
rect -27788 70 -27782 467
rect -27676 70 -27670 467
rect -27788 58 -27670 70
rect -27554 467 -27436 479
rect -27554 70 -27548 467
rect -27442 70 -27436 467
rect -27554 58 -27436 70
rect -27320 467 -27202 479
rect -27320 70 -27314 467
rect -27208 70 -27202 467
rect -27320 58 -27202 70
rect -27086 467 -26968 479
rect -27086 70 -27080 467
rect -26974 70 -26968 467
rect -27086 58 -26968 70
rect -26852 467 -26734 479
rect -26852 70 -26846 467
rect -26740 70 -26734 467
rect -26852 58 -26734 70
rect -26618 467 -26500 479
rect -26618 70 -26612 467
rect -26506 70 -26500 467
rect -26618 58 -26500 70
rect -26384 467 -26266 479
rect -26384 70 -26378 467
rect -26272 70 -26266 467
rect -26384 58 -26266 70
rect -26150 467 -26032 479
rect -26150 70 -26144 467
rect -26038 70 -26032 467
rect -26150 58 -26032 70
rect -25916 467 -25798 479
rect -25916 70 -25910 467
rect -25804 70 -25798 467
rect -25916 58 -25798 70
rect -25682 467 -25564 479
rect -25682 70 -25676 467
rect -25570 70 -25564 467
rect -25682 58 -25564 70
rect -25448 467 -25330 479
rect -25448 70 -25442 467
rect -25336 70 -25330 467
rect -25448 58 -25330 70
rect -25214 467 -25096 479
rect -25214 70 -25208 467
rect -25102 70 -25096 467
rect -25214 58 -25096 70
rect -24980 467 -24862 479
rect -24980 70 -24974 467
rect -24868 70 -24862 467
rect -24980 58 -24862 70
rect -24746 467 -24628 479
rect -24746 70 -24740 467
rect -24634 70 -24628 467
rect -24746 58 -24628 70
rect -24512 467 -24394 479
rect -24512 70 -24506 467
rect -24400 70 -24394 467
rect -24512 58 -24394 70
rect -24278 467 -24160 479
rect -24278 70 -24272 467
rect -24166 70 -24160 467
rect -24278 58 -24160 70
rect -24044 467 -23926 479
rect -24044 70 -24038 467
rect -23932 70 -23926 467
rect -24044 58 -23926 70
rect -23810 467 -23692 479
rect -23810 70 -23804 467
rect -23698 70 -23692 467
rect -23810 58 -23692 70
rect -23576 467 -23458 479
rect -23576 70 -23570 467
rect -23464 70 -23458 467
rect -23576 58 -23458 70
rect -23342 467 -23224 479
rect -23342 70 -23336 467
rect -23230 70 -23224 467
rect -23342 58 -23224 70
rect -23108 467 -22990 479
rect -23108 70 -23102 467
rect -22996 70 -22990 467
rect -23108 58 -22990 70
rect -22874 467 -22756 479
rect -22874 70 -22868 467
rect -22762 70 -22756 467
rect -22874 58 -22756 70
rect -22640 467 -22522 479
rect -22640 70 -22634 467
rect -22528 70 -22522 467
rect -22640 58 -22522 70
rect -22406 467 -22288 479
rect -22406 70 -22400 467
rect -22294 70 -22288 467
rect -22406 58 -22288 70
rect -22172 467 -22054 479
rect -22172 70 -22166 467
rect -22060 70 -22054 467
rect -22172 58 -22054 70
rect -21938 467 -21820 479
rect -21938 70 -21932 467
rect -21826 70 -21820 467
rect -21938 58 -21820 70
rect -21704 467 -21586 479
rect -21704 70 -21698 467
rect -21592 70 -21586 467
rect -21704 58 -21586 70
rect -21470 467 -21352 479
rect -21470 70 -21464 467
rect -21358 70 -21352 467
rect -21470 58 -21352 70
rect -21236 467 -21118 479
rect -21236 70 -21230 467
rect -21124 70 -21118 467
rect -21236 58 -21118 70
rect -21002 467 -20884 479
rect -21002 70 -20996 467
rect -20890 70 -20884 467
rect -21002 58 -20884 70
rect -20768 467 -20650 479
rect -20768 70 -20762 467
rect -20656 70 -20650 467
rect -20768 58 -20650 70
rect -20534 467 -20416 479
rect -20534 70 -20528 467
rect -20422 70 -20416 467
rect -20534 58 -20416 70
rect -20300 467 -20182 479
rect -20300 70 -20294 467
rect -20188 70 -20182 467
rect -20300 58 -20182 70
rect -20066 467 -19948 479
rect -20066 70 -20060 467
rect -19954 70 -19948 467
rect -20066 58 -19948 70
rect -19832 467 -19714 479
rect -19832 70 -19826 467
rect -19720 70 -19714 467
rect -19832 58 -19714 70
rect -19598 467 -19480 479
rect -19598 70 -19592 467
rect -19486 70 -19480 467
rect -19598 58 -19480 70
rect -19364 467 -19246 479
rect -19364 70 -19358 467
rect -19252 70 -19246 467
rect -19364 58 -19246 70
rect -19130 467 -19012 479
rect -19130 70 -19124 467
rect -19018 70 -19012 467
rect -19130 58 -19012 70
rect -18896 467 -18778 479
rect -18896 70 -18890 467
rect -18784 70 -18778 467
rect -18896 58 -18778 70
rect -18662 467 -18544 479
rect -18662 70 -18656 467
rect -18550 70 -18544 467
rect -18662 58 -18544 70
rect -18428 467 -18310 479
rect -18428 70 -18422 467
rect -18316 70 -18310 467
rect -18428 58 -18310 70
rect -18194 467 -18076 479
rect -18194 70 -18188 467
rect -18082 70 -18076 467
rect -18194 58 -18076 70
rect -17960 467 -17842 479
rect -17960 70 -17954 467
rect -17848 70 -17842 467
rect -17960 58 -17842 70
rect -17726 467 -17608 479
rect -17726 70 -17720 467
rect -17614 70 -17608 467
rect -17726 58 -17608 70
rect -17492 467 -17374 479
rect -17492 70 -17486 467
rect -17380 70 -17374 467
rect -17492 58 -17374 70
rect -17258 467 -17140 479
rect -17258 70 -17252 467
rect -17146 70 -17140 467
rect -17258 58 -17140 70
rect -17024 467 -16906 479
rect -17024 70 -17018 467
rect -16912 70 -16906 467
rect -17024 58 -16906 70
rect -16790 467 -16672 479
rect -16790 70 -16784 467
rect -16678 70 -16672 467
rect -16790 58 -16672 70
rect -16556 467 -16438 479
rect -16556 70 -16550 467
rect -16444 70 -16438 467
rect -16556 58 -16438 70
rect -16322 467 -16204 479
rect -16322 70 -16316 467
rect -16210 70 -16204 467
rect -16322 58 -16204 70
rect -16088 467 -15970 479
rect -16088 70 -16082 467
rect -15976 70 -15970 467
rect -16088 58 -15970 70
rect -15854 467 -15736 479
rect -15854 70 -15848 467
rect -15742 70 -15736 467
rect -15854 58 -15736 70
rect -15620 467 -15502 479
rect -15620 70 -15614 467
rect -15508 70 -15502 467
rect -15620 58 -15502 70
rect -15386 467 -15268 479
rect -15386 70 -15380 467
rect -15274 70 -15268 467
rect -15386 58 -15268 70
rect -15152 467 -15034 479
rect -15152 70 -15146 467
rect -15040 70 -15034 467
rect -15152 58 -15034 70
rect -14918 467 -14800 479
rect -14918 70 -14912 467
rect -14806 70 -14800 467
rect -14918 58 -14800 70
rect -14684 467 -14566 479
rect -14684 70 -14678 467
rect -14572 70 -14566 467
rect -14684 58 -14566 70
rect -14450 467 -14332 479
rect -14450 70 -14444 467
rect -14338 70 -14332 467
rect -14450 58 -14332 70
rect -14216 467 -14098 479
rect -14216 70 -14210 467
rect -14104 70 -14098 467
rect -14216 58 -14098 70
rect -13982 467 -13864 479
rect -13982 70 -13976 467
rect -13870 70 -13864 467
rect -13982 58 -13864 70
rect -13748 467 -13630 479
rect -13748 70 -13742 467
rect -13636 70 -13630 467
rect -13748 58 -13630 70
rect -13514 467 -13396 479
rect -13514 70 -13508 467
rect -13402 70 -13396 467
rect -13514 58 -13396 70
rect -13280 467 -13162 479
rect -13280 70 -13274 467
rect -13168 70 -13162 467
rect -13280 58 -13162 70
rect -13046 467 -12928 479
rect -13046 70 -13040 467
rect -12934 70 -12928 467
rect -13046 58 -12928 70
rect -12812 467 -12694 479
rect -12812 70 -12806 467
rect -12700 70 -12694 467
rect -12812 58 -12694 70
rect -12578 467 -12460 479
rect -12578 70 -12572 467
rect -12466 70 -12460 467
rect -12578 58 -12460 70
rect -12344 467 -12226 479
rect -12344 70 -12338 467
rect -12232 70 -12226 467
rect -12344 58 -12226 70
rect -12110 467 -11992 479
rect -12110 70 -12104 467
rect -11998 70 -11992 467
rect -12110 58 -11992 70
rect -11876 467 -11758 479
rect -11876 70 -11870 467
rect -11764 70 -11758 467
rect -11876 58 -11758 70
rect -11642 467 -11524 479
rect -11642 70 -11636 467
rect -11530 70 -11524 467
rect -11642 58 -11524 70
rect -11408 467 -11290 479
rect -11408 70 -11402 467
rect -11296 70 -11290 467
rect -11408 58 -11290 70
rect -11174 467 -11056 479
rect -11174 70 -11168 467
rect -11062 70 -11056 467
rect -11174 58 -11056 70
rect -10940 467 -10822 479
rect -10940 70 -10934 467
rect -10828 70 -10822 467
rect -10940 58 -10822 70
rect -10706 467 -10588 479
rect -10706 70 -10700 467
rect -10594 70 -10588 467
rect -10706 58 -10588 70
rect -10472 467 -10354 479
rect -10472 70 -10466 467
rect -10360 70 -10354 467
rect -10472 58 -10354 70
rect -10238 467 -10120 479
rect -10238 70 -10232 467
rect -10126 70 -10120 467
rect -10238 58 -10120 70
rect -10004 467 -9886 479
rect -10004 70 -9998 467
rect -9892 70 -9886 467
rect -10004 58 -9886 70
rect -9770 467 -9652 479
rect -9770 70 -9764 467
rect -9658 70 -9652 467
rect -9770 58 -9652 70
rect -9536 467 -9418 479
rect -9536 70 -9530 467
rect -9424 70 -9418 467
rect -9536 58 -9418 70
rect -9302 467 -9184 479
rect -9302 70 -9296 467
rect -9190 70 -9184 467
rect -9302 58 -9184 70
rect -9068 467 -8950 479
rect -9068 70 -9062 467
rect -8956 70 -8950 467
rect -9068 58 -8950 70
rect -8834 467 -8716 479
rect -8834 70 -8828 467
rect -8722 70 -8716 467
rect -8834 58 -8716 70
rect -8600 467 -8482 479
rect -8600 70 -8594 467
rect -8488 70 -8482 467
rect -8600 58 -8482 70
rect -8366 467 -8248 479
rect -8366 70 -8360 467
rect -8254 70 -8248 467
rect -8366 58 -8248 70
rect -8132 467 -8014 479
rect -8132 70 -8126 467
rect -8020 70 -8014 467
rect -8132 58 -8014 70
rect -7898 467 -7780 479
rect -7898 70 -7892 467
rect -7786 70 -7780 467
rect -7898 58 -7780 70
rect -7664 467 -7546 479
rect -7664 70 -7658 467
rect -7552 70 -7546 467
rect -7664 58 -7546 70
rect -7430 467 -7312 479
rect -7430 70 -7424 467
rect -7318 70 -7312 467
rect -7430 58 -7312 70
rect -7196 467 -7078 479
rect -7196 70 -7190 467
rect -7084 70 -7078 467
rect -7196 58 -7078 70
rect -6962 467 -6844 479
rect -6962 70 -6956 467
rect -6850 70 -6844 467
rect -6962 58 -6844 70
rect -6728 467 -6610 479
rect -6728 70 -6722 467
rect -6616 70 -6610 467
rect -6728 58 -6610 70
rect -6494 467 -6376 479
rect -6494 70 -6488 467
rect -6382 70 -6376 467
rect -6494 58 -6376 70
rect -6260 467 -6142 479
rect -6260 70 -6254 467
rect -6148 70 -6142 467
rect -6260 58 -6142 70
rect -6026 467 -5908 479
rect -6026 70 -6020 467
rect -5914 70 -5908 467
rect -6026 58 -5908 70
rect -5792 467 -5674 479
rect -5792 70 -5786 467
rect -5680 70 -5674 467
rect -5792 58 -5674 70
rect -5558 467 -5440 479
rect -5558 70 -5552 467
rect -5446 70 -5440 467
rect -5558 58 -5440 70
rect -5324 467 -5206 479
rect -5324 70 -5318 467
rect -5212 70 -5206 467
rect -5324 58 -5206 70
rect -5090 467 -4972 479
rect -5090 70 -5084 467
rect -4978 70 -4972 467
rect -5090 58 -4972 70
rect -4856 467 -4738 479
rect -4856 70 -4850 467
rect -4744 70 -4738 467
rect -4856 58 -4738 70
rect -4622 467 -4504 479
rect -4622 70 -4616 467
rect -4510 70 -4504 467
rect -4622 58 -4504 70
rect -4388 467 -4270 479
rect -4388 70 -4382 467
rect -4276 70 -4270 467
rect -4388 58 -4270 70
rect -4154 467 -4036 479
rect -4154 70 -4148 467
rect -4042 70 -4036 467
rect -4154 58 -4036 70
rect -3920 467 -3802 479
rect -3920 70 -3914 467
rect -3808 70 -3802 467
rect -3920 58 -3802 70
rect -3686 467 -3568 479
rect -3686 70 -3680 467
rect -3574 70 -3568 467
rect -3686 58 -3568 70
rect -3452 467 -3334 479
rect -3452 70 -3446 467
rect -3340 70 -3334 467
rect -3452 58 -3334 70
rect -3218 467 -3100 479
rect -3218 70 -3212 467
rect -3106 70 -3100 467
rect -3218 58 -3100 70
rect -2984 467 -2866 479
rect -2984 70 -2978 467
rect -2872 70 -2866 467
rect -2984 58 -2866 70
rect -2750 467 -2632 479
rect -2750 70 -2744 467
rect -2638 70 -2632 467
rect -2750 58 -2632 70
rect -2516 467 -2398 479
rect -2516 70 -2510 467
rect -2404 70 -2398 467
rect -2516 58 -2398 70
rect -2282 467 -2164 479
rect -2282 70 -2276 467
rect -2170 70 -2164 467
rect -2282 58 -2164 70
rect -2048 467 -1930 479
rect -2048 70 -2042 467
rect -1936 70 -1930 467
rect -2048 58 -1930 70
rect -1814 467 -1696 479
rect -1814 70 -1808 467
rect -1702 70 -1696 467
rect -1814 58 -1696 70
rect -1580 467 -1462 479
rect -1580 70 -1574 467
rect -1468 70 -1462 467
rect -1580 58 -1462 70
rect -1346 467 -1228 479
rect -1346 70 -1340 467
rect -1234 70 -1228 467
rect -1346 58 -1228 70
rect -1112 467 -994 479
rect -1112 70 -1106 467
rect -1000 70 -994 467
rect -1112 58 -994 70
rect -878 467 -760 479
rect -878 70 -872 467
rect -766 70 -760 467
rect -878 58 -760 70
rect -644 467 -526 479
rect -644 70 -638 467
rect -532 70 -526 467
rect -644 58 -526 70
rect -410 467 -292 479
rect -410 70 -404 467
rect -298 70 -292 467
rect -410 58 -292 70
rect -176 467 -58 479
rect -176 70 -170 467
rect -64 70 -58 467
rect -176 58 -58 70
rect 58 467 176 479
rect 58 70 64 467
rect 170 70 176 467
rect 58 58 176 70
rect 292 467 410 479
rect 292 70 298 467
rect 404 70 410 467
rect 292 58 410 70
rect 526 467 644 479
rect 526 70 532 467
rect 638 70 644 467
rect 526 58 644 70
rect 760 467 878 479
rect 760 70 766 467
rect 872 70 878 467
rect 760 58 878 70
rect 994 467 1112 479
rect 994 70 1000 467
rect 1106 70 1112 467
rect 994 58 1112 70
rect 1228 467 1346 479
rect 1228 70 1234 467
rect 1340 70 1346 467
rect 1228 58 1346 70
rect 1462 467 1580 479
rect 1462 70 1468 467
rect 1574 70 1580 467
rect 1462 58 1580 70
rect 1696 467 1814 479
rect 1696 70 1702 467
rect 1808 70 1814 467
rect 1696 58 1814 70
rect 1930 467 2048 479
rect 1930 70 1936 467
rect 2042 70 2048 467
rect 1930 58 2048 70
rect 2164 467 2282 479
rect 2164 70 2170 467
rect 2276 70 2282 467
rect 2164 58 2282 70
rect 2398 467 2516 479
rect 2398 70 2404 467
rect 2510 70 2516 467
rect 2398 58 2516 70
rect 2632 467 2750 479
rect 2632 70 2638 467
rect 2744 70 2750 467
rect 2632 58 2750 70
rect 2866 467 2984 479
rect 2866 70 2872 467
rect 2978 70 2984 467
rect 2866 58 2984 70
rect 3100 467 3218 479
rect 3100 70 3106 467
rect 3212 70 3218 467
rect 3100 58 3218 70
rect 3334 467 3452 479
rect 3334 70 3340 467
rect 3446 70 3452 467
rect 3334 58 3452 70
rect 3568 467 3686 479
rect 3568 70 3574 467
rect 3680 70 3686 467
rect 3568 58 3686 70
rect 3802 467 3920 479
rect 3802 70 3808 467
rect 3914 70 3920 467
rect 3802 58 3920 70
rect 4036 467 4154 479
rect 4036 70 4042 467
rect 4148 70 4154 467
rect 4036 58 4154 70
rect 4270 467 4388 479
rect 4270 70 4276 467
rect 4382 70 4388 467
rect 4270 58 4388 70
rect 4504 467 4622 479
rect 4504 70 4510 467
rect 4616 70 4622 467
rect 4504 58 4622 70
rect 4738 467 4856 479
rect 4738 70 4744 467
rect 4850 70 4856 467
rect 4738 58 4856 70
rect 4972 467 5090 479
rect 4972 70 4978 467
rect 5084 70 5090 467
rect 4972 58 5090 70
rect 5206 467 5324 479
rect 5206 70 5212 467
rect 5318 70 5324 467
rect 5206 58 5324 70
rect 5440 467 5558 479
rect 5440 70 5446 467
rect 5552 70 5558 467
rect 5440 58 5558 70
rect 5674 467 5792 479
rect 5674 70 5680 467
rect 5786 70 5792 467
rect 5674 58 5792 70
rect 5908 467 6026 479
rect 5908 70 5914 467
rect 6020 70 6026 467
rect 5908 58 6026 70
rect 6142 467 6260 479
rect 6142 70 6148 467
rect 6254 70 6260 467
rect 6142 58 6260 70
rect 6376 467 6494 479
rect 6376 70 6382 467
rect 6488 70 6494 467
rect 6376 58 6494 70
rect 6610 467 6728 479
rect 6610 70 6616 467
rect 6722 70 6728 467
rect 6610 58 6728 70
rect 6844 467 6962 479
rect 6844 70 6850 467
rect 6956 70 6962 467
rect 6844 58 6962 70
rect 7078 467 7196 479
rect 7078 70 7084 467
rect 7190 70 7196 467
rect 7078 58 7196 70
rect 7312 467 7430 479
rect 7312 70 7318 467
rect 7424 70 7430 467
rect 7312 58 7430 70
rect 7546 467 7664 479
rect 7546 70 7552 467
rect 7658 70 7664 467
rect 7546 58 7664 70
rect 7780 467 7898 479
rect 7780 70 7786 467
rect 7892 70 7898 467
rect 7780 58 7898 70
rect 8014 467 8132 479
rect 8014 70 8020 467
rect 8126 70 8132 467
rect 8014 58 8132 70
rect 8248 467 8366 479
rect 8248 70 8254 467
rect 8360 70 8366 467
rect 8248 58 8366 70
rect 8482 467 8600 479
rect 8482 70 8488 467
rect 8594 70 8600 467
rect 8482 58 8600 70
rect 8716 467 8834 479
rect 8716 70 8722 467
rect 8828 70 8834 467
rect 8716 58 8834 70
rect 8950 467 9068 479
rect 8950 70 8956 467
rect 9062 70 9068 467
rect 8950 58 9068 70
rect 9184 467 9302 479
rect 9184 70 9190 467
rect 9296 70 9302 467
rect 9184 58 9302 70
rect 9418 467 9536 479
rect 9418 70 9424 467
rect 9530 70 9536 467
rect 9418 58 9536 70
rect 9652 467 9770 479
rect 9652 70 9658 467
rect 9764 70 9770 467
rect 9652 58 9770 70
rect 9886 467 10004 479
rect 9886 70 9892 467
rect 9998 70 10004 467
rect 9886 58 10004 70
rect 10120 467 10238 479
rect 10120 70 10126 467
rect 10232 70 10238 467
rect 10120 58 10238 70
rect 10354 467 10472 479
rect 10354 70 10360 467
rect 10466 70 10472 467
rect 10354 58 10472 70
rect 10588 467 10706 479
rect 10588 70 10594 467
rect 10700 70 10706 467
rect 10588 58 10706 70
rect 10822 467 10940 479
rect 10822 70 10828 467
rect 10934 70 10940 467
rect 10822 58 10940 70
rect 11056 467 11174 479
rect 11056 70 11062 467
rect 11168 70 11174 467
rect 11056 58 11174 70
rect 11290 467 11408 479
rect 11290 70 11296 467
rect 11402 70 11408 467
rect 11290 58 11408 70
rect 11524 467 11642 479
rect 11524 70 11530 467
rect 11636 70 11642 467
rect 11524 58 11642 70
rect 11758 467 11876 479
rect 11758 70 11764 467
rect 11870 70 11876 467
rect 11758 58 11876 70
rect 11992 467 12110 479
rect 11992 70 11998 467
rect 12104 70 12110 467
rect 11992 58 12110 70
rect 12226 467 12344 479
rect 12226 70 12232 467
rect 12338 70 12344 467
rect 12226 58 12344 70
rect 12460 467 12578 479
rect 12460 70 12466 467
rect 12572 70 12578 467
rect 12460 58 12578 70
rect 12694 467 12812 479
rect 12694 70 12700 467
rect 12806 70 12812 467
rect 12694 58 12812 70
rect 12928 467 13046 479
rect 12928 70 12934 467
rect 13040 70 13046 467
rect 12928 58 13046 70
rect 13162 467 13280 479
rect 13162 70 13168 467
rect 13274 70 13280 467
rect 13162 58 13280 70
rect 13396 467 13514 479
rect 13396 70 13402 467
rect 13508 70 13514 467
rect 13396 58 13514 70
rect 13630 467 13748 479
rect 13630 70 13636 467
rect 13742 70 13748 467
rect 13630 58 13748 70
rect 13864 467 13982 479
rect 13864 70 13870 467
rect 13976 70 13982 467
rect 13864 58 13982 70
rect 14098 467 14216 479
rect 14098 70 14104 467
rect 14210 70 14216 467
rect 14098 58 14216 70
rect 14332 467 14450 479
rect 14332 70 14338 467
rect 14444 70 14450 467
rect 14332 58 14450 70
rect 14566 467 14684 479
rect 14566 70 14572 467
rect 14678 70 14684 467
rect 14566 58 14684 70
rect 14800 467 14918 479
rect 14800 70 14806 467
rect 14912 70 14918 467
rect 14800 58 14918 70
rect 15034 467 15152 479
rect 15034 70 15040 467
rect 15146 70 15152 467
rect 15034 58 15152 70
rect 15268 467 15386 479
rect 15268 70 15274 467
rect 15380 70 15386 467
rect 15268 58 15386 70
rect 15502 467 15620 479
rect 15502 70 15508 467
rect 15614 70 15620 467
rect 15502 58 15620 70
rect 15736 467 15854 479
rect 15736 70 15742 467
rect 15848 70 15854 467
rect 15736 58 15854 70
rect 15970 467 16088 479
rect 15970 70 15976 467
rect 16082 70 16088 467
rect 15970 58 16088 70
rect 16204 467 16322 479
rect 16204 70 16210 467
rect 16316 70 16322 467
rect 16204 58 16322 70
rect 16438 467 16556 479
rect 16438 70 16444 467
rect 16550 70 16556 467
rect 16438 58 16556 70
rect 16672 467 16790 479
rect 16672 70 16678 467
rect 16784 70 16790 467
rect 16672 58 16790 70
rect 16906 467 17024 479
rect 16906 70 16912 467
rect 17018 70 17024 467
rect 16906 58 17024 70
rect 17140 467 17258 479
rect 17140 70 17146 467
rect 17252 70 17258 467
rect 17140 58 17258 70
rect 17374 467 17492 479
rect 17374 70 17380 467
rect 17486 70 17492 467
rect 17374 58 17492 70
rect 17608 467 17726 479
rect 17608 70 17614 467
rect 17720 70 17726 467
rect 17608 58 17726 70
rect 17842 467 17960 479
rect 17842 70 17848 467
rect 17954 70 17960 467
rect 17842 58 17960 70
rect 18076 467 18194 479
rect 18076 70 18082 467
rect 18188 70 18194 467
rect 18076 58 18194 70
rect 18310 467 18428 479
rect 18310 70 18316 467
rect 18422 70 18428 467
rect 18310 58 18428 70
rect 18544 467 18662 479
rect 18544 70 18550 467
rect 18656 70 18662 467
rect 18544 58 18662 70
rect 18778 467 18896 479
rect 18778 70 18784 467
rect 18890 70 18896 467
rect 18778 58 18896 70
rect 19012 467 19130 479
rect 19012 70 19018 467
rect 19124 70 19130 467
rect 19012 58 19130 70
rect 19246 467 19364 479
rect 19246 70 19252 467
rect 19358 70 19364 467
rect 19246 58 19364 70
rect 19480 467 19598 479
rect 19480 70 19486 467
rect 19592 70 19598 467
rect 19480 58 19598 70
rect 19714 467 19832 479
rect 19714 70 19720 467
rect 19826 70 19832 467
rect 19714 58 19832 70
rect 19948 467 20066 479
rect 19948 70 19954 467
rect 20060 70 20066 467
rect 19948 58 20066 70
rect 20182 467 20300 479
rect 20182 70 20188 467
rect 20294 70 20300 467
rect 20182 58 20300 70
rect 20416 467 20534 479
rect 20416 70 20422 467
rect 20528 70 20534 467
rect 20416 58 20534 70
rect 20650 467 20768 479
rect 20650 70 20656 467
rect 20762 70 20768 467
rect 20650 58 20768 70
rect 20884 467 21002 479
rect 20884 70 20890 467
rect 20996 70 21002 467
rect 20884 58 21002 70
rect 21118 467 21236 479
rect 21118 70 21124 467
rect 21230 70 21236 467
rect 21118 58 21236 70
rect 21352 467 21470 479
rect 21352 70 21358 467
rect 21464 70 21470 467
rect 21352 58 21470 70
rect 21586 467 21704 479
rect 21586 70 21592 467
rect 21698 70 21704 467
rect 21586 58 21704 70
rect 21820 467 21938 479
rect 21820 70 21826 467
rect 21932 70 21938 467
rect 21820 58 21938 70
rect 22054 467 22172 479
rect 22054 70 22060 467
rect 22166 70 22172 467
rect 22054 58 22172 70
rect 22288 467 22406 479
rect 22288 70 22294 467
rect 22400 70 22406 467
rect 22288 58 22406 70
rect 22522 467 22640 479
rect 22522 70 22528 467
rect 22634 70 22640 467
rect 22522 58 22640 70
rect 22756 467 22874 479
rect 22756 70 22762 467
rect 22868 70 22874 467
rect 22756 58 22874 70
rect 22990 467 23108 479
rect 22990 70 22996 467
rect 23102 70 23108 467
rect 22990 58 23108 70
rect 23224 467 23342 479
rect 23224 70 23230 467
rect 23336 70 23342 467
rect 23224 58 23342 70
rect 23458 467 23576 479
rect 23458 70 23464 467
rect 23570 70 23576 467
rect 23458 58 23576 70
rect 23692 467 23810 479
rect 23692 70 23698 467
rect 23804 70 23810 467
rect 23692 58 23810 70
rect 23926 467 24044 479
rect 23926 70 23932 467
rect 24038 70 24044 467
rect 23926 58 24044 70
rect 24160 467 24278 479
rect 24160 70 24166 467
rect 24272 70 24278 467
rect 24160 58 24278 70
rect 24394 467 24512 479
rect 24394 70 24400 467
rect 24506 70 24512 467
rect 24394 58 24512 70
rect 24628 467 24746 479
rect 24628 70 24634 467
rect 24740 70 24746 467
rect 24628 58 24746 70
rect 24862 467 24980 479
rect 24862 70 24868 467
rect 24974 70 24980 467
rect 24862 58 24980 70
rect 25096 467 25214 479
rect 25096 70 25102 467
rect 25208 70 25214 467
rect 25096 58 25214 70
rect 25330 467 25448 479
rect 25330 70 25336 467
rect 25442 70 25448 467
rect 25330 58 25448 70
rect 25564 467 25682 479
rect 25564 70 25570 467
rect 25676 70 25682 467
rect 25564 58 25682 70
rect 25798 467 25916 479
rect 25798 70 25804 467
rect 25910 70 25916 467
rect 25798 58 25916 70
rect 26032 467 26150 479
rect 26032 70 26038 467
rect 26144 70 26150 467
rect 26032 58 26150 70
rect 26266 467 26384 479
rect 26266 70 26272 467
rect 26378 70 26384 467
rect 26266 58 26384 70
rect 26500 467 26618 479
rect 26500 70 26506 467
rect 26612 70 26618 467
rect 26500 58 26618 70
rect 26734 467 26852 479
rect 26734 70 26740 467
rect 26846 70 26852 467
rect 26734 58 26852 70
rect 26968 467 27086 479
rect 26968 70 26974 467
rect 27080 70 27086 467
rect 26968 58 27086 70
rect 27202 467 27320 479
rect 27202 70 27208 467
rect 27314 70 27320 467
rect 27202 58 27320 70
rect 27436 467 27554 479
rect 27436 70 27442 467
rect 27548 70 27554 467
rect 27436 58 27554 70
rect 27670 467 27788 479
rect 27670 70 27676 467
rect 27782 70 27788 467
rect 27670 58 27788 70
rect 27904 467 28022 479
rect 27904 70 27910 467
rect 28016 70 28022 467
rect 27904 58 28022 70
rect 28138 467 28256 479
rect 28138 70 28144 467
rect 28250 70 28256 467
rect 28138 58 28256 70
rect 28372 467 28490 479
rect 28372 70 28378 467
rect 28484 70 28490 467
rect 28372 58 28490 70
rect 28606 467 28724 479
rect 28606 70 28612 467
rect 28718 70 28724 467
rect 28606 58 28724 70
rect 28840 467 28958 479
rect 28840 70 28846 467
rect 28952 70 28958 467
rect 28840 58 28958 70
rect 29074 467 29192 479
rect 29074 70 29080 467
rect 29186 70 29192 467
rect 29074 58 29192 70
rect 29308 467 29426 479
rect 29308 70 29314 467
rect 29420 70 29426 467
rect 29308 58 29426 70
rect 29542 467 29660 479
rect 29542 70 29548 467
rect 29654 70 29660 467
rect 29542 58 29660 70
rect 29776 467 29894 479
rect 29776 70 29782 467
rect 29888 70 29894 467
rect 29776 58 29894 70
rect -29894 -70 -29776 -58
rect -29894 -467 -29888 -70
rect -29782 -467 -29776 -70
rect -29894 -479 -29776 -467
rect -29660 -70 -29542 -58
rect -29660 -467 -29654 -70
rect -29548 -467 -29542 -70
rect -29660 -479 -29542 -467
rect -29426 -70 -29308 -58
rect -29426 -467 -29420 -70
rect -29314 -467 -29308 -70
rect -29426 -479 -29308 -467
rect -29192 -70 -29074 -58
rect -29192 -467 -29186 -70
rect -29080 -467 -29074 -70
rect -29192 -479 -29074 -467
rect -28958 -70 -28840 -58
rect -28958 -467 -28952 -70
rect -28846 -467 -28840 -70
rect -28958 -479 -28840 -467
rect -28724 -70 -28606 -58
rect -28724 -467 -28718 -70
rect -28612 -467 -28606 -70
rect -28724 -479 -28606 -467
rect -28490 -70 -28372 -58
rect -28490 -467 -28484 -70
rect -28378 -467 -28372 -70
rect -28490 -479 -28372 -467
rect -28256 -70 -28138 -58
rect -28256 -467 -28250 -70
rect -28144 -467 -28138 -70
rect -28256 -479 -28138 -467
rect -28022 -70 -27904 -58
rect -28022 -467 -28016 -70
rect -27910 -467 -27904 -70
rect -28022 -479 -27904 -467
rect -27788 -70 -27670 -58
rect -27788 -467 -27782 -70
rect -27676 -467 -27670 -70
rect -27788 -479 -27670 -467
rect -27554 -70 -27436 -58
rect -27554 -467 -27548 -70
rect -27442 -467 -27436 -70
rect -27554 -479 -27436 -467
rect -27320 -70 -27202 -58
rect -27320 -467 -27314 -70
rect -27208 -467 -27202 -70
rect -27320 -479 -27202 -467
rect -27086 -70 -26968 -58
rect -27086 -467 -27080 -70
rect -26974 -467 -26968 -70
rect -27086 -479 -26968 -467
rect -26852 -70 -26734 -58
rect -26852 -467 -26846 -70
rect -26740 -467 -26734 -70
rect -26852 -479 -26734 -467
rect -26618 -70 -26500 -58
rect -26618 -467 -26612 -70
rect -26506 -467 -26500 -70
rect -26618 -479 -26500 -467
rect -26384 -70 -26266 -58
rect -26384 -467 -26378 -70
rect -26272 -467 -26266 -70
rect -26384 -479 -26266 -467
rect -26150 -70 -26032 -58
rect -26150 -467 -26144 -70
rect -26038 -467 -26032 -70
rect -26150 -479 -26032 -467
rect -25916 -70 -25798 -58
rect -25916 -467 -25910 -70
rect -25804 -467 -25798 -70
rect -25916 -479 -25798 -467
rect -25682 -70 -25564 -58
rect -25682 -467 -25676 -70
rect -25570 -467 -25564 -70
rect -25682 -479 -25564 -467
rect -25448 -70 -25330 -58
rect -25448 -467 -25442 -70
rect -25336 -467 -25330 -70
rect -25448 -479 -25330 -467
rect -25214 -70 -25096 -58
rect -25214 -467 -25208 -70
rect -25102 -467 -25096 -70
rect -25214 -479 -25096 -467
rect -24980 -70 -24862 -58
rect -24980 -467 -24974 -70
rect -24868 -467 -24862 -70
rect -24980 -479 -24862 -467
rect -24746 -70 -24628 -58
rect -24746 -467 -24740 -70
rect -24634 -467 -24628 -70
rect -24746 -479 -24628 -467
rect -24512 -70 -24394 -58
rect -24512 -467 -24506 -70
rect -24400 -467 -24394 -70
rect -24512 -479 -24394 -467
rect -24278 -70 -24160 -58
rect -24278 -467 -24272 -70
rect -24166 -467 -24160 -70
rect -24278 -479 -24160 -467
rect -24044 -70 -23926 -58
rect -24044 -467 -24038 -70
rect -23932 -467 -23926 -70
rect -24044 -479 -23926 -467
rect -23810 -70 -23692 -58
rect -23810 -467 -23804 -70
rect -23698 -467 -23692 -70
rect -23810 -479 -23692 -467
rect -23576 -70 -23458 -58
rect -23576 -467 -23570 -70
rect -23464 -467 -23458 -70
rect -23576 -479 -23458 -467
rect -23342 -70 -23224 -58
rect -23342 -467 -23336 -70
rect -23230 -467 -23224 -70
rect -23342 -479 -23224 -467
rect -23108 -70 -22990 -58
rect -23108 -467 -23102 -70
rect -22996 -467 -22990 -70
rect -23108 -479 -22990 -467
rect -22874 -70 -22756 -58
rect -22874 -467 -22868 -70
rect -22762 -467 -22756 -70
rect -22874 -479 -22756 -467
rect -22640 -70 -22522 -58
rect -22640 -467 -22634 -70
rect -22528 -467 -22522 -70
rect -22640 -479 -22522 -467
rect -22406 -70 -22288 -58
rect -22406 -467 -22400 -70
rect -22294 -467 -22288 -70
rect -22406 -479 -22288 -467
rect -22172 -70 -22054 -58
rect -22172 -467 -22166 -70
rect -22060 -467 -22054 -70
rect -22172 -479 -22054 -467
rect -21938 -70 -21820 -58
rect -21938 -467 -21932 -70
rect -21826 -467 -21820 -70
rect -21938 -479 -21820 -467
rect -21704 -70 -21586 -58
rect -21704 -467 -21698 -70
rect -21592 -467 -21586 -70
rect -21704 -479 -21586 -467
rect -21470 -70 -21352 -58
rect -21470 -467 -21464 -70
rect -21358 -467 -21352 -70
rect -21470 -479 -21352 -467
rect -21236 -70 -21118 -58
rect -21236 -467 -21230 -70
rect -21124 -467 -21118 -70
rect -21236 -479 -21118 -467
rect -21002 -70 -20884 -58
rect -21002 -467 -20996 -70
rect -20890 -467 -20884 -70
rect -21002 -479 -20884 -467
rect -20768 -70 -20650 -58
rect -20768 -467 -20762 -70
rect -20656 -467 -20650 -70
rect -20768 -479 -20650 -467
rect -20534 -70 -20416 -58
rect -20534 -467 -20528 -70
rect -20422 -467 -20416 -70
rect -20534 -479 -20416 -467
rect -20300 -70 -20182 -58
rect -20300 -467 -20294 -70
rect -20188 -467 -20182 -70
rect -20300 -479 -20182 -467
rect -20066 -70 -19948 -58
rect -20066 -467 -20060 -70
rect -19954 -467 -19948 -70
rect -20066 -479 -19948 -467
rect -19832 -70 -19714 -58
rect -19832 -467 -19826 -70
rect -19720 -467 -19714 -70
rect -19832 -479 -19714 -467
rect -19598 -70 -19480 -58
rect -19598 -467 -19592 -70
rect -19486 -467 -19480 -70
rect -19598 -479 -19480 -467
rect -19364 -70 -19246 -58
rect -19364 -467 -19358 -70
rect -19252 -467 -19246 -70
rect -19364 -479 -19246 -467
rect -19130 -70 -19012 -58
rect -19130 -467 -19124 -70
rect -19018 -467 -19012 -70
rect -19130 -479 -19012 -467
rect -18896 -70 -18778 -58
rect -18896 -467 -18890 -70
rect -18784 -467 -18778 -70
rect -18896 -479 -18778 -467
rect -18662 -70 -18544 -58
rect -18662 -467 -18656 -70
rect -18550 -467 -18544 -70
rect -18662 -479 -18544 -467
rect -18428 -70 -18310 -58
rect -18428 -467 -18422 -70
rect -18316 -467 -18310 -70
rect -18428 -479 -18310 -467
rect -18194 -70 -18076 -58
rect -18194 -467 -18188 -70
rect -18082 -467 -18076 -70
rect -18194 -479 -18076 -467
rect -17960 -70 -17842 -58
rect -17960 -467 -17954 -70
rect -17848 -467 -17842 -70
rect -17960 -479 -17842 -467
rect -17726 -70 -17608 -58
rect -17726 -467 -17720 -70
rect -17614 -467 -17608 -70
rect -17726 -479 -17608 -467
rect -17492 -70 -17374 -58
rect -17492 -467 -17486 -70
rect -17380 -467 -17374 -70
rect -17492 -479 -17374 -467
rect -17258 -70 -17140 -58
rect -17258 -467 -17252 -70
rect -17146 -467 -17140 -70
rect -17258 -479 -17140 -467
rect -17024 -70 -16906 -58
rect -17024 -467 -17018 -70
rect -16912 -467 -16906 -70
rect -17024 -479 -16906 -467
rect -16790 -70 -16672 -58
rect -16790 -467 -16784 -70
rect -16678 -467 -16672 -70
rect -16790 -479 -16672 -467
rect -16556 -70 -16438 -58
rect -16556 -467 -16550 -70
rect -16444 -467 -16438 -70
rect -16556 -479 -16438 -467
rect -16322 -70 -16204 -58
rect -16322 -467 -16316 -70
rect -16210 -467 -16204 -70
rect -16322 -479 -16204 -467
rect -16088 -70 -15970 -58
rect -16088 -467 -16082 -70
rect -15976 -467 -15970 -70
rect -16088 -479 -15970 -467
rect -15854 -70 -15736 -58
rect -15854 -467 -15848 -70
rect -15742 -467 -15736 -70
rect -15854 -479 -15736 -467
rect -15620 -70 -15502 -58
rect -15620 -467 -15614 -70
rect -15508 -467 -15502 -70
rect -15620 -479 -15502 -467
rect -15386 -70 -15268 -58
rect -15386 -467 -15380 -70
rect -15274 -467 -15268 -70
rect -15386 -479 -15268 -467
rect -15152 -70 -15034 -58
rect -15152 -467 -15146 -70
rect -15040 -467 -15034 -70
rect -15152 -479 -15034 -467
rect -14918 -70 -14800 -58
rect -14918 -467 -14912 -70
rect -14806 -467 -14800 -70
rect -14918 -479 -14800 -467
rect -14684 -70 -14566 -58
rect -14684 -467 -14678 -70
rect -14572 -467 -14566 -70
rect -14684 -479 -14566 -467
rect -14450 -70 -14332 -58
rect -14450 -467 -14444 -70
rect -14338 -467 -14332 -70
rect -14450 -479 -14332 -467
rect -14216 -70 -14098 -58
rect -14216 -467 -14210 -70
rect -14104 -467 -14098 -70
rect -14216 -479 -14098 -467
rect -13982 -70 -13864 -58
rect -13982 -467 -13976 -70
rect -13870 -467 -13864 -70
rect -13982 -479 -13864 -467
rect -13748 -70 -13630 -58
rect -13748 -467 -13742 -70
rect -13636 -467 -13630 -70
rect -13748 -479 -13630 -467
rect -13514 -70 -13396 -58
rect -13514 -467 -13508 -70
rect -13402 -467 -13396 -70
rect -13514 -479 -13396 -467
rect -13280 -70 -13162 -58
rect -13280 -467 -13274 -70
rect -13168 -467 -13162 -70
rect -13280 -479 -13162 -467
rect -13046 -70 -12928 -58
rect -13046 -467 -13040 -70
rect -12934 -467 -12928 -70
rect -13046 -479 -12928 -467
rect -12812 -70 -12694 -58
rect -12812 -467 -12806 -70
rect -12700 -467 -12694 -70
rect -12812 -479 -12694 -467
rect -12578 -70 -12460 -58
rect -12578 -467 -12572 -70
rect -12466 -467 -12460 -70
rect -12578 -479 -12460 -467
rect -12344 -70 -12226 -58
rect -12344 -467 -12338 -70
rect -12232 -467 -12226 -70
rect -12344 -479 -12226 -467
rect -12110 -70 -11992 -58
rect -12110 -467 -12104 -70
rect -11998 -467 -11992 -70
rect -12110 -479 -11992 -467
rect -11876 -70 -11758 -58
rect -11876 -467 -11870 -70
rect -11764 -467 -11758 -70
rect -11876 -479 -11758 -467
rect -11642 -70 -11524 -58
rect -11642 -467 -11636 -70
rect -11530 -467 -11524 -70
rect -11642 -479 -11524 -467
rect -11408 -70 -11290 -58
rect -11408 -467 -11402 -70
rect -11296 -467 -11290 -70
rect -11408 -479 -11290 -467
rect -11174 -70 -11056 -58
rect -11174 -467 -11168 -70
rect -11062 -467 -11056 -70
rect -11174 -479 -11056 -467
rect -10940 -70 -10822 -58
rect -10940 -467 -10934 -70
rect -10828 -467 -10822 -70
rect -10940 -479 -10822 -467
rect -10706 -70 -10588 -58
rect -10706 -467 -10700 -70
rect -10594 -467 -10588 -70
rect -10706 -479 -10588 -467
rect -10472 -70 -10354 -58
rect -10472 -467 -10466 -70
rect -10360 -467 -10354 -70
rect -10472 -479 -10354 -467
rect -10238 -70 -10120 -58
rect -10238 -467 -10232 -70
rect -10126 -467 -10120 -70
rect -10238 -479 -10120 -467
rect -10004 -70 -9886 -58
rect -10004 -467 -9998 -70
rect -9892 -467 -9886 -70
rect -10004 -479 -9886 -467
rect -9770 -70 -9652 -58
rect -9770 -467 -9764 -70
rect -9658 -467 -9652 -70
rect -9770 -479 -9652 -467
rect -9536 -70 -9418 -58
rect -9536 -467 -9530 -70
rect -9424 -467 -9418 -70
rect -9536 -479 -9418 -467
rect -9302 -70 -9184 -58
rect -9302 -467 -9296 -70
rect -9190 -467 -9184 -70
rect -9302 -479 -9184 -467
rect -9068 -70 -8950 -58
rect -9068 -467 -9062 -70
rect -8956 -467 -8950 -70
rect -9068 -479 -8950 -467
rect -8834 -70 -8716 -58
rect -8834 -467 -8828 -70
rect -8722 -467 -8716 -70
rect -8834 -479 -8716 -467
rect -8600 -70 -8482 -58
rect -8600 -467 -8594 -70
rect -8488 -467 -8482 -70
rect -8600 -479 -8482 -467
rect -8366 -70 -8248 -58
rect -8366 -467 -8360 -70
rect -8254 -467 -8248 -70
rect -8366 -479 -8248 -467
rect -8132 -70 -8014 -58
rect -8132 -467 -8126 -70
rect -8020 -467 -8014 -70
rect -8132 -479 -8014 -467
rect -7898 -70 -7780 -58
rect -7898 -467 -7892 -70
rect -7786 -467 -7780 -70
rect -7898 -479 -7780 -467
rect -7664 -70 -7546 -58
rect -7664 -467 -7658 -70
rect -7552 -467 -7546 -70
rect -7664 -479 -7546 -467
rect -7430 -70 -7312 -58
rect -7430 -467 -7424 -70
rect -7318 -467 -7312 -70
rect -7430 -479 -7312 -467
rect -7196 -70 -7078 -58
rect -7196 -467 -7190 -70
rect -7084 -467 -7078 -70
rect -7196 -479 -7078 -467
rect -6962 -70 -6844 -58
rect -6962 -467 -6956 -70
rect -6850 -467 -6844 -70
rect -6962 -479 -6844 -467
rect -6728 -70 -6610 -58
rect -6728 -467 -6722 -70
rect -6616 -467 -6610 -70
rect -6728 -479 -6610 -467
rect -6494 -70 -6376 -58
rect -6494 -467 -6488 -70
rect -6382 -467 -6376 -70
rect -6494 -479 -6376 -467
rect -6260 -70 -6142 -58
rect -6260 -467 -6254 -70
rect -6148 -467 -6142 -70
rect -6260 -479 -6142 -467
rect -6026 -70 -5908 -58
rect -6026 -467 -6020 -70
rect -5914 -467 -5908 -70
rect -6026 -479 -5908 -467
rect -5792 -70 -5674 -58
rect -5792 -467 -5786 -70
rect -5680 -467 -5674 -70
rect -5792 -479 -5674 -467
rect -5558 -70 -5440 -58
rect -5558 -467 -5552 -70
rect -5446 -467 -5440 -70
rect -5558 -479 -5440 -467
rect -5324 -70 -5206 -58
rect -5324 -467 -5318 -70
rect -5212 -467 -5206 -70
rect -5324 -479 -5206 -467
rect -5090 -70 -4972 -58
rect -5090 -467 -5084 -70
rect -4978 -467 -4972 -70
rect -5090 -479 -4972 -467
rect -4856 -70 -4738 -58
rect -4856 -467 -4850 -70
rect -4744 -467 -4738 -70
rect -4856 -479 -4738 -467
rect -4622 -70 -4504 -58
rect -4622 -467 -4616 -70
rect -4510 -467 -4504 -70
rect -4622 -479 -4504 -467
rect -4388 -70 -4270 -58
rect -4388 -467 -4382 -70
rect -4276 -467 -4270 -70
rect -4388 -479 -4270 -467
rect -4154 -70 -4036 -58
rect -4154 -467 -4148 -70
rect -4042 -467 -4036 -70
rect -4154 -479 -4036 -467
rect -3920 -70 -3802 -58
rect -3920 -467 -3914 -70
rect -3808 -467 -3802 -70
rect -3920 -479 -3802 -467
rect -3686 -70 -3568 -58
rect -3686 -467 -3680 -70
rect -3574 -467 -3568 -70
rect -3686 -479 -3568 -467
rect -3452 -70 -3334 -58
rect -3452 -467 -3446 -70
rect -3340 -467 -3334 -70
rect -3452 -479 -3334 -467
rect -3218 -70 -3100 -58
rect -3218 -467 -3212 -70
rect -3106 -467 -3100 -70
rect -3218 -479 -3100 -467
rect -2984 -70 -2866 -58
rect -2984 -467 -2978 -70
rect -2872 -467 -2866 -70
rect -2984 -479 -2866 -467
rect -2750 -70 -2632 -58
rect -2750 -467 -2744 -70
rect -2638 -467 -2632 -70
rect -2750 -479 -2632 -467
rect -2516 -70 -2398 -58
rect -2516 -467 -2510 -70
rect -2404 -467 -2398 -70
rect -2516 -479 -2398 -467
rect -2282 -70 -2164 -58
rect -2282 -467 -2276 -70
rect -2170 -467 -2164 -70
rect -2282 -479 -2164 -467
rect -2048 -70 -1930 -58
rect -2048 -467 -2042 -70
rect -1936 -467 -1930 -70
rect -2048 -479 -1930 -467
rect -1814 -70 -1696 -58
rect -1814 -467 -1808 -70
rect -1702 -467 -1696 -70
rect -1814 -479 -1696 -467
rect -1580 -70 -1462 -58
rect -1580 -467 -1574 -70
rect -1468 -467 -1462 -70
rect -1580 -479 -1462 -467
rect -1346 -70 -1228 -58
rect -1346 -467 -1340 -70
rect -1234 -467 -1228 -70
rect -1346 -479 -1228 -467
rect -1112 -70 -994 -58
rect -1112 -467 -1106 -70
rect -1000 -467 -994 -70
rect -1112 -479 -994 -467
rect -878 -70 -760 -58
rect -878 -467 -872 -70
rect -766 -467 -760 -70
rect -878 -479 -760 -467
rect -644 -70 -526 -58
rect -644 -467 -638 -70
rect -532 -467 -526 -70
rect -644 -479 -526 -467
rect -410 -70 -292 -58
rect -410 -467 -404 -70
rect -298 -467 -292 -70
rect -410 -479 -292 -467
rect -176 -70 -58 -58
rect -176 -467 -170 -70
rect -64 -467 -58 -70
rect -176 -479 -58 -467
rect 58 -70 176 -58
rect 58 -467 64 -70
rect 170 -467 176 -70
rect 58 -479 176 -467
rect 292 -70 410 -58
rect 292 -467 298 -70
rect 404 -467 410 -70
rect 292 -479 410 -467
rect 526 -70 644 -58
rect 526 -467 532 -70
rect 638 -467 644 -70
rect 526 -479 644 -467
rect 760 -70 878 -58
rect 760 -467 766 -70
rect 872 -467 878 -70
rect 760 -479 878 -467
rect 994 -70 1112 -58
rect 994 -467 1000 -70
rect 1106 -467 1112 -70
rect 994 -479 1112 -467
rect 1228 -70 1346 -58
rect 1228 -467 1234 -70
rect 1340 -467 1346 -70
rect 1228 -479 1346 -467
rect 1462 -70 1580 -58
rect 1462 -467 1468 -70
rect 1574 -467 1580 -70
rect 1462 -479 1580 -467
rect 1696 -70 1814 -58
rect 1696 -467 1702 -70
rect 1808 -467 1814 -70
rect 1696 -479 1814 -467
rect 1930 -70 2048 -58
rect 1930 -467 1936 -70
rect 2042 -467 2048 -70
rect 1930 -479 2048 -467
rect 2164 -70 2282 -58
rect 2164 -467 2170 -70
rect 2276 -467 2282 -70
rect 2164 -479 2282 -467
rect 2398 -70 2516 -58
rect 2398 -467 2404 -70
rect 2510 -467 2516 -70
rect 2398 -479 2516 -467
rect 2632 -70 2750 -58
rect 2632 -467 2638 -70
rect 2744 -467 2750 -70
rect 2632 -479 2750 -467
rect 2866 -70 2984 -58
rect 2866 -467 2872 -70
rect 2978 -467 2984 -70
rect 2866 -479 2984 -467
rect 3100 -70 3218 -58
rect 3100 -467 3106 -70
rect 3212 -467 3218 -70
rect 3100 -479 3218 -467
rect 3334 -70 3452 -58
rect 3334 -467 3340 -70
rect 3446 -467 3452 -70
rect 3334 -479 3452 -467
rect 3568 -70 3686 -58
rect 3568 -467 3574 -70
rect 3680 -467 3686 -70
rect 3568 -479 3686 -467
rect 3802 -70 3920 -58
rect 3802 -467 3808 -70
rect 3914 -467 3920 -70
rect 3802 -479 3920 -467
rect 4036 -70 4154 -58
rect 4036 -467 4042 -70
rect 4148 -467 4154 -70
rect 4036 -479 4154 -467
rect 4270 -70 4388 -58
rect 4270 -467 4276 -70
rect 4382 -467 4388 -70
rect 4270 -479 4388 -467
rect 4504 -70 4622 -58
rect 4504 -467 4510 -70
rect 4616 -467 4622 -70
rect 4504 -479 4622 -467
rect 4738 -70 4856 -58
rect 4738 -467 4744 -70
rect 4850 -467 4856 -70
rect 4738 -479 4856 -467
rect 4972 -70 5090 -58
rect 4972 -467 4978 -70
rect 5084 -467 5090 -70
rect 4972 -479 5090 -467
rect 5206 -70 5324 -58
rect 5206 -467 5212 -70
rect 5318 -467 5324 -70
rect 5206 -479 5324 -467
rect 5440 -70 5558 -58
rect 5440 -467 5446 -70
rect 5552 -467 5558 -70
rect 5440 -479 5558 -467
rect 5674 -70 5792 -58
rect 5674 -467 5680 -70
rect 5786 -467 5792 -70
rect 5674 -479 5792 -467
rect 5908 -70 6026 -58
rect 5908 -467 5914 -70
rect 6020 -467 6026 -70
rect 5908 -479 6026 -467
rect 6142 -70 6260 -58
rect 6142 -467 6148 -70
rect 6254 -467 6260 -70
rect 6142 -479 6260 -467
rect 6376 -70 6494 -58
rect 6376 -467 6382 -70
rect 6488 -467 6494 -70
rect 6376 -479 6494 -467
rect 6610 -70 6728 -58
rect 6610 -467 6616 -70
rect 6722 -467 6728 -70
rect 6610 -479 6728 -467
rect 6844 -70 6962 -58
rect 6844 -467 6850 -70
rect 6956 -467 6962 -70
rect 6844 -479 6962 -467
rect 7078 -70 7196 -58
rect 7078 -467 7084 -70
rect 7190 -467 7196 -70
rect 7078 -479 7196 -467
rect 7312 -70 7430 -58
rect 7312 -467 7318 -70
rect 7424 -467 7430 -70
rect 7312 -479 7430 -467
rect 7546 -70 7664 -58
rect 7546 -467 7552 -70
rect 7658 -467 7664 -70
rect 7546 -479 7664 -467
rect 7780 -70 7898 -58
rect 7780 -467 7786 -70
rect 7892 -467 7898 -70
rect 7780 -479 7898 -467
rect 8014 -70 8132 -58
rect 8014 -467 8020 -70
rect 8126 -467 8132 -70
rect 8014 -479 8132 -467
rect 8248 -70 8366 -58
rect 8248 -467 8254 -70
rect 8360 -467 8366 -70
rect 8248 -479 8366 -467
rect 8482 -70 8600 -58
rect 8482 -467 8488 -70
rect 8594 -467 8600 -70
rect 8482 -479 8600 -467
rect 8716 -70 8834 -58
rect 8716 -467 8722 -70
rect 8828 -467 8834 -70
rect 8716 -479 8834 -467
rect 8950 -70 9068 -58
rect 8950 -467 8956 -70
rect 9062 -467 9068 -70
rect 8950 -479 9068 -467
rect 9184 -70 9302 -58
rect 9184 -467 9190 -70
rect 9296 -467 9302 -70
rect 9184 -479 9302 -467
rect 9418 -70 9536 -58
rect 9418 -467 9424 -70
rect 9530 -467 9536 -70
rect 9418 -479 9536 -467
rect 9652 -70 9770 -58
rect 9652 -467 9658 -70
rect 9764 -467 9770 -70
rect 9652 -479 9770 -467
rect 9886 -70 10004 -58
rect 9886 -467 9892 -70
rect 9998 -467 10004 -70
rect 9886 -479 10004 -467
rect 10120 -70 10238 -58
rect 10120 -467 10126 -70
rect 10232 -467 10238 -70
rect 10120 -479 10238 -467
rect 10354 -70 10472 -58
rect 10354 -467 10360 -70
rect 10466 -467 10472 -70
rect 10354 -479 10472 -467
rect 10588 -70 10706 -58
rect 10588 -467 10594 -70
rect 10700 -467 10706 -70
rect 10588 -479 10706 -467
rect 10822 -70 10940 -58
rect 10822 -467 10828 -70
rect 10934 -467 10940 -70
rect 10822 -479 10940 -467
rect 11056 -70 11174 -58
rect 11056 -467 11062 -70
rect 11168 -467 11174 -70
rect 11056 -479 11174 -467
rect 11290 -70 11408 -58
rect 11290 -467 11296 -70
rect 11402 -467 11408 -70
rect 11290 -479 11408 -467
rect 11524 -70 11642 -58
rect 11524 -467 11530 -70
rect 11636 -467 11642 -70
rect 11524 -479 11642 -467
rect 11758 -70 11876 -58
rect 11758 -467 11764 -70
rect 11870 -467 11876 -70
rect 11758 -479 11876 -467
rect 11992 -70 12110 -58
rect 11992 -467 11998 -70
rect 12104 -467 12110 -70
rect 11992 -479 12110 -467
rect 12226 -70 12344 -58
rect 12226 -467 12232 -70
rect 12338 -467 12344 -70
rect 12226 -479 12344 -467
rect 12460 -70 12578 -58
rect 12460 -467 12466 -70
rect 12572 -467 12578 -70
rect 12460 -479 12578 -467
rect 12694 -70 12812 -58
rect 12694 -467 12700 -70
rect 12806 -467 12812 -70
rect 12694 -479 12812 -467
rect 12928 -70 13046 -58
rect 12928 -467 12934 -70
rect 13040 -467 13046 -70
rect 12928 -479 13046 -467
rect 13162 -70 13280 -58
rect 13162 -467 13168 -70
rect 13274 -467 13280 -70
rect 13162 -479 13280 -467
rect 13396 -70 13514 -58
rect 13396 -467 13402 -70
rect 13508 -467 13514 -70
rect 13396 -479 13514 -467
rect 13630 -70 13748 -58
rect 13630 -467 13636 -70
rect 13742 -467 13748 -70
rect 13630 -479 13748 -467
rect 13864 -70 13982 -58
rect 13864 -467 13870 -70
rect 13976 -467 13982 -70
rect 13864 -479 13982 -467
rect 14098 -70 14216 -58
rect 14098 -467 14104 -70
rect 14210 -467 14216 -70
rect 14098 -479 14216 -467
rect 14332 -70 14450 -58
rect 14332 -467 14338 -70
rect 14444 -467 14450 -70
rect 14332 -479 14450 -467
rect 14566 -70 14684 -58
rect 14566 -467 14572 -70
rect 14678 -467 14684 -70
rect 14566 -479 14684 -467
rect 14800 -70 14918 -58
rect 14800 -467 14806 -70
rect 14912 -467 14918 -70
rect 14800 -479 14918 -467
rect 15034 -70 15152 -58
rect 15034 -467 15040 -70
rect 15146 -467 15152 -70
rect 15034 -479 15152 -467
rect 15268 -70 15386 -58
rect 15268 -467 15274 -70
rect 15380 -467 15386 -70
rect 15268 -479 15386 -467
rect 15502 -70 15620 -58
rect 15502 -467 15508 -70
rect 15614 -467 15620 -70
rect 15502 -479 15620 -467
rect 15736 -70 15854 -58
rect 15736 -467 15742 -70
rect 15848 -467 15854 -70
rect 15736 -479 15854 -467
rect 15970 -70 16088 -58
rect 15970 -467 15976 -70
rect 16082 -467 16088 -70
rect 15970 -479 16088 -467
rect 16204 -70 16322 -58
rect 16204 -467 16210 -70
rect 16316 -467 16322 -70
rect 16204 -479 16322 -467
rect 16438 -70 16556 -58
rect 16438 -467 16444 -70
rect 16550 -467 16556 -70
rect 16438 -479 16556 -467
rect 16672 -70 16790 -58
rect 16672 -467 16678 -70
rect 16784 -467 16790 -70
rect 16672 -479 16790 -467
rect 16906 -70 17024 -58
rect 16906 -467 16912 -70
rect 17018 -467 17024 -70
rect 16906 -479 17024 -467
rect 17140 -70 17258 -58
rect 17140 -467 17146 -70
rect 17252 -467 17258 -70
rect 17140 -479 17258 -467
rect 17374 -70 17492 -58
rect 17374 -467 17380 -70
rect 17486 -467 17492 -70
rect 17374 -479 17492 -467
rect 17608 -70 17726 -58
rect 17608 -467 17614 -70
rect 17720 -467 17726 -70
rect 17608 -479 17726 -467
rect 17842 -70 17960 -58
rect 17842 -467 17848 -70
rect 17954 -467 17960 -70
rect 17842 -479 17960 -467
rect 18076 -70 18194 -58
rect 18076 -467 18082 -70
rect 18188 -467 18194 -70
rect 18076 -479 18194 -467
rect 18310 -70 18428 -58
rect 18310 -467 18316 -70
rect 18422 -467 18428 -70
rect 18310 -479 18428 -467
rect 18544 -70 18662 -58
rect 18544 -467 18550 -70
rect 18656 -467 18662 -70
rect 18544 -479 18662 -467
rect 18778 -70 18896 -58
rect 18778 -467 18784 -70
rect 18890 -467 18896 -70
rect 18778 -479 18896 -467
rect 19012 -70 19130 -58
rect 19012 -467 19018 -70
rect 19124 -467 19130 -70
rect 19012 -479 19130 -467
rect 19246 -70 19364 -58
rect 19246 -467 19252 -70
rect 19358 -467 19364 -70
rect 19246 -479 19364 -467
rect 19480 -70 19598 -58
rect 19480 -467 19486 -70
rect 19592 -467 19598 -70
rect 19480 -479 19598 -467
rect 19714 -70 19832 -58
rect 19714 -467 19720 -70
rect 19826 -467 19832 -70
rect 19714 -479 19832 -467
rect 19948 -70 20066 -58
rect 19948 -467 19954 -70
rect 20060 -467 20066 -70
rect 19948 -479 20066 -467
rect 20182 -70 20300 -58
rect 20182 -467 20188 -70
rect 20294 -467 20300 -70
rect 20182 -479 20300 -467
rect 20416 -70 20534 -58
rect 20416 -467 20422 -70
rect 20528 -467 20534 -70
rect 20416 -479 20534 -467
rect 20650 -70 20768 -58
rect 20650 -467 20656 -70
rect 20762 -467 20768 -70
rect 20650 -479 20768 -467
rect 20884 -70 21002 -58
rect 20884 -467 20890 -70
rect 20996 -467 21002 -70
rect 20884 -479 21002 -467
rect 21118 -70 21236 -58
rect 21118 -467 21124 -70
rect 21230 -467 21236 -70
rect 21118 -479 21236 -467
rect 21352 -70 21470 -58
rect 21352 -467 21358 -70
rect 21464 -467 21470 -70
rect 21352 -479 21470 -467
rect 21586 -70 21704 -58
rect 21586 -467 21592 -70
rect 21698 -467 21704 -70
rect 21586 -479 21704 -467
rect 21820 -70 21938 -58
rect 21820 -467 21826 -70
rect 21932 -467 21938 -70
rect 21820 -479 21938 -467
rect 22054 -70 22172 -58
rect 22054 -467 22060 -70
rect 22166 -467 22172 -70
rect 22054 -479 22172 -467
rect 22288 -70 22406 -58
rect 22288 -467 22294 -70
rect 22400 -467 22406 -70
rect 22288 -479 22406 -467
rect 22522 -70 22640 -58
rect 22522 -467 22528 -70
rect 22634 -467 22640 -70
rect 22522 -479 22640 -467
rect 22756 -70 22874 -58
rect 22756 -467 22762 -70
rect 22868 -467 22874 -70
rect 22756 -479 22874 -467
rect 22990 -70 23108 -58
rect 22990 -467 22996 -70
rect 23102 -467 23108 -70
rect 22990 -479 23108 -467
rect 23224 -70 23342 -58
rect 23224 -467 23230 -70
rect 23336 -467 23342 -70
rect 23224 -479 23342 -467
rect 23458 -70 23576 -58
rect 23458 -467 23464 -70
rect 23570 -467 23576 -70
rect 23458 -479 23576 -467
rect 23692 -70 23810 -58
rect 23692 -467 23698 -70
rect 23804 -467 23810 -70
rect 23692 -479 23810 -467
rect 23926 -70 24044 -58
rect 23926 -467 23932 -70
rect 24038 -467 24044 -70
rect 23926 -479 24044 -467
rect 24160 -70 24278 -58
rect 24160 -467 24166 -70
rect 24272 -467 24278 -70
rect 24160 -479 24278 -467
rect 24394 -70 24512 -58
rect 24394 -467 24400 -70
rect 24506 -467 24512 -70
rect 24394 -479 24512 -467
rect 24628 -70 24746 -58
rect 24628 -467 24634 -70
rect 24740 -467 24746 -70
rect 24628 -479 24746 -467
rect 24862 -70 24980 -58
rect 24862 -467 24868 -70
rect 24974 -467 24980 -70
rect 24862 -479 24980 -467
rect 25096 -70 25214 -58
rect 25096 -467 25102 -70
rect 25208 -467 25214 -70
rect 25096 -479 25214 -467
rect 25330 -70 25448 -58
rect 25330 -467 25336 -70
rect 25442 -467 25448 -70
rect 25330 -479 25448 -467
rect 25564 -70 25682 -58
rect 25564 -467 25570 -70
rect 25676 -467 25682 -70
rect 25564 -479 25682 -467
rect 25798 -70 25916 -58
rect 25798 -467 25804 -70
rect 25910 -467 25916 -70
rect 25798 -479 25916 -467
rect 26032 -70 26150 -58
rect 26032 -467 26038 -70
rect 26144 -467 26150 -70
rect 26032 -479 26150 -467
rect 26266 -70 26384 -58
rect 26266 -467 26272 -70
rect 26378 -467 26384 -70
rect 26266 -479 26384 -467
rect 26500 -70 26618 -58
rect 26500 -467 26506 -70
rect 26612 -467 26618 -70
rect 26500 -479 26618 -467
rect 26734 -70 26852 -58
rect 26734 -467 26740 -70
rect 26846 -467 26852 -70
rect 26734 -479 26852 -467
rect 26968 -70 27086 -58
rect 26968 -467 26974 -70
rect 27080 -467 27086 -70
rect 26968 -479 27086 -467
rect 27202 -70 27320 -58
rect 27202 -467 27208 -70
rect 27314 -467 27320 -70
rect 27202 -479 27320 -467
rect 27436 -70 27554 -58
rect 27436 -467 27442 -70
rect 27548 -467 27554 -70
rect 27436 -479 27554 -467
rect 27670 -70 27788 -58
rect 27670 -467 27676 -70
rect 27782 -467 27788 -70
rect 27670 -479 27788 -467
rect 27904 -70 28022 -58
rect 27904 -467 27910 -70
rect 28016 -467 28022 -70
rect 27904 -479 28022 -467
rect 28138 -70 28256 -58
rect 28138 -467 28144 -70
rect 28250 -467 28256 -70
rect 28138 -479 28256 -467
rect 28372 -70 28490 -58
rect 28372 -467 28378 -70
rect 28484 -467 28490 -70
rect 28372 -479 28490 -467
rect 28606 -70 28724 -58
rect 28606 -467 28612 -70
rect 28718 -467 28724 -70
rect 28606 -479 28724 -467
rect 28840 -70 28958 -58
rect 28840 -467 28846 -70
rect 28952 -467 28958 -70
rect 28840 -479 28958 -467
rect 29074 -70 29192 -58
rect 29074 -467 29080 -70
rect 29186 -467 29192 -70
rect 29074 -479 29192 -467
rect 29308 -70 29426 -58
rect 29308 -467 29314 -70
rect 29420 -467 29426 -70
rect 29308 -479 29426 -467
rect 29542 -70 29660 -58
rect 29542 -467 29548 -70
rect 29654 -467 29660 -70
rect 29542 -479 29660 -467
rect 29776 -70 29894 -58
rect 29776 -467 29782 -70
rect 29888 -467 29894 -70
rect 29776 -479 29894 -467
rect -29894 -5469 -29776 -5457
rect -29894 -5866 -29888 -5469
rect -29782 -5866 -29776 -5469
rect -29894 -5878 -29776 -5866
rect -29660 -5469 -29542 -5457
rect -29660 -5866 -29654 -5469
rect -29548 -5866 -29542 -5469
rect -29660 -5878 -29542 -5866
rect -29426 -5469 -29308 -5457
rect -29426 -5866 -29420 -5469
rect -29314 -5866 -29308 -5469
rect -29426 -5878 -29308 -5866
rect -29192 -5469 -29074 -5457
rect -29192 -5866 -29186 -5469
rect -29080 -5866 -29074 -5469
rect -29192 -5878 -29074 -5866
rect -28958 -5469 -28840 -5457
rect -28958 -5866 -28952 -5469
rect -28846 -5866 -28840 -5469
rect -28958 -5878 -28840 -5866
rect -28724 -5469 -28606 -5457
rect -28724 -5866 -28718 -5469
rect -28612 -5866 -28606 -5469
rect -28724 -5878 -28606 -5866
rect -28490 -5469 -28372 -5457
rect -28490 -5866 -28484 -5469
rect -28378 -5866 -28372 -5469
rect -28490 -5878 -28372 -5866
rect -28256 -5469 -28138 -5457
rect -28256 -5866 -28250 -5469
rect -28144 -5866 -28138 -5469
rect -28256 -5878 -28138 -5866
rect -28022 -5469 -27904 -5457
rect -28022 -5866 -28016 -5469
rect -27910 -5866 -27904 -5469
rect -28022 -5878 -27904 -5866
rect -27788 -5469 -27670 -5457
rect -27788 -5866 -27782 -5469
rect -27676 -5866 -27670 -5469
rect -27788 -5878 -27670 -5866
rect -27554 -5469 -27436 -5457
rect -27554 -5866 -27548 -5469
rect -27442 -5866 -27436 -5469
rect -27554 -5878 -27436 -5866
rect -27320 -5469 -27202 -5457
rect -27320 -5866 -27314 -5469
rect -27208 -5866 -27202 -5469
rect -27320 -5878 -27202 -5866
rect -27086 -5469 -26968 -5457
rect -27086 -5866 -27080 -5469
rect -26974 -5866 -26968 -5469
rect -27086 -5878 -26968 -5866
rect -26852 -5469 -26734 -5457
rect -26852 -5866 -26846 -5469
rect -26740 -5866 -26734 -5469
rect -26852 -5878 -26734 -5866
rect -26618 -5469 -26500 -5457
rect -26618 -5866 -26612 -5469
rect -26506 -5866 -26500 -5469
rect -26618 -5878 -26500 -5866
rect -26384 -5469 -26266 -5457
rect -26384 -5866 -26378 -5469
rect -26272 -5866 -26266 -5469
rect -26384 -5878 -26266 -5866
rect -26150 -5469 -26032 -5457
rect -26150 -5866 -26144 -5469
rect -26038 -5866 -26032 -5469
rect -26150 -5878 -26032 -5866
rect -25916 -5469 -25798 -5457
rect -25916 -5866 -25910 -5469
rect -25804 -5866 -25798 -5469
rect -25916 -5878 -25798 -5866
rect -25682 -5469 -25564 -5457
rect -25682 -5866 -25676 -5469
rect -25570 -5866 -25564 -5469
rect -25682 -5878 -25564 -5866
rect -25448 -5469 -25330 -5457
rect -25448 -5866 -25442 -5469
rect -25336 -5866 -25330 -5469
rect -25448 -5878 -25330 -5866
rect -25214 -5469 -25096 -5457
rect -25214 -5866 -25208 -5469
rect -25102 -5866 -25096 -5469
rect -25214 -5878 -25096 -5866
rect -24980 -5469 -24862 -5457
rect -24980 -5866 -24974 -5469
rect -24868 -5866 -24862 -5469
rect -24980 -5878 -24862 -5866
rect -24746 -5469 -24628 -5457
rect -24746 -5866 -24740 -5469
rect -24634 -5866 -24628 -5469
rect -24746 -5878 -24628 -5866
rect -24512 -5469 -24394 -5457
rect -24512 -5866 -24506 -5469
rect -24400 -5866 -24394 -5469
rect -24512 -5878 -24394 -5866
rect -24278 -5469 -24160 -5457
rect -24278 -5866 -24272 -5469
rect -24166 -5866 -24160 -5469
rect -24278 -5878 -24160 -5866
rect -24044 -5469 -23926 -5457
rect -24044 -5866 -24038 -5469
rect -23932 -5866 -23926 -5469
rect -24044 -5878 -23926 -5866
rect -23810 -5469 -23692 -5457
rect -23810 -5866 -23804 -5469
rect -23698 -5866 -23692 -5469
rect -23810 -5878 -23692 -5866
rect -23576 -5469 -23458 -5457
rect -23576 -5866 -23570 -5469
rect -23464 -5866 -23458 -5469
rect -23576 -5878 -23458 -5866
rect -23342 -5469 -23224 -5457
rect -23342 -5866 -23336 -5469
rect -23230 -5866 -23224 -5469
rect -23342 -5878 -23224 -5866
rect -23108 -5469 -22990 -5457
rect -23108 -5866 -23102 -5469
rect -22996 -5866 -22990 -5469
rect -23108 -5878 -22990 -5866
rect -22874 -5469 -22756 -5457
rect -22874 -5866 -22868 -5469
rect -22762 -5866 -22756 -5469
rect -22874 -5878 -22756 -5866
rect -22640 -5469 -22522 -5457
rect -22640 -5866 -22634 -5469
rect -22528 -5866 -22522 -5469
rect -22640 -5878 -22522 -5866
rect -22406 -5469 -22288 -5457
rect -22406 -5866 -22400 -5469
rect -22294 -5866 -22288 -5469
rect -22406 -5878 -22288 -5866
rect -22172 -5469 -22054 -5457
rect -22172 -5866 -22166 -5469
rect -22060 -5866 -22054 -5469
rect -22172 -5878 -22054 -5866
rect -21938 -5469 -21820 -5457
rect -21938 -5866 -21932 -5469
rect -21826 -5866 -21820 -5469
rect -21938 -5878 -21820 -5866
rect -21704 -5469 -21586 -5457
rect -21704 -5866 -21698 -5469
rect -21592 -5866 -21586 -5469
rect -21704 -5878 -21586 -5866
rect -21470 -5469 -21352 -5457
rect -21470 -5866 -21464 -5469
rect -21358 -5866 -21352 -5469
rect -21470 -5878 -21352 -5866
rect -21236 -5469 -21118 -5457
rect -21236 -5866 -21230 -5469
rect -21124 -5866 -21118 -5469
rect -21236 -5878 -21118 -5866
rect -21002 -5469 -20884 -5457
rect -21002 -5866 -20996 -5469
rect -20890 -5866 -20884 -5469
rect -21002 -5878 -20884 -5866
rect -20768 -5469 -20650 -5457
rect -20768 -5866 -20762 -5469
rect -20656 -5866 -20650 -5469
rect -20768 -5878 -20650 -5866
rect -20534 -5469 -20416 -5457
rect -20534 -5866 -20528 -5469
rect -20422 -5866 -20416 -5469
rect -20534 -5878 -20416 -5866
rect -20300 -5469 -20182 -5457
rect -20300 -5866 -20294 -5469
rect -20188 -5866 -20182 -5469
rect -20300 -5878 -20182 -5866
rect -20066 -5469 -19948 -5457
rect -20066 -5866 -20060 -5469
rect -19954 -5866 -19948 -5469
rect -20066 -5878 -19948 -5866
rect -19832 -5469 -19714 -5457
rect -19832 -5866 -19826 -5469
rect -19720 -5866 -19714 -5469
rect -19832 -5878 -19714 -5866
rect -19598 -5469 -19480 -5457
rect -19598 -5866 -19592 -5469
rect -19486 -5866 -19480 -5469
rect -19598 -5878 -19480 -5866
rect -19364 -5469 -19246 -5457
rect -19364 -5866 -19358 -5469
rect -19252 -5866 -19246 -5469
rect -19364 -5878 -19246 -5866
rect -19130 -5469 -19012 -5457
rect -19130 -5866 -19124 -5469
rect -19018 -5866 -19012 -5469
rect -19130 -5878 -19012 -5866
rect -18896 -5469 -18778 -5457
rect -18896 -5866 -18890 -5469
rect -18784 -5866 -18778 -5469
rect -18896 -5878 -18778 -5866
rect -18662 -5469 -18544 -5457
rect -18662 -5866 -18656 -5469
rect -18550 -5866 -18544 -5469
rect -18662 -5878 -18544 -5866
rect -18428 -5469 -18310 -5457
rect -18428 -5866 -18422 -5469
rect -18316 -5866 -18310 -5469
rect -18428 -5878 -18310 -5866
rect -18194 -5469 -18076 -5457
rect -18194 -5866 -18188 -5469
rect -18082 -5866 -18076 -5469
rect -18194 -5878 -18076 -5866
rect -17960 -5469 -17842 -5457
rect -17960 -5866 -17954 -5469
rect -17848 -5866 -17842 -5469
rect -17960 -5878 -17842 -5866
rect -17726 -5469 -17608 -5457
rect -17726 -5866 -17720 -5469
rect -17614 -5866 -17608 -5469
rect -17726 -5878 -17608 -5866
rect -17492 -5469 -17374 -5457
rect -17492 -5866 -17486 -5469
rect -17380 -5866 -17374 -5469
rect -17492 -5878 -17374 -5866
rect -17258 -5469 -17140 -5457
rect -17258 -5866 -17252 -5469
rect -17146 -5866 -17140 -5469
rect -17258 -5878 -17140 -5866
rect -17024 -5469 -16906 -5457
rect -17024 -5866 -17018 -5469
rect -16912 -5866 -16906 -5469
rect -17024 -5878 -16906 -5866
rect -16790 -5469 -16672 -5457
rect -16790 -5866 -16784 -5469
rect -16678 -5866 -16672 -5469
rect -16790 -5878 -16672 -5866
rect -16556 -5469 -16438 -5457
rect -16556 -5866 -16550 -5469
rect -16444 -5866 -16438 -5469
rect -16556 -5878 -16438 -5866
rect -16322 -5469 -16204 -5457
rect -16322 -5866 -16316 -5469
rect -16210 -5866 -16204 -5469
rect -16322 -5878 -16204 -5866
rect -16088 -5469 -15970 -5457
rect -16088 -5866 -16082 -5469
rect -15976 -5866 -15970 -5469
rect -16088 -5878 -15970 -5866
rect -15854 -5469 -15736 -5457
rect -15854 -5866 -15848 -5469
rect -15742 -5866 -15736 -5469
rect -15854 -5878 -15736 -5866
rect -15620 -5469 -15502 -5457
rect -15620 -5866 -15614 -5469
rect -15508 -5866 -15502 -5469
rect -15620 -5878 -15502 -5866
rect -15386 -5469 -15268 -5457
rect -15386 -5866 -15380 -5469
rect -15274 -5866 -15268 -5469
rect -15386 -5878 -15268 -5866
rect -15152 -5469 -15034 -5457
rect -15152 -5866 -15146 -5469
rect -15040 -5866 -15034 -5469
rect -15152 -5878 -15034 -5866
rect -14918 -5469 -14800 -5457
rect -14918 -5866 -14912 -5469
rect -14806 -5866 -14800 -5469
rect -14918 -5878 -14800 -5866
rect -14684 -5469 -14566 -5457
rect -14684 -5866 -14678 -5469
rect -14572 -5866 -14566 -5469
rect -14684 -5878 -14566 -5866
rect -14450 -5469 -14332 -5457
rect -14450 -5866 -14444 -5469
rect -14338 -5866 -14332 -5469
rect -14450 -5878 -14332 -5866
rect -14216 -5469 -14098 -5457
rect -14216 -5866 -14210 -5469
rect -14104 -5866 -14098 -5469
rect -14216 -5878 -14098 -5866
rect -13982 -5469 -13864 -5457
rect -13982 -5866 -13976 -5469
rect -13870 -5866 -13864 -5469
rect -13982 -5878 -13864 -5866
rect -13748 -5469 -13630 -5457
rect -13748 -5866 -13742 -5469
rect -13636 -5866 -13630 -5469
rect -13748 -5878 -13630 -5866
rect -13514 -5469 -13396 -5457
rect -13514 -5866 -13508 -5469
rect -13402 -5866 -13396 -5469
rect -13514 -5878 -13396 -5866
rect -13280 -5469 -13162 -5457
rect -13280 -5866 -13274 -5469
rect -13168 -5866 -13162 -5469
rect -13280 -5878 -13162 -5866
rect -13046 -5469 -12928 -5457
rect -13046 -5866 -13040 -5469
rect -12934 -5866 -12928 -5469
rect -13046 -5878 -12928 -5866
rect -12812 -5469 -12694 -5457
rect -12812 -5866 -12806 -5469
rect -12700 -5866 -12694 -5469
rect -12812 -5878 -12694 -5866
rect -12578 -5469 -12460 -5457
rect -12578 -5866 -12572 -5469
rect -12466 -5866 -12460 -5469
rect -12578 -5878 -12460 -5866
rect -12344 -5469 -12226 -5457
rect -12344 -5866 -12338 -5469
rect -12232 -5866 -12226 -5469
rect -12344 -5878 -12226 -5866
rect -12110 -5469 -11992 -5457
rect -12110 -5866 -12104 -5469
rect -11998 -5866 -11992 -5469
rect -12110 -5878 -11992 -5866
rect -11876 -5469 -11758 -5457
rect -11876 -5866 -11870 -5469
rect -11764 -5866 -11758 -5469
rect -11876 -5878 -11758 -5866
rect -11642 -5469 -11524 -5457
rect -11642 -5866 -11636 -5469
rect -11530 -5866 -11524 -5469
rect -11642 -5878 -11524 -5866
rect -11408 -5469 -11290 -5457
rect -11408 -5866 -11402 -5469
rect -11296 -5866 -11290 -5469
rect -11408 -5878 -11290 -5866
rect -11174 -5469 -11056 -5457
rect -11174 -5866 -11168 -5469
rect -11062 -5866 -11056 -5469
rect -11174 -5878 -11056 -5866
rect -10940 -5469 -10822 -5457
rect -10940 -5866 -10934 -5469
rect -10828 -5866 -10822 -5469
rect -10940 -5878 -10822 -5866
rect -10706 -5469 -10588 -5457
rect -10706 -5866 -10700 -5469
rect -10594 -5866 -10588 -5469
rect -10706 -5878 -10588 -5866
rect -10472 -5469 -10354 -5457
rect -10472 -5866 -10466 -5469
rect -10360 -5866 -10354 -5469
rect -10472 -5878 -10354 -5866
rect -10238 -5469 -10120 -5457
rect -10238 -5866 -10232 -5469
rect -10126 -5866 -10120 -5469
rect -10238 -5878 -10120 -5866
rect -10004 -5469 -9886 -5457
rect -10004 -5866 -9998 -5469
rect -9892 -5866 -9886 -5469
rect -10004 -5878 -9886 -5866
rect -9770 -5469 -9652 -5457
rect -9770 -5866 -9764 -5469
rect -9658 -5866 -9652 -5469
rect -9770 -5878 -9652 -5866
rect -9536 -5469 -9418 -5457
rect -9536 -5866 -9530 -5469
rect -9424 -5866 -9418 -5469
rect -9536 -5878 -9418 -5866
rect -9302 -5469 -9184 -5457
rect -9302 -5866 -9296 -5469
rect -9190 -5866 -9184 -5469
rect -9302 -5878 -9184 -5866
rect -9068 -5469 -8950 -5457
rect -9068 -5866 -9062 -5469
rect -8956 -5866 -8950 -5469
rect -9068 -5878 -8950 -5866
rect -8834 -5469 -8716 -5457
rect -8834 -5866 -8828 -5469
rect -8722 -5866 -8716 -5469
rect -8834 -5878 -8716 -5866
rect -8600 -5469 -8482 -5457
rect -8600 -5866 -8594 -5469
rect -8488 -5866 -8482 -5469
rect -8600 -5878 -8482 -5866
rect -8366 -5469 -8248 -5457
rect -8366 -5866 -8360 -5469
rect -8254 -5866 -8248 -5469
rect -8366 -5878 -8248 -5866
rect -8132 -5469 -8014 -5457
rect -8132 -5866 -8126 -5469
rect -8020 -5866 -8014 -5469
rect -8132 -5878 -8014 -5866
rect -7898 -5469 -7780 -5457
rect -7898 -5866 -7892 -5469
rect -7786 -5866 -7780 -5469
rect -7898 -5878 -7780 -5866
rect -7664 -5469 -7546 -5457
rect -7664 -5866 -7658 -5469
rect -7552 -5866 -7546 -5469
rect -7664 -5878 -7546 -5866
rect -7430 -5469 -7312 -5457
rect -7430 -5866 -7424 -5469
rect -7318 -5866 -7312 -5469
rect -7430 -5878 -7312 -5866
rect -7196 -5469 -7078 -5457
rect -7196 -5866 -7190 -5469
rect -7084 -5866 -7078 -5469
rect -7196 -5878 -7078 -5866
rect -6962 -5469 -6844 -5457
rect -6962 -5866 -6956 -5469
rect -6850 -5866 -6844 -5469
rect -6962 -5878 -6844 -5866
rect -6728 -5469 -6610 -5457
rect -6728 -5866 -6722 -5469
rect -6616 -5866 -6610 -5469
rect -6728 -5878 -6610 -5866
rect -6494 -5469 -6376 -5457
rect -6494 -5866 -6488 -5469
rect -6382 -5866 -6376 -5469
rect -6494 -5878 -6376 -5866
rect -6260 -5469 -6142 -5457
rect -6260 -5866 -6254 -5469
rect -6148 -5866 -6142 -5469
rect -6260 -5878 -6142 -5866
rect -6026 -5469 -5908 -5457
rect -6026 -5866 -6020 -5469
rect -5914 -5866 -5908 -5469
rect -6026 -5878 -5908 -5866
rect -5792 -5469 -5674 -5457
rect -5792 -5866 -5786 -5469
rect -5680 -5866 -5674 -5469
rect -5792 -5878 -5674 -5866
rect -5558 -5469 -5440 -5457
rect -5558 -5866 -5552 -5469
rect -5446 -5866 -5440 -5469
rect -5558 -5878 -5440 -5866
rect -5324 -5469 -5206 -5457
rect -5324 -5866 -5318 -5469
rect -5212 -5866 -5206 -5469
rect -5324 -5878 -5206 -5866
rect -5090 -5469 -4972 -5457
rect -5090 -5866 -5084 -5469
rect -4978 -5866 -4972 -5469
rect -5090 -5878 -4972 -5866
rect -4856 -5469 -4738 -5457
rect -4856 -5866 -4850 -5469
rect -4744 -5866 -4738 -5469
rect -4856 -5878 -4738 -5866
rect -4622 -5469 -4504 -5457
rect -4622 -5866 -4616 -5469
rect -4510 -5866 -4504 -5469
rect -4622 -5878 -4504 -5866
rect -4388 -5469 -4270 -5457
rect -4388 -5866 -4382 -5469
rect -4276 -5866 -4270 -5469
rect -4388 -5878 -4270 -5866
rect -4154 -5469 -4036 -5457
rect -4154 -5866 -4148 -5469
rect -4042 -5866 -4036 -5469
rect -4154 -5878 -4036 -5866
rect -3920 -5469 -3802 -5457
rect -3920 -5866 -3914 -5469
rect -3808 -5866 -3802 -5469
rect -3920 -5878 -3802 -5866
rect -3686 -5469 -3568 -5457
rect -3686 -5866 -3680 -5469
rect -3574 -5866 -3568 -5469
rect -3686 -5878 -3568 -5866
rect -3452 -5469 -3334 -5457
rect -3452 -5866 -3446 -5469
rect -3340 -5866 -3334 -5469
rect -3452 -5878 -3334 -5866
rect -3218 -5469 -3100 -5457
rect -3218 -5866 -3212 -5469
rect -3106 -5866 -3100 -5469
rect -3218 -5878 -3100 -5866
rect -2984 -5469 -2866 -5457
rect -2984 -5866 -2978 -5469
rect -2872 -5866 -2866 -5469
rect -2984 -5878 -2866 -5866
rect -2750 -5469 -2632 -5457
rect -2750 -5866 -2744 -5469
rect -2638 -5866 -2632 -5469
rect -2750 -5878 -2632 -5866
rect -2516 -5469 -2398 -5457
rect -2516 -5866 -2510 -5469
rect -2404 -5866 -2398 -5469
rect -2516 -5878 -2398 -5866
rect -2282 -5469 -2164 -5457
rect -2282 -5866 -2276 -5469
rect -2170 -5866 -2164 -5469
rect -2282 -5878 -2164 -5866
rect -2048 -5469 -1930 -5457
rect -2048 -5866 -2042 -5469
rect -1936 -5866 -1930 -5469
rect -2048 -5878 -1930 -5866
rect -1814 -5469 -1696 -5457
rect -1814 -5866 -1808 -5469
rect -1702 -5866 -1696 -5469
rect -1814 -5878 -1696 -5866
rect -1580 -5469 -1462 -5457
rect -1580 -5866 -1574 -5469
rect -1468 -5866 -1462 -5469
rect -1580 -5878 -1462 -5866
rect -1346 -5469 -1228 -5457
rect -1346 -5866 -1340 -5469
rect -1234 -5866 -1228 -5469
rect -1346 -5878 -1228 -5866
rect -1112 -5469 -994 -5457
rect -1112 -5866 -1106 -5469
rect -1000 -5866 -994 -5469
rect -1112 -5878 -994 -5866
rect -878 -5469 -760 -5457
rect -878 -5866 -872 -5469
rect -766 -5866 -760 -5469
rect -878 -5878 -760 -5866
rect -644 -5469 -526 -5457
rect -644 -5866 -638 -5469
rect -532 -5866 -526 -5469
rect -644 -5878 -526 -5866
rect -410 -5469 -292 -5457
rect -410 -5866 -404 -5469
rect -298 -5866 -292 -5469
rect -410 -5878 -292 -5866
rect -176 -5469 -58 -5457
rect -176 -5866 -170 -5469
rect -64 -5866 -58 -5469
rect -176 -5878 -58 -5866
rect 58 -5469 176 -5457
rect 58 -5866 64 -5469
rect 170 -5866 176 -5469
rect 58 -5878 176 -5866
rect 292 -5469 410 -5457
rect 292 -5866 298 -5469
rect 404 -5866 410 -5469
rect 292 -5878 410 -5866
rect 526 -5469 644 -5457
rect 526 -5866 532 -5469
rect 638 -5866 644 -5469
rect 526 -5878 644 -5866
rect 760 -5469 878 -5457
rect 760 -5866 766 -5469
rect 872 -5866 878 -5469
rect 760 -5878 878 -5866
rect 994 -5469 1112 -5457
rect 994 -5866 1000 -5469
rect 1106 -5866 1112 -5469
rect 994 -5878 1112 -5866
rect 1228 -5469 1346 -5457
rect 1228 -5866 1234 -5469
rect 1340 -5866 1346 -5469
rect 1228 -5878 1346 -5866
rect 1462 -5469 1580 -5457
rect 1462 -5866 1468 -5469
rect 1574 -5866 1580 -5469
rect 1462 -5878 1580 -5866
rect 1696 -5469 1814 -5457
rect 1696 -5866 1702 -5469
rect 1808 -5866 1814 -5469
rect 1696 -5878 1814 -5866
rect 1930 -5469 2048 -5457
rect 1930 -5866 1936 -5469
rect 2042 -5866 2048 -5469
rect 1930 -5878 2048 -5866
rect 2164 -5469 2282 -5457
rect 2164 -5866 2170 -5469
rect 2276 -5866 2282 -5469
rect 2164 -5878 2282 -5866
rect 2398 -5469 2516 -5457
rect 2398 -5866 2404 -5469
rect 2510 -5866 2516 -5469
rect 2398 -5878 2516 -5866
rect 2632 -5469 2750 -5457
rect 2632 -5866 2638 -5469
rect 2744 -5866 2750 -5469
rect 2632 -5878 2750 -5866
rect 2866 -5469 2984 -5457
rect 2866 -5866 2872 -5469
rect 2978 -5866 2984 -5469
rect 2866 -5878 2984 -5866
rect 3100 -5469 3218 -5457
rect 3100 -5866 3106 -5469
rect 3212 -5866 3218 -5469
rect 3100 -5878 3218 -5866
rect 3334 -5469 3452 -5457
rect 3334 -5866 3340 -5469
rect 3446 -5866 3452 -5469
rect 3334 -5878 3452 -5866
rect 3568 -5469 3686 -5457
rect 3568 -5866 3574 -5469
rect 3680 -5866 3686 -5469
rect 3568 -5878 3686 -5866
rect 3802 -5469 3920 -5457
rect 3802 -5866 3808 -5469
rect 3914 -5866 3920 -5469
rect 3802 -5878 3920 -5866
rect 4036 -5469 4154 -5457
rect 4036 -5866 4042 -5469
rect 4148 -5866 4154 -5469
rect 4036 -5878 4154 -5866
rect 4270 -5469 4388 -5457
rect 4270 -5866 4276 -5469
rect 4382 -5866 4388 -5469
rect 4270 -5878 4388 -5866
rect 4504 -5469 4622 -5457
rect 4504 -5866 4510 -5469
rect 4616 -5866 4622 -5469
rect 4504 -5878 4622 -5866
rect 4738 -5469 4856 -5457
rect 4738 -5866 4744 -5469
rect 4850 -5866 4856 -5469
rect 4738 -5878 4856 -5866
rect 4972 -5469 5090 -5457
rect 4972 -5866 4978 -5469
rect 5084 -5866 5090 -5469
rect 4972 -5878 5090 -5866
rect 5206 -5469 5324 -5457
rect 5206 -5866 5212 -5469
rect 5318 -5866 5324 -5469
rect 5206 -5878 5324 -5866
rect 5440 -5469 5558 -5457
rect 5440 -5866 5446 -5469
rect 5552 -5866 5558 -5469
rect 5440 -5878 5558 -5866
rect 5674 -5469 5792 -5457
rect 5674 -5866 5680 -5469
rect 5786 -5866 5792 -5469
rect 5674 -5878 5792 -5866
rect 5908 -5469 6026 -5457
rect 5908 -5866 5914 -5469
rect 6020 -5866 6026 -5469
rect 5908 -5878 6026 -5866
rect 6142 -5469 6260 -5457
rect 6142 -5866 6148 -5469
rect 6254 -5866 6260 -5469
rect 6142 -5878 6260 -5866
rect 6376 -5469 6494 -5457
rect 6376 -5866 6382 -5469
rect 6488 -5866 6494 -5469
rect 6376 -5878 6494 -5866
rect 6610 -5469 6728 -5457
rect 6610 -5866 6616 -5469
rect 6722 -5866 6728 -5469
rect 6610 -5878 6728 -5866
rect 6844 -5469 6962 -5457
rect 6844 -5866 6850 -5469
rect 6956 -5866 6962 -5469
rect 6844 -5878 6962 -5866
rect 7078 -5469 7196 -5457
rect 7078 -5866 7084 -5469
rect 7190 -5866 7196 -5469
rect 7078 -5878 7196 -5866
rect 7312 -5469 7430 -5457
rect 7312 -5866 7318 -5469
rect 7424 -5866 7430 -5469
rect 7312 -5878 7430 -5866
rect 7546 -5469 7664 -5457
rect 7546 -5866 7552 -5469
rect 7658 -5866 7664 -5469
rect 7546 -5878 7664 -5866
rect 7780 -5469 7898 -5457
rect 7780 -5866 7786 -5469
rect 7892 -5866 7898 -5469
rect 7780 -5878 7898 -5866
rect 8014 -5469 8132 -5457
rect 8014 -5866 8020 -5469
rect 8126 -5866 8132 -5469
rect 8014 -5878 8132 -5866
rect 8248 -5469 8366 -5457
rect 8248 -5866 8254 -5469
rect 8360 -5866 8366 -5469
rect 8248 -5878 8366 -5866
rect 8482 -5469 8600 -5457
rect 8482 -5866 8488 -5469
rect 8594 -5866 8600 -5469
rect 8482 -5878 8600 -5866
rect 8716 -5469 8834 -5457
rect 8716 -5866 8722 -5469
rect 8828 -5866 8834 -5469
rect 8716 -5878 8834 -5866
rect 8950 -5469 9068 -5457
rect 8950 -5866 8956 -5469
rect 9062 -5866 9068 -5469
rect 8950 -5878 9068 -5866
rect 9184 -5469 9302 -5457
rect 9184 -5866 9190 -5469
rect 9296 -5866 9302 -5469
rect 9184 -5878 9302 -5866
rect 9418 -5469 9536 -5457
rect 9418 -5866 9424 -5469
rect 9530 -5866 9536 -5469
rect 9418 -5878 9536 -5866
rect 9652 -5469 9770 -5457
rect 9652 -5866 9658 -5469
rect 9764 -5866 9770 -5469
rect 9652 -5878 9770 -5866
rect 9886 -5469 10004 -5457
rect 9886 -5866 9892 -5469
rect 9998 -5866 10004 -5469
rect 9886 -5878 10004 -5866
rect 10120 -5469 10238 -5457
rect 10120 -5866 10126 -5469
rect 10232 -5866 10238 -5469
rect 10120 -5878 10238 -5866
rect 10354 -5469 10472 -5457
rect 10354 -5866 10360 -5469
rect 10466 -5866 10472 -5469
rect 10354 -5878 10472 -5866
rect 10588 -5469 10706 -5457
rect 10588 -5866 10594 -5469
rect 10700 -5866 10706 -5469
rect 10588 -5878 10706 -5866
rect 10822 -5469 10940 -5457
rect 10822 -5866 10828 -5469
rect 10934 -5866 10940 -5469
rect 10822 -5878 10940 -5866
rect 11056 -5469 11174 -5457
rect 11056 -5866 11062 -5469
rect 11168 -5866 11174 -5469
rect 11056 -5878 11174 -5866
rect 11290 -5469 11408 -5457
rect 11290 -5866 11296 -5469
rect 11402 -5866 11408 -5469
rect 11290 -5878 11408 -5866
rect 11524 -5469 11642 -5457
rect 11524 -5866 11530 -5469
rect 11636 -5866 11642 -5469
rect 11524 -5878 11642 -5866
rect 11758 -5469 11876 -5457
rect 11758 -5866 11764 -5469
rect 11870 -5866 11876 -5469
rect 11758 -5878 11876 -5866
rect 11992 -5469 12110 -5457
rect 11992 -5866 11998 -5469
rect 12104 -5866 12110 -5469
rect 11992 -5878 12110 -5866
rect 12226 -5469 12344 -5457
rect 12226 -5866 12232 -5469
rect 12338 -5866 12344 -5469
rect 12226 -5878 12344 -5866
rect 12460 -5469 12578 -5457
rect 12460 -5866 12466 -5469
rect 12572 -5866 12578 -5469
rect 12460 -5878 12578 -5866
rect 12694 -5469 12812 -5457
rect 12694 -5866 12700 -5469
rect 12806 -5866 12812 -5469
rect 12694 -5878 12812 -5866
rect 12928 -5469 13046 -5457
rect 12928 -5866 12934 -5469
rect 13040 -5866 13046 -5469
rect 12928 -5878 13046 -5866
rect 13162 -5469 13280 -5457
rect 13162 -5866 13168 -5469
rect 13274 -5866 13280 -5469
rect 13162 -5878 13280 -5866
rect 13396 -5469 13514 -5457
rect 13396 -5866 13402 -5469
rect 13508 -5866 13514 -5469
rect 13396 -5878 13514 -5866
rect 13630 -5469 13748 -5457
rect 13630 -5866 13636 -5469
rect 13742 -5866 13748 -5469
rect 13630 -5878 13748 -5866
rect 13864 -5469 13982 -5457
rect 13864 -5866 13870 -5469
rect 13976 -5866 13982 -5469
rect 13864 -5878 13982 -5866
rect 14098 -5469 14216 -5457
rect 14098 -5866 14104 -5469
rect 14210 -5866 14216 -5469
rect 14098 -5878 14216 -5866
rect 14332 -5469 14450 -5457
rect 14332 -5866 14338 -5469
rect 14444 -5866 14450 -5469
rect 14332 -5878 14450 -5866
rect 14566 -5469 14684 -5457
rect 14566 -5866 14572 -5469
rect 14678 -5866 14684 -5469
rect 14566 -5878 14684 -5866
rect 14800 -5469 14918 -5457
rect 14800 -5866 14806 -5469
rect 14912 -5866 14918 -5469
rect 14800 -5878 14918 -5866
rect 15034 -5469 15152 -5457
rect 15034 -5866 15040 -5469
rect 15146 -5866 15152 -5469
rect 15034 -5878 15152 -5866
rect 15268 -5469 15386 -5457
rect 15268 -5866 15274 -5469
rect 15380 -5866 15386 -5469
rect 15268 -5878 15386 -5866
rect 15502 -5469 15620 -5457
rect 15502 -5866 15508 -5469
rect 15614 -5866 15620 -5469
rect 15502 -5878 15620 -5866
rect 15736 -5469 15854 -5457
rect 15736 -5866 15742 -5469
rect 15848 -5866 15854 -5469
rect 15736 -5878 15854 -5866
rect 15970 -5469 16088 -5457
rect 15970 -5866 15976 -5469
rect 16082 -5866 16088 -5469
rect 15970 -5878 16088 -5866
rect 16204 -5469 16322 -5457
rect 16204 -5866 16210 -5469
rect 16316 -5866 16322 -5469
rect 16204 -5878 16322 -5866
rect 16438 -5469 16556 -5457
rect 16438 -5866 16444 -5469
rect 16550 -5866 16556 -5469
rect 16438 -5878 16556 -5866
rect 16672 -5469 16790 -5457
rect 16672 -5866 16678 -5469
rect 16784 -5866 16790 -5469
rect 16672 -5878 16790 -5866
rect 16906 -5469 17024 -5457
rect 16906 -5866 16912 -5469
rect 17018 -5866 17024 -5469
rect 16906 -5878 17024 -5866
rect 17140 -5469 17258 -5457
rect 17140 -5866 17146 -5469
rect 17252 -5866 17258 -5469
rect 17140 -5878 17258 -5866
rect 17374 -5469 17492 -5457
rect 17374 -5866 17380 -5469
rect 17486 -5866 17492 -5469
rect 17374 -5878 17492 -5866
rect 17608 -5469 17726 -5457
rect 17608 -5866 17614 -5469
rect 17720 -5866 17726 -5469
rect 17608 -5878 17726 -5866
rect 17842 -5469 17960 -5457
rect 17842 -5866 17848 -5469
rect 17954 -5866 17960 -5469
rect 17842 -5878 17960 -5866
rect 18076 -5469 18194 -5457
rect 18076 -5866 18082 -5469
rect 18188 -5866 18194 -5469
rect 18076 -5878 18194 -5866
rect 18310 -5469 18428 -5457
rect 18310 -5866 18316 -5469
rect 18422 -5866 18428 -5469
rect 18310 -5878 18428 -5866
rect 18544 -5469 18662 -5457
rect 18544 -5866 18550 -5469
rect 18656 -5866 18662 -5469
rect 18544 -5878 18662 -5866
rect 18778 -5469 18896 -5457
rect 18778 -5866 18784 -5469
rect 18890 -5866 18896 -5469
rect 18778 -5878 18896 -5866
rect 19012 -5469 19130 -5457
rect 19012 -5866 19018 -5469
rect 19124 -5866 19130 -5469
rect 19012 -5878 19130 -5866
rect 19246 -5469 19364 -5457
rect 19246 -5866 19252 -5469
rect 19358 -5866 19364 -5469
rect 19246 -5878 19364 -5866
rect 19480 -5469 19598 -5457
rect 19480 -5866 19486 -5469
rect 19592 -5866 19598 -5469
rect 19480 -5878 19598 -5866
rect 19714 -5469 19832 -5457
rect 19714 -5866 19720 -5469
rect 19826 -5866 19832 -5469
rect 19714 -5878 19832 -5866
rect 19948 -5469 20066 -5457
rect 19948 -5866 19954 -5469
rect 20060 -5866 20066 -5469
rect 19948 -5878 20066 -5866
rect 20182 -5469 20300 -5457
rect 20182 -5866 20188 -5469
rect 20294 -5866 20300 -5469
rect 20182 -5878 20300 -5866
rect 20416 -5469 20534 -5457
rect 20416 -5866 20422 -5469
rect 20528 -5866 20534 -5469
rect 20416 -5878 20534 -5866
rect 20650 -5469 20768 -5457
rect 20650 -5866 20656 -5469
rect 20762 -5866 20768 -5469
rect 20650 -5878 20768 -5866
rect 20884 -5469 21002 -5457
rect 20884 -5866 20890 -5469
rect 20996 -5866 21002 -5469
rect 20884 -5878 21002 -5866
rect 21118 -5469 21236 -5457
rect 21118 -5866 21124 -5469
rect 21230 -5866 21236 -5469
rect 21118 -5878 21236 -5866
rect 21352 -5469 21470 -5457
rect 21352 -5866 21358 -5469
rect 21464 -5866 21470 -5469
rect 21352 -5878 21470 -5866
rect 21586 -5469 21704 -5457
rect 21586 -5866 21592 -5469
rect 21698 -5866 21704 -5469
rect 21586 -5878 21704 -5866
rect 21820 -5469 21938 -5457
rect 21820 -5866 21826 -5469
rect 21932 -5866 21938 -5469
rect 21820 -5878 21938 -5866
rect 22054 -5469 22172 -5457
rect 22054 -5866 22060 -5469
rect 22166 -5866 22172 -5469
rect 22054 -5878 22172 -5866
rect 22288 -5469 22406 -5457
rect 22288 -5866 22294 -5469
rect 22400 -5866 22406 -5469
rect 22288 -5878 22406 -5866
rect 22522 -5469 22640 -5457
rect 22522 -5866 22528 -5469
rect 22634 -5866 22640 -5469
rect 22522 -5878 22640 -5866
rect 22756 -5469 22874 -5457
rect 22756 -5866 22762 -5469
rect 22868 -5866 22874 -5469
rect 22756 -5878 22874 -5866
rect 22990 -5469 23108 -5457
rect 22990 -5866 22996 -5469
rect 23102 -5866 23108 -5469
rect 22990 -5878 23108 -5866
rect 23224 -5469 23342 -5457
rect 23224 -5866 23230 -5469
rect 23336 -5866 23342 -5469
rect 23224 -5878 23342 -5866
rect 23458 -5469 23576 -5457
rect 23458 -5866 23464 -5469
rect 23570 -5866 23576 -5469
rect 23458 -5878 23576 -5866
rect 23692 -5469 23810 -5457
rect 23692 -5866 23698 -5469
rect 23804 -5866 23810 -5469
rect 23692 -5878 23810 -5866
rect 23926 -5469 24044 -5457
rect 23926 -5866 23932 -5469
rect 24038 -5866 24044 -5469
rect 23926 -5878 24044 -5866
rect 24160 -5469 24278 -5457
rect 24160 -5866 24166 -5469
rect 24272 -5866 24278 -5469
rect 24160 -5878 24278 -5866
rect 24394 -5469 24512 -5457
rect 24394 -5866 24400 -5469
rect 24506 -5866 24512 -5469
rect 24394 -5878 24512 -5866
rect 24628 -5469 24746 -5457
rect 24628 -5866 24634 -5469
rect 24740 -5866 24746 -5469
rect 24628 -5878 24746 -5866
rect 24862 -5469 24980 -5457
rect 24862 -5866 24868 -5469
rect 24974 -5866 24980 -5469
rect 24862 -5878 24980 -5866
rect 25096 -5469 25214 -5457
rect 25096 -5866 25102 -5469
rect 25208 -5866 25214 -5469
rect 25096 -5878 25214 -5866
rect 25330 -5469 25448 -5457
rect 25330 -5866 25336 -5469
rect 25442 -5866 25448 -5469
rect 25330 -5878 25448 -5866
rect 25564 -5469 25682 -5457
rect 25564 -5866 25570 -5469
rect 25676 -5866 25682 -5469
rect 25564 -5878 25682 -5866
rect 25798 -5469 25916 -5457
rect 25798 -5866 25804 -5469
rect 25910 -5866 25916 -5469
rect 25798 -5878 25916 -5866
rect 26032 -5469 26150 -5457
rect 26032 -5866 26038 -5469
rect 26144 -5866 26150 -5469
rect 26032 -5878 26150 -5866
rect 26266 -5469 26384 -5457
rect 26266 -5866 26272 -5469
rect 26378 -5866 26384 -5469
rect 26266 -5878 26384 -5866
rect 26500 -5469 26618 -5457
rect 26500 -5866 26506 -5469
rect 26612 -5866 26618 -5469
rect 26500 -5878 26618 -5866
rect 26734 -5469 26852 -5457
rect 26734 -5866 26740 -5469
rect 26846 -5866 26852 -5469
rect 26734 -5878 26852 -5866
rect 26968 -5469 27086 -5457
rect 26968 -5866 26974 -5469
rect 27080 -5866 27086 -5469
rect 26968 -5878 27086 -5866
rect 27202 -5469 27320 -5457
rect 27202 -5866 27208 -5469
rect 27314 -5866 27320 -5469
rect 27202 -5878 27320 -5866
rect 27436 -5469 27554 -5457
rect 27436 -5866 27442 -5469
rect 27548 -5866 27554 -5469
rect 27436 -5878 27554 -5866
rect 27670 -5469 27788 -5457
rect 27670 -5866 27676 -5469
rect 27782 -5866 27788 -5469
rect 27670 -5878 27788 -5866
rect 27904 -5469 28022 -5457
rect 27904 -5866 27910 -5469
rect 28016 -5866 28022 -5469
rect 27904 -5878 28022 -5866
rect 28138 -5469 28256 -5457
rect 28138 -5866 28144 -5469
rect 28250 -5866 28256 -5469
rect 28138 -5878 28256 -5866
rect 28372 -5469 28490 -5457
rect 28372 -5866 28378 -5469
rect 28484 -5866 28490 -5469
rect 28372 -5878 28490 -5866
rect 28606 -5469 28724 -5457
rect 28606 -5866 28612 -5469
rect 28718 -5866 28724 -5469
rect 28606 -5878 28724 -5866
rect 28840 -5469 28958 -5457
rect 28840 -5866 28846 -5469
rect 28952 -5866 28958 -5469
rect 28840 -5878 28958 -5866
rect 29074 -5469 29192 -5457
rect 29074 -5866 29080 -5469
rect 29186 -5866 29192 -5469
rect 29074 -5878 29192 -5866
rect 29308 -5469 29426 -5457
rect 29308 -5866 29314 -5469
rect 29420 -5866 29426 -5469
rect 29308 -5878 29426 -5866
rect 29542 -5469 29660 -5457
rect 29542 -5866 29548 -5469
rect 29654 -5866 29660 -5469
rect 29542 -5878 29660 -5866
rect 29776 -5469 29894 -5457
rect 29776 -5866 29782 -5469
rect 29888 -5866 29894 -5469
rect 29776 -5878 29894 -5866
<< properties >>
string FIXED_BBOX -30017 -5997 30017 5997
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 25.0 m 2 nx 256 wmin 0.690 lmin 0.50 class resistor rho 319.8 val 12.151k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
