magic
tech sky130A
magscale 1 2
timestamp 1730743893
<< error_p >>
rect 10828 30694 10886 30700
rect 10828 30660 10840 30694
rect 10828 30654 10886 30660
rect 11438 30648 11496 30654
rect 11438 30614 11450 30648
rect 11438 30608 11496 30614
rect 19690 29890 19748 29896
rect 19690 29856 19702 29890
rect 19690 29850 19748 29856
rect 10828 29084 10886 29090
rect 10828 29050 10840 29084
rect 10828 29044 10886 29050
rect 11438 29038 11496 29044
rect 11438 29004 11450 29038
rect 11438 28998 11496 29004
rect 19690 28280 19748 28286
rect 19690 28246 19702 28280
rect 19690 28240 19748 28246
rect 19742 27682 19800 27688
rect 19742 27648 19754 27682
rect 19742 27642 19800 27648
rect 15594 27268 18158 27270
rect 19742 26072 19800 26078
rect 19742 26038 19754 26072
rect 19742 26032 19800 26038
rect 19630 21168 19688 21174
rect 19630 21134 19642 21168
rect 19630 21128 19688 21134
rect 4428 15098 4478 18216
rect 7554 15148 10540 15162
rect 2118 13364 2176 13370
rect 2118 13330 2130 13364
rect 2118 13324 2176 13330
rect 2118 11754 2176 11760
rect 2118 11720 2130 11754
rect 2118 11714 2176 11720
rect 2184 11150 2242 11156
rect 2184 11116 2196 11150
rect 2184 11110 2242 11116
rect 2184 9540 2242 9546
rect 2184 9506 2196 9540
rect 2184 9500 2242 9506
rect 4468 5834 4518 8272
<< error_s >>
rect 19630 19558 19688 19564
rect 4428 19476 4478 19536
rect 19630 19524 19642 19558
rect 19630 19518 19688 19524
rect 19682 18960 19740 18966
rect 19682 18926 19694 18960
rect 19682 18920 19740 18926
rect 19682 17350 19740 17356
rect 19682 17316 19694 17350
rect 19682 17310 19740 17316
rect 2158 490 2216 496
rect 2158 456 2170 490
rect 2158 450 2216 456
rect 2224 -114 2282 -108
rect 2224 -148 2236 -114
rect 2224 -154 2282 -148
rect 2224 -1724 2282 -1718
rect 2224 -1758 2236 -1724
rect 2224 -1764 2282 -1758
<< error_ps >>
rect 4428 18216 4478 19476
rect 4468 3834 4518 5834
rect 7594 3884 10580 3898
rect 2158 2100 2216 2106
rect 2158 2066 2170 2100
rect 2158 2060 2216 2066
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
rect 0 -6400 200 -6200
rect 0 -6800 200 -6600
use Parallel_10B_Block2  x1
timestamp 1730743893
transform 1 0 0 0 1 -6800
box 0 -6800 37772 26360
use Input_Stage_v1  x2
timestamp 1730739923
transform 1 0 1472 0 1 23250
box 0 -19414 36640 8756
use vbias_gen_pga  x3
timestamp 1729620069
transform 1 0 1355 0 1 25173
box -65 -865 591 651
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {V\[9\]}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 {V\[8\]}
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 {V\[7\]}
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 {V\[6\]}
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 {V\[5\]}
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 {V\[4\]}
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 {V\[3\]}
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 {V\[2\]}
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 {V\[1\]}
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 {V\[0\]}
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 VCM
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 IBIAS
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 AVDD
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 VIN
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 DVDD
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 256 0 0 0 VOUT
port 15 nsew
flabel metal1 0 -6400 200 -6200 0 FreeSans 256 0 0 0 AVSS
port 16 nsew
flabel metal1 0 -6800 200 -6600 0 FreeSans 256 0 0 0 DVSS
port 17 nsew
<< end >>
