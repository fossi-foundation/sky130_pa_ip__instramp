magic
tech sky130A
magscale 1 2
timestamp 1730737834
<< pwell >>
rect -5875 -2978 5875 2978
<< mvnmos >>
rect -5647 1720 -5447 2720
rect -5389 1720 -5189 2720
rect -5131 1720 -4931 2720
rect -4873 1720 -4673 2720
rect -4615 1720 -4415 2720
rect -4357 1720 -4157 2720
rect -4099 1720 -3899 2720
rect -3841 1720 -3641 2720
rect -3583 1720 -3383 2720
rect -3325 1720 -3125 2720
rect -3067 1720 -2867 2720
rect -2809 1720 -2609 2720
rect -2551 1720 -2351 2720
rect -2293 1720 -2093 2720
rect -2035 1720 -1835 2720
rect -1777 1720 -1577 2720
rect -1519 1720 -1319 2720
rect -1261 1720 -1061 2720
rect -1003 1720 -803 2720
rect -745 1720 -545 2720
rect -487 1720 -287 2720
rect -229 1720 -29 2720
rect 29 1720 229 2720
rect 287 1720 487 2720
rect 545 1720 745 2720
rect 803 1720 1003 2720
rect 1061 1720 1261 2720
rect 1319 1720 1519 2720
rect 1577 1720 1777 2720
rect 1835 1720 2035 2720
rect 2093 1720 2293 2720
rect 2351 1720 2551 2720
rect 2609 1720 2809 2720
rect 2867 1720 3067 2720
rect 3125 1720 3325 2720
rect 3383 1720 3583 2720
rect 3641 1720 3841 2720
rect 3899 1720 4099 2720
rect 4157 1720 4357 2720
rect 4415 1720 4615 2720
rect 4673 1720 4873 2720
rect 4931 1720 5131 2720
rect 5189 1720 5389 2720
rect 5447 1720 5647 2720
rect -5647 610 -5447 1610
rect -5389 610 -5189 1610
rect -5131 610 -4931 1610
rect -4873 610 -4673 1610
rect -4615 610 -4415 1610
rect -4357 610 -4157 1610
rect -4099 610 -3899 1610
rect -3841 610 -3641 1610
rect -3583 610 -3383 1610
rect -3325 610 -3125 1610
rect -3067 610 -2867 1610
rect -2809 610 -2609 1610
rect -2551 610 -2351 1610
rect -2293 610 -2093 1610
rect -2035 610 -1835 1610
rect -1777 610 -1577 1610
rect -1519 610 -1319 1610
rect -1261 610 -1061 1610
rect -1003 610 -803 1610
rect -745 610 -545 1610
rect -487 610 -287 1610
rect -229 610 -29 1610
rect 29 610 229 1610
rect 287 610 487 1610
rect 545 610 745 1610
rect 803 610 1003 1610
rect 1061 610 1261 1610
rect 1319 610 1519 1610
rect 1577 610 1777 1610
rect 1835 610 2035 1610
rect 2093 610 2293 1610
rect 2351 610 2551 1610
rect 2609 610 2809 1610
rect 2867 610 3067 1610
rect 3125 610 3325 1610
rect 3383 610 3583 1610
rect 3641 610 3841 1610
rect 3899 610 4099 1610
rect 4157 610 4357 1610
rect 4415 610 4615 1610
rect 4673 610 4873 1610
rect 4931 610 5131 1610
rect 5189 610 5389 1610
rect 5447 610 5647 1610
rect -5647 -500 -5447 500
rect -5389 -500 -5189 500
rect -5131 -500 -4931 500
rect -4873 -500 -4673 500
rect -4615 -500 -4415 500
rect -4357 -500 -4157 500
rect -4099 -500 -3899 500
rect -3841 -500 -3641 500
rect -3583 -500 -3383 500
rect -3325 -500 -3125 500
rect -3067 -500 -2867 500
rect -2809 -500 -2609 500
rect -2551 -500 -2351 500
rect -2293 -500 -2093 500
rect -2035 -500 -1835 500
rect -1777 -500 -1577 500
rect -1519 -500 -1319 500
rect -1261 -500 -1061 500
rect -1003 -500 -803 500
rect -745 -500 -545 500
rect -487 -500 -287 500
rect -229 -500 -29 500
rect 29 -500 229 500
rect 287 -500 487 500
rect 545 -500 745 500
rect 803 -500 1003 500
rect 1061 -500 1261 500
rect 1319 -500 1519 500
rect 1577 -500 1777 500
rect 1835 -500 2035 500
rect 2093 -500 2293 500
rect 2351 -500 2551 500
rect 2609 -500 2809 500
rect 2867 -500 3067 500
rect 3125 -500 3325 500
rect 3383 -500 3583 500
rect 3641 -500 3841 500
rect 3899 -500 4099 500
rect 4157 -500 4357 500
rect 4415 -500 4615 500
rect 4673 -500 4873 500
rect 4931 -500 5131 500
rect 5189 -500 5389 500
rect 5447 -500 5647 500
rect -5647 -1610 -5447 -610
rect -5389 -1610 -5189 -610
rect -5131 -1610 -4931 -610
rect -4873 -1610 -4673 -610
rect -4615 -1610 -4415 -610
rect -4357 -1610 -4157 -610
rect -4099 -1610 -3899 -610
rect -3841 -1610 -3641 -610
rect -3583 -1610 -3383 -610
rect -3325 -1610 -3125 -610
rect -3067 -1610 -2867 -610
rect -2809 -1610 -2609 -610
rect -2551 -1610 -2351 -610
rect -2293 -1610 -2093 -610
rect -2035 -1610 -1835 -610
rect -1777 -1610 -1577 -610
rect -1519 -1610 -1319 -610
rect -1261 -1610 -1061 -610
rect -1003 -1610 -803 -610
rect -745 -1610 -545 -610
rect -487 -1610 -287 -610
rect -229 -1610 -29 -610
rect 29 -1610 229 -610
rect 287 -1610 487 -610
rect 545 -1610 745 -610
rect 803 -1610 1003 -610
rect 1061 -1610 1261 -610
rect 1319 -1610 1519 -610
rect 1577 -1610 1777 -610
rect 1835 -1610 2035 -610
rect 2093 -1610 2293 -610
rect 2351 -1610 2551 -610
rect 2609 -1610 2809 -610
rect 2867 -1610 3067 -610
rect 3125 -1610 3325 -610
rect 3383 -1610 3583 -610
rect 3641 -1610 3841 -610
rect 3899 -1610 4099 -610
rect 4157 -1610 4357 -610
rect 4415 -1610 4615 -610
rect 4673 -1610 4873 -610
rect 4931 -1610 5131 -610
rect 5189 -1610 5389 -610
rect 5447 -1610 5647 -610
rect -5647 -2720 -5447 -1720
rect -5389 -2720 -5189 -1720
rect -5131 -2720 -4931 -1720
rect -4873 -2720 -4673 -1720
rect -4615 -2720 -4415 -1720
rect -4357 -2720 -4157 -1720
rect -4099 -2720 -3899 -1720
rect -3841 -2720 -3641 -1720
rect -3583 -2720 -3383 -1720
rect -3325 -2720 -3125 -1720
rect -3067 -2720 -2867 -1720
rect -2809 -2720 -2609 -1720
rect -2551 -2720 -2351 -1720
rect -2293 -2720 -2093 -1720
rect -2035 -2720 -1835 -1720
rect -1777 -2720 -1577 -1720
rect -1519 -2720 -1319 -1720
rect -1261 -2720 -1061 -1720
rect -1003 -2720 -803 -1720
rect -745 -2720 -545 -1720
rect -487 -2720 -287 -1720
rect -229 -2720 -29 -1720
rect 29 -2720 229 -1720
rect 287 -2720 487 -1720
rect 545 -2720 745 -1720
rect 803 -2720 1003 -1720
rect 1061 -2720 1261 -1720
rect 1319 -2720 1519 -1720
rect 1577 -2720 1777 -1720
rect 1835 -2720 2035 -1720
rect 2093 -2720 2293 -1720
rect 2351 -2720 2551 -1720
rect 2609 -2720 2809 -1720
rect 2867 -2720 3067 -1720
rect 3125 -2720 3325 -1720
rect 3383 -2720 3583 -1720
rect 3641 -2720 3841 -1720
rect 3899 -2720 4099 -1720
rect 4157 -2720 4357 -1720
rect 4415 -2720 4615 -1720
rect 4673 -2720 4873 -1720
rect 4931 -2720 5131 -1720
rect 5189 -2720 5389 -1720
rect 5447 -2720 5647 -1720
<< mvndiff >>
rect -5705 2708 -5647 2720
rect -5705 1732 -5693 2708
rect -5659 1732 -5647 2708
rect -5705 1720 -5647 1732
rect -5447 2708 -5389 2720
rect -5447 1732 -5435 2708
rect -5401 1732 -5389 2708
rect -5447 1720 -5389 1732
rect -5189 2708 -5131 2720
rect -5189 1732 -5177 2708
rect -5143 1732 -5131 2708
rect -5189 1720 -5131 1732
rect -4931 2708 -4873 2720
rect -4931 1732 -4919 2708
rect -4885 1732 -4873 2708
rect -4931 1720 -4873 1732
rect -4673 2708 -4615 2720
rect -4673 1732 -4661 2708
rect -4627 1732 -4615 2708
rect -4673 1720 -4615 1732
rect -4415 2708 -4357 2720
rect -4415 1732 -4403 2708
rect -4369 1732 -4357 2708
rect -4415 1720 -4357 1732
rect -4157 2708 -4099 2720
rect -4157 1732 -4145 2708
rect -4111 1732 -4099 2708
rect -4157 1720 -4099 1732
rect -3899 2708 -3841 2720
rect -3899 1732 -3887 2708
rect -3853 1732 -3841 2708
rect -3899 1720 -3841 1732
rect -3641 2708 -3583 2720
rect -3641 1732 -3629 2708
rect -3595 1732 -3583 2708
rect -3641 1720 -3583 1732
rect -3383 2708 -3325 2720
rect -3383 1732 -3371 2708
rect -3337 1732 -3325 2708
rect -3383 1720 -3325 1732
rect -3125 2708 -3067 2720
rect -3125 1732 -3113 2708
rect -3079 1732 -3067 2708
rect -3125 1720 -3067 1732
rect -2867 2708 -2809 2720
rect -2867 1732 -2855 2708
rect -2821 1732 -2809 2708
rect -2867 1720 -2809 1732
rect -2609 2708 -2551 2720
rect -2609 1732 -2597 2708
rect -2563 1732 -2551 2708
rect -2609 1720 -2551 1732
rect -2351 2708 -2293 2720
rect -2351 1732 -2339 2708
rect -2305 1732 -2293 2708
rect -2351 1720 -2293 1732
rect -2093 2708 -2035 2720
rect -2093 1732 -2081 2708
rect -2047 1732 -2035 2708
rect -2093 1720 -2035 1732
rect -1835 2708 -1777 2720
rect -1835 1732 -1823 2708
rect -1789 1732 -1777 2708
rect -1835 1720 -1777 1732
rect -1577 2708 -1519 2720
rect -1577 1732 -1565 2708
rect -1531 1732 -1519 2708
rect -1577 1720 -1519 1732
rect -1319 2708 -1261 2720
rect -1319 1732 -1307 2708
rect -1273 1732 -1261 2708
rect -1319 1720 -1261 1732
rect -1061 2708 -1003 2720
rect -1061 1732 -1049 2708
rect -1015 1732 -1003 2708
rect -1061 1720 -1003 1732
rect -803 2708 -745 2720
rect -803 1732 -791 2708
rect -757 1732 -745 2708
rect -803 1720 -745 1732
rect -545 2708 -487 2720
rect -545 1732 -533 2708
rect -499 1732 -487 2708
rect -545 1720 -487 1732
rect -287 2708 -229 2720
rect -287 1732 -275 2708
rect -241 1732 -229 2708
rect -287 1720 -229 1732
rect -29 2708 29 2720
rect -29 1732 -17 2708
rect 17 1732 29 2708
rect -29 1720 29 1732
rect 229 2708 287 2720
rect 229 1732 241 2708
rect 275 1732 287 2708
rect 229 1720 287 1732
rect 487 2708 545 2720
rect 487 1732 499 2708
rect 533 1732 545 2708
rect 487 1720 545 1732
rect 745 2708 803 2720
rect 745 1732 757 2708
rect 791 1732 803 2708
rect 745 1720 803 1732
rect 1003 2708 1061 2720
rect 1003 1732 1015 2708
rect 1049 1732 1061 2708
rect 1003 1720 1061 1732
rect 1261 2708 1319 2720
rect 1261 1732 1273 2708
rect 1307 1732 1319 2708
rect 1261 1720 1319 1732
rect 1519 2708 1577 2720
rect 1519 1732 1531 2708
rect 1565 1732 1577 2708
rect 1519 1720 1577 1732
rect 1777 2708 1835 2720
rect 1777 1732 1789 2708
rect 1823 1732 1835 2708
rect 1777 1720 1835 1732
rect 2035 2708 2093 2720
rect 2035 1732 2047 2708
rect 2081 1732 2093 2708
rect 2035 1720 2093 1732
rect 2293 2708 2351 2720
rect 2293 1732 2305 2708
rect 2339 1732 2351 2708
rect 2293 1720 2351 1732
rect 2551 2708 2609 2720
rect 2551 1732 2563 2708
rect 2597 1732 2609 2708
rect 2551 1720 2609 1732
rect 2809 2708 2867 2720
rect 2809 1732 2821 2708
rect 2855 1732 2867 2708
rect 2809 1720 2867 1732
rect 3067 2708 3125 2720
rect 3067 1732 3079 2708
rect 3113 1732 3125 2708
rect 3067 1720 3125 1732
rect 3325 2708 3383 2720
rect 3325 1732 3337 2708
rect 3371 1732 3383 2708
rect 3325 1720 3383 1732
rect 3583 2708 3641 2720
rect 3583 1732 3595 2708
rect 3629 1732 3641 2708
rect 3583 1720 3641 1732
rect 3841 2708 3899 2720
rect 3841 1732 3853 2708
rect 3887 1732 3899 2708
rect 3841 1720 3899 1732
rect 4099 2708 4157 2720
rect 4099 1732 4111 2708
rect 4145 1732 4157 2708
rect 4099 1720 4157 1732
rect 4357 2708 4415 2720
rect 4357 1732 4369 2708
rect 4403 1732 4415 2708
rect 4357 1720 4415 1732
rect 4615 2708 4673 2720
rect 4615 1732 4627 2708
rect 4661 1732 4673 2708
rect 4615 1720 4673 1732
rect 4873 2708 4931 2720
rect 4873 1732 4885 2708
rect 4919 1732 4931 2708
rect 4873 1720 4931 1732
rect 5131 2708 5189 2720
rect 5131 1732 5143 2708
rect 5177 1732 5189 2708
rect 5131 1720 5189 1732
rect 5389 2708 5447 2720
rect 5389 1732 5401 2708
rect 5435 1732 5447 2708
rect 5389 1720 5447 1732
rect 5647 2708 5705 2720
rect 5647 1732 5659 2708
rect 5693 1732 5705 2708
rect 5647 1720 5705 1732
rect -5705 1598 -5647 1610
rect -5705 622 -5693 1598
rect -5659 622 -5647 1598
rect -5705 610 -5647 622
rect -5447 1598 -5389 1610
rect -5447 622 -5435 1598
rect -5401 622 -5389 1598
rect -5447 610 -5389 622
rect -5189 1598 -5131 1610
rect -5189 622 -5177 1598
rect -5143 622 -5131 1598
rect -5189 610 -5131 622
rect -4931 1598 -4873 1610
rect -4931 622 -4919 1598
rect -4885 622 -4873 1598
rect -4931 610 -4873 622
rect -4673 1598 -4615 1610
rect -4673 622 -4661 1598
rect -4627 622 -4615 1598
rect -4673 610 -4615 622
rect -4415 1598 -4357 1610
rect -4415 622 -4403 1598
rect -4369 622 -4357 1598
rect -4415 610 -4357 622
rect -4157 1598 -4099 1610
rect -4157 622 -4145 1598
rect -4111 622 -4099 1598
rect -4157 610 -4099 622
rect -3899 1598 -3841 1610
rect -3899 622 -3887 1598
rect -3853 622 -3841 1598
rect -3899 610 -3841 622
rect -3641 1598 -3583 1610
rect -3641 622 -3629 1598
rect -3595 622 -3583 1598
rect -3641 610 -3583 622
rect -3383 1598 -3325 1610
rect -3383 622 -3371 1598
rect -3337 622 -3325 1598
rect -3383 610 -3325 622
rect -3125 1598 -3067 1610
rect -3125 622 -3113 1598
rect -3079 622 -3067 1598
rect -3125 610 -3067 622
rect -2867 1598 -2809 1610
rect -2867 622 -2855 1598
rect -2821 622 -2809 1598
rect -2867 610 -2809 622
rect -2609 1598 -2551 1610
rect -2609 622 -2597 1598
rect -2563 622 -2551 1598
rect -2609 610 -2551 622
rect -2351 1598 -2293 1610
rect -2351 622 -2339 1598
rect -2305 622 -2293 1598
rect -2351 610 -2293 622
rect -2093 1598 -2035 1610
rect -2093 622 -2081 1598
rect -2047 622 -2035 1598
rect -2093 610 -2035 622
rect -1835 1598 -1777 1610
rect -1835 622 -1823 1598
rect -1789 622 -1777 1598
rect -1835 610 -1777 622
rect -1577 1598 -1519 1610
rect -1577 622 -1565 1598
rect -1531 622 -1519 1598
rect -1577 610 -1519 622
rect -1319 1598 -1261 1610
rect -1319 622 -1307 1598
rect -1273 622 -1261 1598
rect -1319 610 -1261 622
rect -1061 1598 -1003 1610
rect -1061 622 -1049 1598
rect -1015 622 -1003 1598
rect -1061 610 -1003 622
rect -803 1598 -745 1610
rect -803 622 -791 1598
rect -757 622 -745 1598
rect -803 610 -745 622
rect -545 1598 -487 1610
rect -545 622 -533 1598
rect -499 622 -487 1598
rect -545 610 -487 622
rect -287 1598 -229 1610
rect -287 622 -275 1598
rect -241 622 -229 1598
rect -287 610 -229 622
rect -29 1598 29 1610
rect -29 622 -17 1598
rect 17 622 29 1598
rect -29 610 29 622
rect 229 1598 287 1610
rect 229 622 241 1598
rect 275 622 287 1598
rect 229 610 287 622
rect 487 1598 545 1610
rect 487 622 499 1598
rect 533 622 545 1598
rect 487 610 545 622
rect 745 1598 803 1610
rect 745 622 757 1598
rect 791 622 803 1598
rect 745 610 803 622
rect 1003 1598 1061 1610
rect 1003 622 1015 1598
rect 1049 622 1061 1598
rect 1003 610 1061 622
rect 1261 1598 1319 1610
rect 1261 622 1273 1598
rect 1307 622 1319 1598
rect 1261 610 1319 622
rect 1519 1598 1577 1610
rect 1519 622 1531 1598
rect 1565 622 1577 1598
rect 1519 610 1577 622
rect 1777 1598 1835 1610
rect 1777 622 1789 1598
rect 1823 622 1835 1598
rect 1777 610 1835 622
rect 2035 1598 2093 1610
rect 2035 622 2047 1598
rect 2081 622 2093 1598
rect 2035 610 2093 622
rect 2293 1598 2351 1610
rect 2293 622 2305 1598
rect 2339 622 2351 1598
rect 2293 610 2351 622
rect 2551 1598 2609 1610
rect 2551 622 2563 1598
rect 2597 622 2609 1598
rect 2551 610 2609 622
rect 2809 1598 2867 1610
rect 2809 622 2821 1598
rect 2855 622 2867 1598
rect 2809 610 2867 622
rect 3067 1598 3125 1610
rect 3067 622 3079 1598
rect 3113 622 3125 1598
rect 3067 610 3125 622
rect 3325 1598 3383 1610
rect 3325 622 3337 1598
rect 3371 622 3383 1598
rect 3325 610 3383 622
rect 3583 1598 3641 1610
rect 3583 622 3595 1598
rect 3629 622 3641 1598
rect 3583 610 3641 622
rect 3841 1598 3899 1610
rect 3841 622 3853 1598
rect 3887 622 3899 1598
rect 3841 610 3899 622
rect 4099 1598 4157 1610
rect 4099 622 4111 1598
rect 4145 622 4157 1598
rect 4099 610 4157 622
rect 4357 1598 4415 1610
rect 4357 622 4369 1598
rect 4403 622 4415 1598
rect 4357 610 4415 622
rect 4615 1598 4673 1610
rect 4615 622 4627 1598
rect 4661 622 4673 1598
rect 4615 610 4673 622
rect 4873 1598 4931 1610
rect 4873 622 4885 1598
rect 4919 622 4931 1598
rect 4873 610 4931 622
rect 5131 1598 5189 1610
rect 5131 622 5143 1598
rect 5177 622 5189 1598
rect 5131 610 5189 622
rect 5389 1598 5447 1610
rect 5389 622 5401 1598
rect 5435 622 5447 1598
rect 5389 610 5447 622
rect 5647 1598 5705 1610
rect 5647 622 5659 1598
rect 5693 622 5705 1598
rect 5647 610 5705 622
rect -5705 488 -5647 500
rect -5705 -488 -5693 488
rect -5659 -488 -5647 488
rect -5705 -500 -5647 -488
rect -5447 488 -5389 500
rect -5447 -488 -5435 488
rect -5401 -488 -5389 488
rect -5447 -500 -5389 -488
rect -5189 488 -5131 500
rect -5189 -488 -5177 488
rect -5143 -488 -5131 488
rect -5189 -500 -5131 -488
rect -4931 488 -4873 500
rect -4931 -488 -4919 488
rect -4885 -488 -4873 488
rect -4931 -500 -4873 -488
rect -4673 488 -4615 500
rect -4673 -488 -4661 488
rect -4627 -488 -4615 488
rect -4673 -500 -4615 -488
rect -4415 488 -4357 500
rect -4415 -488 -4403 488
rect -4369 -488 -4357 488
rect -4415 -500 -4357 -488
rect -4157 488 -4099 500
rect -4157 -488 -4145 488
rect -4111 -488 -4099 488
rect -4157 -500 -4099 -488
rect -3899 488 -3841 500
rect -3899 -488 -3887 488
rect -3853 -488 -3841 488
rect -3899 -500 -3841 -488
rect -3641 488 -3583 500
rect -3641 -488 -3629 488
rect -3595 -488 -3583 488
rect -3641 -500 -3583 -488
rect -3383 488 -3325 500
rect -3383 -488 -3371 488
rect -3337 -488 -3325 488
rect -3383 -500 -3325 -488
rect -3125 488 -3067 500
rect -3125 -488 -3113 488
rect -3079 -488 -3067 488
rect -3125 -500 -3067 -488
rect -2867 488 -2809 500
rect -2867 -488 -2855 488
rect -2821 -488 -2809 488
rect -2867 -500 -2809 -488
rect -2609 488 -2551 500
rect -2609 -488 -2597 488
rect -2563 -488 -2551 488
rect -2609 -500 -2551 -488
rect -2351 488 -2293 500
rect -2351 -488 -2339 488
rect -2305 -488 -2293 488
rect -2351 -500 -2293 -488
rect -2093 488 -2035 500
rect -2093 -488 -2081 488
rect -2047 -488 -2035 488
rect -2093 -500 -2035 -488
rect -1835 488 -1777 500
rect -1835 -488 -1823 488
rect -1789 -488 -1777 488
rect -1835 -500 -1777 -488
rect -1577 488 -1519 500
rect -1577 -488 -1565 488
rect -1531 -488 -1519 488
rect -1577 -500 -1519 -488
rect -1319 488 -1261 500
rect -1319 -488 -1307 488
rect -1273 -488 -1261 488
rect -1319 -500 -1261 -488
rect -1061 488 -1003 500
rect -1061 -488 -1049 488
rect -1015 -488 -1003 488
rect -1061 -500 -1003 -488
rect -803 488 -745 500
rect -803 -488 -791 488
rect -757 -488 -745 488
rect -803 -500 -745 -488
rect -545 488 -487 500
rect -545 -488 -533 488
rect -499 -488 -487 488
rect -545 -500 -487 -488
rect -287 488 -229 500
rect -287 -488 -275 488
rect -241 -488 -229 488
rect -287 -500 -229 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 229 488 287 500
rect 229 -488 241 488
rect 275 -488 287 488
rect 229 -500 287 -488
rect 487 488 545 500
rect 487 -488 499 488
rect 533 -488 545 488
rect 487 -500 545 -488
rect 745 488 803 500
rect 745 -488 757 488
rect 791 -488 803 488
rect 745 -500 803 -488
rect 1003 488 1061 500
rect 1003 -488 1015 488
rect 1049 -488 1061 488
rect 1003 -500 1061 -488
rect 1261 488 1319 500
rect 1261 -488 1273 488
rect 1307 -488 1319 488
rect 1261 -500 1319 -488
rect 1519 488 1577 500
rect 1519 -488 1531 488
rect 1565 -488 1577 488
rect 1519 -500 1577 -488
rect 1777 488 1835 500
rect 1777 -488 1789 488
rect 1823 -488 1835 488
rect 1777 -500 1835 -488
rect 2035 488 2093 500
rect 2035 -488 2047 488
rect 2081 -488 2093 488
rect 2035 -500 2093 -488
rect 2293 488 2351 500
rect 2293 -488 2305 488
rect 2339 -488 2351 488
rect 2293 -500 2351 -488
rect 2551 488 2609 500
rect 2551 -488 2563 488
rect 2597 -488 2609 488
rect 2551 -500 2609 -488
rect 2809 488 2867 500
rect 2809 -488 2821 488
rect 2855 -488 2867 488
rect 2809 -500 2867 -488
rect 3067 488 3125 500
rect 3067 -488 3079 488
rect 3113 -488 3125 488
rect 3067 -500 3125 -488
rect 3325 488 3383 500
rect 3325 -488 3337 488
rect 3371 -488 3383 488
rect 3325 -500 3383 -488
rect 3583 488 3641 500
rect 3583 -488 3595 488
rect 3629 -488 3641 488
rect 3583 -500 3641 -488
rect 3841 488 3899 500
rect 3841 -488 3853 488
rect 3887 -488 3899 488
rect 3841 -500 3899 -488
rect 4099 488 4157 500
rect 4099 -488 4111 488
rect 4145 -488 4157 488
rect 4099 -500 4157 -488
rect 4357 488 4415 500
rect 4357 -488 4369 488
rect 4403 -488 4415 488
rect 4357 -500 4415 -488
rect 4615 488 4673 500
rect 4615 -488 4627 488
rect 4661 -488 4673 488
rect 4615 -500 4673 -488
rect 4873 488 4931 500
rect 4873 -488 4885 488
rect 4919 -488 4931 488
rect 4873 -500 4931 -488
rect 5131 488 5189 500
rect 5131 -488 5143 488
rect 5177 -488 5189 488
rect 5131 -500 5189 -488
rect 5389 488 5447 500
rect 5389 -488 5401 488
rect 5435 -488 5447 488
rect 5389 -500 5447 -488
rect 5647 488 5705 500
rect 5647 -488 5659 488
rect 5693 -488 5705 488
rect 5647 -500 5705 -488
rect -5705 -622 -5647 -610
rect -5705 -1598 -5693 -622
rect -5659 -1598 -5647 -622
rect -5705 -1610 -5647 -1598
rect -5447 -622 -5389 -610
rect -5447 -1598 -5435 -622
rect -5401 -1598 -5389 -622
rect -5447 -1610 -5389 -1598
rect -5189 -622 -5131 -610
rect -5189 -1598 -5177 -622
rect -5143 -1598 -5131 -622
rect -5189 -1610 -5131 -1598
rect -4931 -622 -4873 -610
rect -4931 -1598 -4919 -622
rect -4885 -1598 -4873 -622
rect -4931 -1610 -4873 -1598
rect -4673 -622 -4615 -610
rect -4673 -1598 -4661 -622
rect -4627 -1598 -4615 -622
rect -4673 -1610 -4615 -1598
rect -4415 -622 -4357 -610
rect -4415 -1598 -4403 -622
rect -4369 -1598 -4357 -622
rect -4415 -1610 -4357 -1598
rect -4157 -622 -4099 -610
rect -4157 -1598 -4145 -622
rect -4111 -1598 -4099 -622
rect -4157 -1610 -4099 -1598
rect -3899 -622 -3841 -610
rect -3899 -1598 -3887 -622
rect -3853 -1598 -3841 -622
rect -3899 -1610 -3841 -1598
rect -3641 -622 -3583 -610
rect -3641 -1598 -3629 -622
rect -3595 -1598 -3583 -622
rect -3641 -1610 -3583 -1598
rect -3383 -622 -3325 -610
rect -3383 -1598 -3371 -622
rect -3337 -1598 -3325 -622
rect -3383 -1610 -3325 -1598
rect -3125 -622 -3067 -610
rect -3125 -1598 -3113 -622
rect -3079 -1598 -3067 -622
rect -3125 -1610 -3067 -1598
rect -2867 -622 -2809 -610
rect -2867 -1598 -2855 -622
rect -2821 -1598 -2809 -622
rect -2867 -1610 -2809 -1598
rect -2609 -622 -2551 -610
rect -2609 -1598 -2597 -622
rect -2563 -1598 -2551 -622
rect -2609 -1610 -2551 -1598
rect -2351 -622 -2293 -610
rect -2351 -1598 -2339 -622
rect -2305 -1598 -2293 -622
rect -2351 -1610 -2293 -1598
rect -2093 -622 -2035 -610
rect -2093 -1598 -2081 -622
rect -2047 -1598 -2035 -622
rect -2093 -1610 -2035 -1598
rect -1835 -622 -1777 -610
rect -1835 -1598 -1823 -622
rect -1789 -1598 -1777 -622
rect -1835 -1610 -1777 -1598
rect -1577 -622 -1519 -610
rect -1577 -1598 -1565 -622
rect -1531 -1598 -1519 -622
rect -1577 -1610 -1519 -1598
rect -1319 -622 -1261 -610
rect -1319 -1598 -1307 -622
rect -1273 -1598 -1261 -622
rect -1319 -1610 -1261 -1598
rect -1061 -622 -1003 -610
rect -1061 -1598 -1049 -622
rect -1015 -1598 -1003 -622
rect -1061 -1610 -1003 -1598
rect -803 -622 -745 -610
rect -803 -1598 -791 -622
rect -757 -1598 -745 -622
rect -803 -1610 -745 -1598
rect -545 -622 -487 -610
rect -545 -1598 -533 -622
rect -499 -1598 -487 -622
rect -545 -1610 -487 -1598
rect -287 -622 -229 -610
rect -287 -1598 -275 -622
rect -241 -1598 -229 -622
rect -287 -1610 -229 -1598
rect -29 -622 29 -610
rect -29 -1598 -17 -622
rect 17 -1598 29 -622
rect -29 -1610 29 -1598
rect 229 -622 287 -610
rect 229 -1598 241 -622
rect 275 -1598 287 -622
rect 229 -1610 287 -1598
rect 487 -622 545 -610
rect 487 -1598 499 -622
rect 533 -1598 545 -622
rect 487 -1610 545 -1598
rect 745 -622 803 -610
rect 745 -1598 757 -622
rect 791 -1598 803 -622
rect 745 -1610 803 -1598
rect 1003 -622 1061 -610
rect 1003 -1598 1015 -622
rect 1049 -1598 1061 -622
rect 1003 -1610 1061 -1598
rect 1261 -622 1319 -610
rect 1261 -1598 1273 -622
rect 1307 -1598 1319 -622
rect 1261 -1610 1319 -1598
rect 1519 -622 1577 -610
rect 1519 -1598 1531 -622
rect 1565 -1598 1577 -622
rect 1519 -1610 1577 -1598
rect 1777 -622 1835 -610
rect 1777 -1598 1789 -622
rect 1823 -1598 1835 -622
rect 1777 -1610 1835 -1598
rect 2035 -622 2093 -610
rect 2035 -1598 2047 -622
rect 2081 -1598 2093 -622
rect 2035 -1610 2093 -1598
rect 2293 -622 2351 -610
rect 2293 -1598 2305 -622
rect 2339 -1598 2351 -622
rect 2293 -1610 2351 -1598
rect 2551 -622 2609 -610
rect 2551 -1598 2563 -622
rect 2597 -1598 2609 -622
rect 2551 -1610 2609 -1598
rect 2809 -622 2867 -610
rect 2809 -1598 2821 -622
rect 2855 -1598 2867 -622
rect 2809 -1610 2867 -1598
rect 3067 -622 3125 -610
rect 3067 -1598 3079 -622
rect 3113 -1598 3125 -622
rect 3067 -1610 3125 -1598
rect 3325 -622 3383 -610
rect 3325 -1598 3337 -622
rect 3371 -1598 3383 -622
rect 3325 -1610 3383 -1598
rect 3583 -622 3641 -610
rect 3583 -1598 3595 -622
rect 3629 -1598 3641 -622
rect 3583 -1610 3641 -1598
rect 3841 -622 3899 -610
rect 3841 -1598 3853 -622
rect 3887 -1598 3899 -622
rect 3841 -1610 3899 -1598
rect 4099 -622 4157 -610
rect 4099 -1598 4111 -622
rect 4145 -1598 4157 -622
rect 4099 -1610 4157 -1598
rect 4357 -622 4415 -610
rect 4357 -1598 4369 -622
rect 4403 -1598 4415 -622
rect 4357 -1610 4415 -1598
rect 4615 -622 4673 -610
rect 4615 -1598 4627 -622
rect 4661 -1598 4673 -622
rect 4615 -1610 4673 -1598
rect 4873 -622 4931 -610
rect 4873 -1598 4885 -622
rect 4919 -1598 4931 -622
rect 4873 -1610 4931 -1598
rect 5131 -622 5189 -610
rect 5131 -1598 5143 -622
rect 5177 -1598 5189 -622
rect 5131 -1610 5189 -1598
rect 5389 -622 5447 -610
rect 5389 -1598 5401 -622
rect 5435 -1598 5447 -622
rect 5389 -1610 5447 -1598
rect 5647 -622 5705 -610
rect 5647 -1598 5659 -622
rect 5693 -1598 5705 -622
rect 5647 -1610 5705 -1598
rect -5705 -1732 -5647 -1720
rect -5705 -2708 -5693 -1732
rect -5659 -2708 -5647 -1732
rect -5705 -2720 -5647 -2708
rect -5447 -1732 -5389 -1720
rect -5447 -2708 -5435 -1732
rect -5401 -2708 -5389 -1732
rect -5447 -2720 -5389 -2708
rect -5189 -1732 -5131 -1720
rect -5189 -2708 -5177 -1732
rect -5143 -2708 -5131 -1732
rect -5189 -2720 -5131 -2708
rect -4931 -1732 -4873 -1720
rect -4931 -2708 -4919 -1732
rect -4885 -2708 -4873 -1732
rect -4931 -2720 -4873 -2708
rect -4673 -1732 -4615 -1720
rect -4673 -2708 -4661 -1732
rect -4627 -2708 -4615 -1732
rect -4673 -2720 -4615 -2708
rect -4415 -1732 -4357 -1720
rect -4415 -2708 -4403 -1732
rect -4369 -2708 -4357 -1732
rect -4415 -2720 -4357 -2708
rect -4157 -1732 -4099 -1720
rect -4157 -2708 -4145 -1732
rect -4111 -2708 -4099 -1732
rect -4157 -2720 -4099 -2708
rect -3899 -1732 -3841 -1720
rect -3899 -2708 -3887 -1732
rect -3853 -2708 -3841 -1732
rect -3899 -2720 -3841 -2708
rect -3641 -1732 -3583 -1720
rect -3641 -2708 -3629 -1732
rect -3595 -2708 -3583 -1732
rect -3641 -2720 -3583 -2708
rect -3383 -1732 -3325 -1720
rect -3383 -2708 -3371 -1732
rect -3337 -2708 -3325 -1732
rect -3383 -2720 -3325 -2708
rect -3125 -1732 -3067 -1720
rect -3125 -2708 -3113 -1732
rect -3079 -2708 -3067 -1732
rect -3125 -2720 -3067 -2708
rect -2867 -1732 -2809 -1720
rect -2867 -2708 -2855 -1732
rect -2821 -2708 -2809 -1732
rect -2867 -2720 -2809 -2708
rect -2609 -1732 -2551 -1720
rect -2609 -2708 -2597 -1732
rect -2563 -2708 -2551 -1732
rect -2609 -2720 -2551 -2708
rect -2351 -1732 -2293 -1720
rect -2351 -2708 -2339 -1732
rect -2305 -2708 -2293 -1732
rect -2351 -2720 -2293 -2708
rect -2093 -1732 -2035 -1720
rect -2093 -2708 -2081 -1732
rect -2047 -2708 -2035 -1732
rect -2093 -2720 -2035 -2708
rect -1835 -1732 -1777 -1720
rect -1835 -2708 -1823 -1732
rect -1789 -2708 -1777 -1732
rect -1835 -2720 -1777 -2708
rect -1577 -1732 -1519 -1720
rect -1577 -2708 -1565 -1732
rect -1531 -2708 -1519 -1732
rect -1577 -2720 -1519 -2708
rect -1319 -1732 -1261 -1720
rect -1319 -2708 -1307 -1732
rect -1273 -2708 -1261 -1732
rect -1319 -2720 -1261 -2708
rect -1061 -1732 -1003 -1720
rect -1061 -2708 -1049 -1732
rect -1015 -2708 -1003 -1732
rect -1061 -2720 -1003 -2708
rect -803 -1732 -745 -1720
rect -803 -2708 -791 -1732
rect -757 -2708 -745 -1732
rect -803 -2720 -745 -2708
rect -545 -1732 -487 -1720
rect -545 -2708 -533 -1732
rect -499 -2708 -487 -1732
rect -545 -2720 -487 -2708
rect -287 -1732 -229 -1720
rect -287 -2708 -275 -1732
rect -241 -2708 -229 -1732
rect -287 -2720 -229 -2708
rect -29 -1732 29 -1720
rect -29 -2708 -17 -1732
rect 17 -2708 29 -1732
rect -29 -2720 29 -2708
rect 229 -1732 287 -1720
rect 229 -2708 241 -1732
rect 275 -2708 287 -1732
rect 229 -2720 287 -2708
rect 487 -1732 545 -1720
rect 487 -2708 499 -1732
rect 533 -2708 545 -1732
rect 487 -2720 545 -2708
rect 745 -1732 803 -1720
rect 745 -2708 757 -1732
rect 791 -2708 803 -1732
rect 745 -2720 803 -2708
rect 1003 -1732 1061 -1720
rect 1003 -2708 1015 -1732
rect 1049 -2708 1061 -1732
rect 1003 -2720 1061 -2708
rect 1261 -1732 1319 -1720
rect 1261 -2708 1273 -1732
rect 1307 -2708 1319 -1732
rect 1261 -2720 1319 -2708
rect 1519 -1732 1577 -1720
rect 1519 -2708 1531 -1732
rect 1565 -2708 1577 -1732
rect 1519 -2720 1577 -2708
rect 1777 -1732 1835 -1720
rect 1777 -2708 1789 -1732
rect 1823 -2708 1835 -1732
rect 1777 -2720 1835 -2708
rect 2035 -1732 2093 -1720
rect 2035 -2708 2047 -1732
rect 2081 -2708 2093 -1732
rect 2035 -2720 2093 -2708
rect 2293 -1732 2351 -1720
rect 2293 -2708 2305 -1732
rect 2339 -2708 2351 -1732
rect 2293 -2720 2351 -2708
rect 2551 -1732 2609 -1720
rect 2551 -2708 2563 -1732
rect 2597 -2708 2609 -1732
rect 2551 -2720 2609 -2708
rect 2809 -1732 2867 -1720
rect 2809 -2708 2821 -1732
rect 2855 -2708 2867 -1732
rect 2809 -2720 2867 -2708
rect 3067 -1732 3125 -1720
rect 3067 -2708 3079 -1732
rect 3113 -2708 3125 -1732
rect 3067 -2720 3125 -2708
rect 3325 -1732 3383 -1720
rect 3325 -2708 3337 -1732
rect 3371 -2708 3383 -1732
rect 3325 -2720 3383 -2708
rect 3583 -1732 3641 -1720
rect 3583 -2708 3595 -1732
rect 3629 -2708 3641 -1732
rect 3583 -2720 3641 -2708
rect 3841 -1732 3899 -1720
rect 3841 -2708 3853 -1732
rect 3887 -2708 3899 -1732
rect 3841 -2720 3899 -2708
rect 4099 -1732 4157 -1720
rect 4099 -2708 4111 -1732
rect 4145 -2708 4157 -1732
rect 4099 -2720 4157 -2708
rect 4357 -1732 4415 -1720
rect 4357 -2708 4369 -1732
rect 4403 -2708 4415 -1732
rect 4357 -2720 4415 -2708
rect 4615 -1732 4673 -1720
rect 4615 -2708 4627 -1732
rect 4661 -2708 4673 -1732
rect 4615 -2720 4673 -2708
rect 4873 -1732 4931 -1720
rect 4873 -2708 4885 -1732
rect 4919 -2708 4931 -1732
rect 4873 -2720 4931 -2708
rect 5131 -1732 5189 -1720
rect 5131 -2708 5143 -1732
rect 5177 -2708 5189 -1732
rect 5131 -2720 5189 -2708
rect 5389 -1732 5447 -1720
rect 5389 -2708 5401 -1732
rect 5435 -2708 5447 -1732
rect 5389 -2720 5447 -2708
rect 5647 -1732 5705 -1720
rect 5647 -2708 5659 -1732
rect 5693 -2708 5705 -1732
rect 5647 -2720 5705 -2708
<< mvndiffc >>
rect -5693 1732 -5659 2708
rect -5435 1732 -5401 2708
rect -5177 1732 -5143 2708
rect -4919 1732 -4885 2708
rect -4661 1732 -4627 2708
rect -4403 1732 -4369 2708
rect -4145 1732 -4111 2708
rect -3887 1732 -3853 2708
rect -3629 1732 -3595 2708
rect -3371 1732 -3337 2708
rect -3113 1732 -3079 2708
rect -2855 1732 -2821 2708
rect -2597 1732 -2563 2708
rect -2339 1732 -2305 2708
rect -2081 1732 -2047 2708
rect -1823 1732 -1789 2708
rect -1565 1732 -1531 2708
rect -1307 1732 -1273 2708
rect -1049 1732 -1015 2708
rect -791 1732 -757 2708
rect -533 1732 -499 2708
rect -275 1732 -241 2708
rect -17 1732 17 2708
rect 241 1732 275 2708
rect 499 1732 533 2708
rect 757 1732 791 2708
rect 1015 1732 1049 2708
rect 1273 1732 1307 2708
rect 1531 1732 1565 2708
rect 1789 1732 1823 2708
rect 2047 1732 2081 2708
rect 2305 1732 2339 2708
rect 2563 1732 2597 2708
rect 2821 1732 2855 2708
rect 3079 1732 3113 2708
rect 3337 1732 3371 2708
rect 3595 1732 3629 2708
rect 3853 1732 3887 2708
rect 4111 1732 4145 2708
rect 4369 1732 4403 2708
rect 4627 1732 4661 2708
rect 4885 1732 4919 2708
rect 5143 1732 5177 2708
rect 5401 1732 5435 2708
rect 5659 1732 5693 2708
rect -5693 622 -5659 1598
rect -5435 622 -5401 1598
rect -5177 622 -5143 1598
rect -4919 622 -4885 1598
rect -4661 622 -4627 1598
rect -4403 622 -4369 1598
rect -4145 622 -4111 1598
rect -3887 622 -3853 1598
rect -3629 622 -3595 1598
rect -3371 622 -3337 1598
rect -3113 622 -3079 1598
rect -2855 622 -2821 1598
rect -2597 622 -2563 1598
rect -2339 622 -2305 1598
rect -2081 622 -2047 1598
rect -1823 622 -1789 1598
rect -1565 622 -1531 1598
rect -1307 622 -1273 1598
rect -1049 622 -1015 1598
rect -791 622 -757 1598
rect -533 622 -499 1598
rect -275 622 -241 1598
rect -17 622 17 1598
rect 241 622 275 1598
rect 499 622 533 1598
rect 757 622 791 1598
rect 1015 622 1049 1598
rect 1273 622 1307 1598
rect 1531 622 1565 1598
rect 1789 622 1823 1598
rect 2047 622 2081 1598
rect 2305 622 2339 1598
rect 2563 622 2597 1598
rect 2821 622 2855 1598
rect 3079 622 3113 1598
rect 3337 622 3371 1598
rect 3595 622 3629 1598
rect 3853 622 3887 1598
rect 4111 622 4145 1598
rect 4369 622 4403 1598
rect 4627 622 4661 1598
rect 4885 622 4919 1598
rect 5143 622 5177 1598
rect 5401 622 5435 1598
rect 5659 622 5693 1598
rect -5693 -488 -5659 488
rect -5435 -488 -5401 488
rect -5177 -488 -5143 488
rect -4919 -488 -4885 488
rect -4661 -488 -4627 488
rect -4403 -488 -4369 488
rect -4145 -488 -4111 488
rect -3887 -488 -3853 488
rect -3629 -488 -3595 488
rect -3371 -488 -3337 488
rect -3113 -488 -3079 488
rect -2855 -488 -2821 488
rect -2597 -488 -2563 488
rect -2339 -488 -2305 488
rect -2081 -488 -2047 488
rect -1823 -488 -1789 488
rect -1565 -488 -1531 488
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
rect 1531 -488 1565 488
rect 1789 -488 1823 488
rect 2047 -488 2081 488
rect 2305 -488 2339 488
rect 2563 -488 2597 488
rect 2821 -488 2855 488
rect 3079 -488 3113 488
rect 3337 -488 3371 488
rect 3595 -488 3629 488
rect 3853 -488 3887 488
rect 4111 -488 4145 488
rect 4369 -488 4403 488
rect 4627 -488 4661 488
rect 4885 -488 4919 488
rect 5143 -488 5177 488
rect 5401 -488 5435 488
rect 5659 -488 5693 488
rect -5693 -1598 -5659 -622
rect -5435 -1598 -5401 -622
rect -5177 -1598 -5143 -622
rect -4919 -1598 -4885 -622
rect -4661 -1598 -4627 -622
rect -4403 -1598 -4369 -622
rect -4145 -1598 -4111 -622
rect -3887 -1598 -3853 -622
rect -3629 -1598 -3595 -622
rect -3371 -1598 -3337 -622
rect -3113 -1598 -3079 -622
rect -2855 -1598 -2821 -622
rect -2597 -1598 -2563 -622
rect -2339 -1598 -2305 -622
rect -2081 -1598 -2047 -622
rect -1823 -1598 -1789 -622
rect -1565 -1598 -1531 -622
rect -1307 -1598 -1273 -622
rect -1049 -1598 -1015 -622
rect -791 -1598 -757 -622
rect -533 -1598 -499 -622
rect -275 -1598 -241 -622
rect -17 -1598 17 -622
rect 241 -1598 275 -622
rect 499 -1598 533 -622
rect 757 -1598 791 -622
rect 1015 -1598 1049 -622
rect 1273 -1598 1307 -622
rect 1531 -1598 1565 -622
rect 1789 -1598 1823 -622
rect 2047 -1598 2081 -622
rect 2305 -1598 2339 -622
rect 2563 -1598 2597 -622
rect 2821 -1598 2855 -622
rect 3079 -1598 3113 -622
rect 3337 -1598 3371 -622
rect 3595 -1598 3629 -622
rect 3853 -1598 3887 -622
rect 4111 -1598 4145 -622
rect 4369 -1598 4403 -622
rect 4627 -1598 4661 -622
rect 4885 -1598 4919 -622
rect 5143 -1598 5177 -622
rect 5401 -1598 5435 -622
rect 5659 -1598 5693 -622
rect -5693 -2708 -5659 -1732
rect -5435 -2708 -5401 -1732
rect -5177 -2708 -5143 -1732
rect -4919 -2708 -4885 -1732
rect -4661 -2708 -4627 -1732
rect -4403 -2708 -4369 -1732
rect -4145 -2708 -4111 -1732
rect -3887 -2708 -3853 -1732
rect -3629 -2708 -3595 -1732
rect -3371 -2708 -3337 -1732
rect -3113 -2708 -3079 -1732
rect -2855 -2708 -2821 -1732
rect -2597 -2708 -2563 -1732
rect -2339 -2708 -2305 -1732
rect -2081 -2708 -2047 -1732
rect -1823 -2708 -1789 -1732
rect -1565 -2708 -1531 -1732
rect -1307 -2708 -1273 -1732
rect -1049 -2708 -1015 -1732
rect -791 -2708 -757 -1732
rect -533 -2708 -499 -1732
rect -275 -2708 -241 -1732
rect -17 -2708 17 -1732
rect 241 -2708 275 -1732
rect 499 -2708 533 -1732
rect 757 -2708 791 -1732
rect 1015 -2708 1049 -1732
rect 1273 -2708 1307 -1732
rect 1531 -2708 1565 -1732
rect 1789 -2708 1823 -1732
rect 2047 -2708 2081 -1732
rect 2305 -2708 2339 -1732
rect 2563 -2708 2597 -1732
rect 2821 -2708 2855 -1732
rect 3079 -2708 3113 -1732
rect 3337 -2708 3371 -1732
rect 3595 -2708 3629 -1732
rect 3853 -2708 3887 -1732
rect 4111 -2708 4145 -1732
rect 4369 -2708 4403 -1732
rect 4627 -2708 4661 -1732
rect 4885 -2708 4919 -1732
rect 5143 -2708 5177 -1732
rect 5401 -2708 5435 -1732
rect 5659 -2708 5693 -1732
<< mvpsubdiff >>
rect -5839 2930 5839 2942
rect -5839 2896 -5731 2930
rect 5731 2896 5839 2930
rect -5839 2884 5839 2896
rect -5839 2834 -5781 2884
rect -5839 -2834 -5827 2834
rect -5793 -2834 -5781 2834
rect 5781 2834 5839 2884
rect -5839 -2884 -5781 -2834
rect 5781 -2834 5793 2834
rect 5827 -2834 5839 2834
rect 5781 -2884 5839 -2834
rect -5839 -2896 5839 -2884
rect -5839 -2930 -5731 -2896
rect 5731 -2930 5839 -2896
rect -5839 -2942 5839 -2930
<< mvpsubdiffcont >>
rect -5731 2896 5731 2930
rect -5827 -2834 -5793 2834
rect 5793 -2834 5827 2834
rect -5731 -2930 5731 -2896
<< poly >>
rect -5647 2792 -5447 2808
rect -5647 2758 -5631 2792
rect -5463 2758 -5447 2792
rect -5647 2720 -5447 2758
rect -5389 2792 -5189 2808
rect -5389 2758 -5373 2792
rect -5205 2758 -5189 2792
rect -5389 2720 -5189 2758
rect -5131 2792 -4931 2808
rect -5131 2758 -5115 2792
rect -4947 2758 -4931 2792
rect -5131 2720 -4931 2758
rect -4873 2792 -4673 2808
rect -4873 2758 -4857 2792
rect -4689 2758 -4673 2792
rect -4873 2720 -4673 2758
rect -4615 2792 -4415 2808
rect -4615 2758 -4599 2792
rect -4431 2758 -4415 2792
rect -4615 2720 -4415 2758
rect -4357 2792 -4157 2808
rect -4357 2758 -4341 2792
rect -4173 2758 -4157 2792
rect -4357 2720 -4157 2758
rect -4099 2792 -3899 2808
rect -4099 2758 -4083 2792
rect -3915 2758 -3899 2792
rect -4099 2720 -3899 2758
rect -3841 2792 -3641 2808
rect -3841 2758 -3825 2792
rect -3657 2758 -3641 2792
rect -3841 2720 -3641 2758
rect -3583 2792 -3383 2808
rect -3583 2758 -3567 2792
rect -3399 2758 -3383 2792
rect -3583 2720 -3383 2758
rect -3325 2792 -3125 2808
rect -3325 2758 -3309 2792
rect -3141 2758 -3125 2792
rect -3325 2720 -3125 2758
rect -3067 2792 -2867 2808
rect -3067 2758 -3051 2792
rect -2883 2758 -2867 2792
rect -3067 2720 -2867 2758
rect -2809 2792 -2609 2808
rect -2809 2758 -2793 2792
rect -2625 2758 -2609 2792
rect -2809 2720 -2609 2758
rect -2551 2792 -2351 2808
rect -2551 2758 -2535 2792
rect -2367 2758 -2351 2792
rect -2551 2720 -2351 2758
rect -2293 2792 -2093 2808
rect -2293 2758 -2277 2792
rect -2109 2758 -2093 2792
rect -2293 2720 -2093 2758
rect -2035 2792 -1835 2808
rect -2035 2758 -2019 2792
rect -1851 2758 -1835 2792
rect -2035 2720 -1835 2758
rect -1777 2792 -1577 2808
rect -1777 2758 -1761 2792
rect -1593 2758 -1577 2792
rect -1777 2720 -1577 2758
rect -1519 2792 -1319 2808
rect -1519 2758 -1503 2792
rect -1335 2758 -1319 2792
rect -1519 2720 -1319 2758
rect -1261 2792 -1061 2808
rect -1261 2758 -1245 2792
rect -1077 2758 -1061 2792
rect -1261 2720 -1061 2758
rect -1003 2792 -803 2808
rect -1003 2758 -987 2792
rect -819 2758 -803 2792
rect -1003 2720 -803 2758
rect -745 2792 -545 2808
rect -745 2758 -729 2792
rect -561 2758 -545 2792
rect -745 2720 -545 2758
rect -487 2792 -287 2808
rect -487 2758 -471 2792
rect -303 2758 -287 2792
rect -487 2720 -287 2758
rect -229 2792 -29 2808
rect -229 2758 -213 2792
rect -45 2758 -29 2792
rect -229 2720 -29 2758
rect 29 2792 229 2808
rect 29 2758 45 2792
rect 213 2758 229 2792
rect 29 2720 229 2758
rect 287 2792 487 2808
rect 287 2758 303 2792
rect 471 2758 487 2792
rect 287 2720 487 2758
rect 545 2792 745 2808
rect 545 2758 561 2792
rect 729 2758 745 2792
rect 545 2720 745 2758
rect 803 2792 1003 2808
rect 803 2758 819 2792
rect 987 2758 1003 2792
rect 803 2720 1003 2758
rect 1061 2792 1261 2808
rect 1061 2758 1077 2792
rect 1245 2758 1261 2792
rect 1061 2720 1261 2758
rect 1319 2792 1519 2808
rect 1319 2758 1335 2792
rect 1503 2758 1519 2792
rect 1319 2720 1519 2758
rect 1577 2792 1777 2808
rect 1577 2758 1593 2792
rect 1761 2758 1777 2792
rect 1577 2720 1777 2758
rect 1835 2792 2035 2808
rect 1835 2758 1851 2792
rect 2019 2758 2035 2792
rect 1835 2720 2035 2758
rect 2093 2792 2293 2808
rect 2093 2758 2109 2792
rect 2277 2758 2293 2792
rect 2093 2720 2293 2758
rect 2351 2792 2551 2808
rect 2351 2758 2367 2792
rect 2535 2758 2551 2792
rect 2351 2720 2551 2758
rect 2609 2792 2809 2808
rect 2609 2758 2625 2792
rect 2793 2758 2809 2792
rect 2609 2720 2809 2758
rect 2867 2792 3067 2808
rect 2867 2758 2883 2792
rect 3051 2758 3067 2792
rect 2867 2720 3067 2758
rect 3125 2792 3325 2808
rect 3125 2758 3141 2792
rect 3309 2758 3325 2792
rect 3125 2720 3325 2758
rect 3383 2792 3583 2808
rect 3383 2758 3399 2792
rect 3567 2758 3583 2792
rect 3383 2720 3583 2758
rect 3641 2792 3841 2808
rect 3641 2758 3657 2792
rect 3825 2758 3841 2792
rect 3641 2720 3841 2758
rect 3899 2792 4099 2808
rect 3899 2758 3915 2792
rect 4083 2758 4099 2792
rect 3899 2720 4099 2758
rect 4157 2792 4357 2808
rect 4157 2758 4173 2792
rect 4341 2758 4357 2792
rect 4157 2720 4357 2758
rect 4415 2792 4615 2808
rect 4415 2758 4431 2792
rect 4599 2758 4615 2792
rect 4415 2720 4615 2758
rect 4673 2792 4873 2808
rect 4673 2758 4689 2792
rect 4857 2758 4873 2792
rect 4673 2720 4873 2758
rect 4931 2792 5131 2808
rect 4931 2758 4947 2792
rect 5115 2758 5131 2792
rect 4931 2720 5131 2758
rect 5189 2792 5389 2808
rect 5189 2758 5205 2792
rect 5373 2758 5389 2792
rect 5189 2720 5389 2758
rect 5447 2792 5647 2808
rect 5447 2758 5463 2792
rect 5631 2758 5647 2792
rect 5447 2720 5647 2758
rect -5647 1682 -5447 1720
rect -5647 1648 -5631 1682
rect -5463 1648 -5447 1682
rect -5647 1610 -5447 1648
rect -5389 1682 -5189 1720
rect -5389 1648 -5373 1682
rect -5205 1648 -5189 1682
rect -5389 1610 -5189 1648
rect -5131 1682 -4931 1720
rect -5131 1648 -5115 1682
rect -4947 1648 -4931 1682
rect -5131 1610 -4931 1648
rect -4873 1682 -4673 1720
rect -4873 1648 -4857 1682
rect -4689 1648 -4673 1682
rect -4873 1610 -4673 1648
rect -4615 1682 -4415 1720
rect -4615 1648 -4599 1682
rect -4431 1648 -4415 1682
rect -4615 1610 -4415 1648
rect -4357 1682 -4157 1720
rect -4357 1648 -4341 1682
rect -4173 1648 -4157 1682
rect -4357 1610 -4157 1648
rect -4099 1682 -3899 1720
rect -4099 1648 -4083 1682
rect -3915 1648 -3899 1682
rect -4099 1610 -3899 1648
rect -3841 1682 -3641 1720
rect -3841 1648 -3825 1682
rect -3657 1648 -3641 1682
rect -3841 1610 -3641 1648
rect -3583 1682 -3383 1720
rect -3583 1648 -3567 1682
rect -3399 1648 -3383 1682
rect -3583 1610 -3383 1648
rect -3325 1682 -3125 1720
rect -3325 1648 -3309 1682
rect -3141 1648 -3125 1682
rect -3325 1610 -3125 1648
rect -3067 1682 -2867 1720
rect -3067 1648 -3051 1682
rect -2883 1648 -2867 1682
rect -3067 1610 -2867 1648
rect -2809 1682 -2609 1720
rect -2809 1648 -2793 1682
rect -2625 1648 -2609 1682
rect -2809 1610 -2609 1648
rect -2551 1682 -2351 1720
rect -2551 1648 -2535 1682
rect -2367 1648 -2351 1682
rect -2551 1610 -2351 1648
rect -2293 1682 -2093 1720
rect -2293 1648 -2277 1682
rect -2109 1648 -2093 1682
rect -2293 1610 -2093 1648
rect -2035 1682 -1835 1720
rect -2035 1648 -2019 1682
rect -1851 1648 -1835 1682
rect -2035 1610 -1835 1648
rect -1777 1682 -1577 1720
rect -1777 1648 -1761 1682
rect -1593 1648 -1577 1682
rect -1777 1610 -1577 1648
rect -1519 1682 -1319 1720
rect -1519 1648 -1503 1682
rect -1335 1648 -1319 1682
rect -1519 1610 -1319 1648
rect -1261 1682 -1061 1720
rect -1261 1648 -1245 1682
rect -1077 1648 -1061 1682
rect -1261 1610 -1061 1648
rect -1003 1682 -803 1720
rect -1003 1648 -987 1682
rect -819 1648 -803 1682
rect -1003 1610 -803 1648
rect -745 1682 -545 1720
rect -745 1648 -729 1682
rect -561 1648 -545 1682
rect -745 1610 -545 1648
rect -487 1682 -287 1720
rect -487 1648 -471 1682
rect -303 1648 -287 1682
rect -487 1610 -287 1648
rect -229 1682 -29 1720
rect -229 1648 -213 1682
rect -45 1648 -29 1682
rect -229 1610 -29 1648
rect 29 1682 229 1720
rect 29 1648 45 1682
rect 213 1648 229 1682
rect 29 1610 229 1648
rect 287 1682 487 1720
rect 287 1648 303 1682
rect 471 1648 487 1682
rect 287 1610 487 1648
rect 545 1682 745 1720
rect 545 1648 561 1682
rect 729 1648 745 1682
rect 545 1610 745 1648
rect 803 1682 1003 1720
rect 803 1648 819 1682
rect 987 1648 1003 1682
rect 803 1610 1003 1648
rect 1061 1682 1261 1720
rect 1061 1648 1077 1682
rect 1245 1648 1261 1682
rect 1061 1610 1261 1648
rect 1319 1682 1519 1720
rect 1319 1648 1335 1682
rect 1503 1648 1519 1682
rect 1319 1610 1519 1648
rect 1577 1682 1777 1720
rect 1577 1648 1593 1682
rect 1761 1648 1777 1682
rect 1577 1610 1777 1648
rect 1835 1682 2035 1720
rect 1835 1648 1851 1682
rect 2019 1648 2035 1682
rect 1835 1610 2035 1648
rect 2093 1682 2293 1720
rect 2093 1648 2109 1682
rect 2277 1648 2293 1682
rect 2093 1610 2293 1648
rect 2351 1682 2551 1720
rect 2351 1648 2367 1682
rect 2535 1648 2551 1682
rect 2351 1610 2551 1648
rect 2609 1682 2809 1720
rect 2609 1648 2625 1682
rect 2793 1648 2809 1682
rect 2609 1610 2809 1648
rect 2867 1682 3067 1720
rect 2867 1648 2883 1682
rect 3051 1648 3067 1682
rect 2867 1610 3067 1648
rect 3125 1682 3325 1720
rect 3125 1648 3141 1682
rect 3309 1648 3325 1682
rect 3125 1610 3325 1648
rect 3383 1682 3583 1720
rect 3383 1648 3399 1682
rect 3567 1648 3583 1682
rect 3383 1610 3583 1648
rect 3641 1682 3841 1720
rect 3641 1648 3657 1682
rect 3825 1648 3841 1682
rect 3641 1610 3841 1648
rect 3899 1682 4099 1720
rect 3899 1648 3915 1682
rect 4083 1648 4099 1682
rect 3899 1610 4099 1648
rect 4157 1682 4357 1720
rect 4157 1648 4173 1682
rect 4341 1648 4357 1682
rect 4157 1610 4357 1648
rect 4415 1682 4615 1720
rect 4415 1648 4431 1682
rect 4599 1648 4615 1682
rect 4415 1610 4615 1648
rect 4673 1682 4873 1720
rect 4673 1648 4689 1682
rect 4857 1648 4873 1682
rect 4673 1610 4873 1648
rect 4931 1682 5131 1720
rect 4931 1648 4947 1682
rect 5115 1648 5131 1682
rect 4931 1610 5131 1648
rect 5189 1682 5389 1720
rect 5189 1648 5205 1682
rect 5373 1648 5389 1682
rect 5189 1610 5389 1648
rect 5447 1682 5647 1720
rect 5447 1648 5463 1682
rect 5631 1648 5647 1682
rect 5447 1610 5647 1648
rect -5647 572 -5447 610
rect -5647 538 -5631 572
rect -5463 538 -5447 572
rect -5647 500 -5447 538
rect -5389 572 -5189 610
rect -5389 538 -5373 572
rect -5205 538 -5189 572
rect -5389 500 -5189 538
rect -5131 572 -4931 610
rect -5131 538 -5115 572
rect -4947 538 -4931 572
rect -5131 500 -4931 538
rect -4873 572 -4673 610
rect -4873 538 -4857 572
rect -4689 538 -4673 572
rect -4873 500 -4673 538
rect -4615 572 -4415 610
rect -4615 538 -4599 572
rect -4431 538 -4415 572
rect -4615 500 -4415 538
rect -4357 572 -4157 610
rect -4357 538 -4341 572
rect -4173 538 -4157 572
rect -4357 500 -4157 538
rect -4099 572 -3899 610
rect -4099 538 -4083 572
rect -3915 538 -3899 572
rect -4099 500 -3899 538
rect -3841 572 -3641 610
rect -3841 538 -3825 572
rect -3657 538 -3641 572
rect -3841 500 -3641 538
rect -3583 572 -3383 610
rect -3583 538 -3567 572
rect -3399 538 -3383 572
rect -3583 500 -3383 538
rect -3325 572 -3125 610
rect -3325 538 -3309 572
rect -3141 538 -3125 572
rect -3325 500 -3125 538
rect -3067 572 -2867 610
rect -3067 538 -3051 572
rect -2883 538 -2867 572
rect -3067 500 -2867 538
rect -2809 572 -2609 610
rect -2809 538 -2793 572
rect -2625 538 -2609 572
rect -2809 500 -2609 538
rect -2551 572 -2351 610
rect -2551 538 -2535 572
rect -2367 538 -2351 572
rect -2551 500 -2351 538
rect -2293 572 -2093 610
rect -2293 538 -2277 572
rect -2109 538 -2093 572
rect -2293 500 -2093 538
rect -2035 572 -1835 610
rect -2035 538 -2019 572
rect -1851 538 -1835 572
rect -2035 500 -1835 538
rect -1777 572 -1577 610
rect -1777 538 -1761 572
rect -1593 538 -1577 572
rect -1777 500 -1577 538
rect -1519 572 -1319 610
rect -1519 538 -1503 572
rect -1335 538 -1319 572
rect -1519 500 -1319 538
rect -1261 572 -1061 610
rect -1261 538 -1245 572
rect -1077 538 -1061 572
rect -1261 500 -1061 538
rect -1003 572 -803 610
rect -1003 538 -987 572
rect -819 538 -803 572
rect -1003 500 -803 538
rect -745 572 -545 610
rect -745 538 -729 572
rect -561 538 -545 572
rect -745 500 -545 538
rect -487 572 -287 610
rect -487 538 -471 572
rect -303 538 -287 572
rect -487 500 -287 538
rect -229 572 -29 610
rect -229 538 -213 572
rect -45 538 -29 572
rect -229 500 -29 538
rect 29 572 229 610
rect 29 538 45 572
rect 213 538 229 572
rect 29 500 229 538
rect 287 572 487 610
rect 287 538 303 572
rect 471 538 487 572
rect 287 500 487 538
rect 545 572 745 610
rect 545 538 561 572
rect 729 538 745 572
rect 545 500 745 538
rect 803 572 1003 610
rect 803 538 819 572
rect 987 538 1003 572
rect 803 500 1003 538
rect 1061 572 1261 610
rect 1061 538 1077 572
rect 1245 538 1261 572
rect 1061 500 1261 538
rect 1319 572 1519 610
rect 1319 538 1335 572
rect 1503 538 1519 572
rect 1319 500 1519 538
rect 1577 572 1777 610
rect 1577 538 1593 572
rect 1761 538 1777 572
rect 1577 500 1777 538
rect 1835 572 2035 610
rect 1835 538 1851 572
rect 2019 538 2035 572
rect 1835 500 2035 538
rect 2093 572 2293 610
rect 2093 538 2109 572
rect 2277 538 2293 572
rect 2093 500 2293 538
rect 2351 572 2551 610
rect 2351 538 2367 572
rect 2535 538 2551 572
rect 2351 500 2551 538
rect 2609 572 2809 610
rect 2609 538 2625 572
rect 2793 538 2809 572
rect 2609 500 2809 538
rect 2867 572 3067 610
rect 2867 538 2883 572
rect 3051 538 3067 572
rect 2867 500 3067 538
rect 3125 572 3325 610
rect 3125 538 3141 572
rect 3309 538 3325 572
rect 3125 500 3325 538
rect 3383 572 3583 610
rect 3383 538 3399 572
rect 3567 538 3583 572
rect 3383 500 3583 538
rect 3641 572 3841 610
rect 3641 538 3657 572
rect 3825 538 3841 572
rect 3641 500 3841 538
rect 3899 572 4099 610
rect 3899 538 3915 572
rect 4083 538 4099 572
rect 3899 500 4099 538
rect 4157 572 4357 610
rect 4157 538 4173 572
rect 4341 538 4357 572
rect 4157 500 4357 538
rect 4415 572 4615 610
rect 4415 538 4431 572
rect 4599 538 4615 572
rect 4415 500 4615 538
rect 4673 572 4873 610
rect 4673 538 4689 572
rect 4857 538 4873 572
rect 4673 500 4873 538
rect 4931 572 5131 610
rect 4931 538 4947 572
rect 5115 538 5131 572
rect 4931 500 5131 538
rect 5189 572 5389 610
rect 5189 538 5205 572
rect 5373 538 5389 572
rect 5189 500 5389 538
rect 5447 572 5647 610
rect 5447 538 5463 572
rect 5631 538 5647 572
rect 5447 500 5647 538
rect -5647 -538 -5447 -500
rect -5647 -572 -5631 -538
rect -5463 -572 -5447 -538
rect -5647 -610 -5447 -572
rect -5389 -538 -5189 -500
rect -5389 -572 -5373 -538
rect -5205 -572 -5189 -538
rect -5389 -610 -5189 -572
rect -5131 -538 -4931 -500
rect -5131 -572 -5115 -538
rect -4947 -572 -4931 -538
rect -5131 -610 -4931 -572
rect -4873 -538 -4673 -500
rect -4873 -572 -4857 -538
rect -4689 -572 -4673 -538
rect -4873 -610 -4673 -572
rect -4615 -538 -4415 -500
rect -4615 -572 -4599 -538
rect -4431 -572 -4415 -538
rect -4615 -610 -4415 -572
rect -4357 -538 -4157 -500
rect -4357 -572 -4341 -538
rect -4173 -572 -4157 -538
rect -4357 -610 -4157 -572
rect -4099 -538 -3899 -500
rect -4099 -572 -4083 -538
rect -3915 -572 -3899 -538
rect -4099 -610 -3899 -572
rect -3841 -538 -3641 -500
rect -3841 -572 -3825 -538
rect -3657 -572 -3641 -538
rect -3841 -610 -3641 -572
rect -3583 -538 -3383 -500
rect -3583 -572 -3567 -538
rect -3399 -572 -3383 -538
rect -3583 -610 -3383 -572
rect -3325 -538 -3125 -500
rect -3325 -572 -3309 -538
rect -3141 -572 -3125 -538
rect -3325 -610 -3125 -572
rect -3067 -538 -2867 -500
rect -3067 -572 -3051 -538
rect -2883 -572 -2867 -538
rect -3067 -610 -2867 -572
rect -2809 -538 -2609 -500
rect -2809 -572 -2793 -538
rect -2625 -572 -2609 -538
rect -2809 -610 -2609 -572
rect -2551 -538 -2351 -500
rect -2551 -572 -2535 -538
rect -2367 -572 -2351 -538
rect -2551 -610 -2351 -572
rect -2293 -538 -2093 -500
rect -2293 -572 -2277 -538
rect -2109 -572 -2093 -538
rect -2293 -610 -2093 -572
rect -2035 -538 -1835 -500
rect -2035 -572 -2019 -538
rect -1851 -572 -1835 -538
rect -2035 -610 -1835 -572
rect -1777 -538 -1577 -500
rect -1777 -572 -1761 -538
rect -1593 -572 -1577 -538
rect -1777 -610 -1577 -572
rect -1519 -538 -1319 -500
rect -1519 -572 -1503 -538
rect -1335 -572 -1319 -538
rect -1519 -610 -1319 -572
rect -1261 -538 -1061 -500
rect -1261 -572 -1245 -538
rect -1077 -572 -1061 -538
rect -1261 -610 -1061 -572
rect -1003 -538 -803 -500
rect -1003 -572 -987 -538
rect -819 -572 -803 -538
rect -1003 -610 -803 -572
rect -745 -538 -545 -500
rect -745 -572 -729 -538
rect -561 -572 -545 -538
rect -745 -610 -545 -572
rect -487 -538 -287 -500
rect -487 -572 -471 -538
rect -303 -572 -287 -538
rect -487 -610 -287 -572
rect -229 -538 -29 -500
rect -229 -572 -213 -538
rect -45 -572 -29 -538
rect -229 -610 -29 -572
rect 29 -538 229 -500
rect 29 -572 45 -538
rect 213 -572 229 -538
rect 29 -610 229 -572
rect 287 -538 487 -500
rect 287 -572 303 -538
rect 471 -572 487 -538
rect 287 -610 487 -572
rect 545 -538 745 -500
rect 545 -572 561 -538
rect 729 -572 745 -538
rect 545 -610 745 -572
rect 803 -538 1003 -500
rect 803 -572 819 -538
rect 987 -572 1003 -538
rect 803 -610 1003 -572
rect 1061 -538 1261 -500
rect 1061 -572 1077 -538
rect 1245 -572 1261 -538
rect 1061 -610 1261 -572
rect 1319 -538 1519 -500
rect 1319 -572 1335 -538
rect 1503 -572 1519 -538
rect 1319 -610 1519 -572
rect 1577 -538 1777 -500
rect 1577 -572 1593 -538
rect 1761 -572 1777 -538
rect 1577 -610 1777 -572
rect 1835 -538 2035 -500
rect 1835 -572 1851 -538
rect 2019 -572 2035 -538
rect 1835 -610 2035 -572
rect 2093 -538 2293 -500
rect 2093 -572 2109 -538
rect 2277 -572 2293 -538
rect 2093 -610 2293 -572
rect 2351 -538 2551 -500
rect 2351 -572 2367 -538
rect 2535 -572 2551 -538
rect 2351 -610 2551 -572
rect 2609 -538 2809 -500
rect 2609 -572 2625 -538
rect 2793 -572 2809 -538
rect 2609 -610 2809 -572
rect 2867 -538 3067 -500
rect 2867 -572 2883 -538
rect 3051 -572 3067 -538
rect 2867 -610 3067 -572
rect 3125 -538 3325 -500
rect 3125 -572 3141 -538
rect 3309 -572 3325 -538
rect 3125 -610 3325 -572
rect 3383 -538 3583 -500
rect 3383 -572 3399 -538
rect 3567 -572 3583 -538
rect 3383 -610 3583 -572
rect 3641 -538 3841 -500
rect 3641 -572 3657 -538
rect 3825 -572 3841 -538
rect 3641 -610 3841 -572
rect 3899 -538 4099 -500
rect 3899 -572 3915 -538
rect 4083 -572 4099 -538
rect 3899 -610 4099 -572
rect 4157 -538 4357 -500
rect 4157 -572 4173 -538
rect 4341 -572 4357 -538
rect 4157 -610 4357 -572
rect 4415 -538 4615 -500
rect 4415 -572 4431 -538
rect 4599 -572 4615 -538
rect 4415 -610 4615 -572
rect 4673 -538 4873 -500
rect 4673 -572 4689 -538
rect 4857 -572 4873 -538
rect 4673 -610 4873 -572
rect 4931 -538 5131 -500
rect 4931 -572 4947 -538
rect 5115 -572 5131 -538
rect 4931 -610 5131 -572
rect 5189 -538 5389 -500
rect 5189 -572 5205 -538
rect 5373 -572 5389 -538
rect 5189 -610 5389 -572
rect 5447 -538 5647 -500
rect 5447 -572 5463 -538
rect 5631 -572 5647 -538
rect 5447 -610 5647 -572
rect -5647 -1648 -5447 -1610
rect -5647 -1682 -5631 -1648
rect -5463 -1682 -5447 -1648
rect -5647 -1720 -5447 -1682
rect -5389 -1648 -5189 -1610
rect -5389 -1682 -5373 -1648
rect -5205 -1682 -5189 -1648
rect -5389 -1720 -5189 -1682
rect -5131 -1648 -4931 -1610
rect -5131 -1682 -5115 -1648
rect -4947 -1682 -4931 -1648
rect -5131 -1720 -4931 -1682
rect -4873 -1648 -4673 -1610
rect -4873 -1682 -4857 -1648
rect -4689 -1682 -4673 -1648
rect -4873 -1720 -4673 -1682
rect -4615 -1648 -4415 -1610
rect -4615 -1682 -4599 -1648
rect -4431 -1682 -4415 -1648
rect -4615 -1720 -4415 -1682
rect -4357 -1648 -4157 -1610
rect -4357 -1682 -4341 -1648
rect -4173 -1682 -4157 -1648
rect -4357 -1720 -4157 -1682
rect -4099 -1648 -3899 -1610
rect -4099 -1682 -4083 -1648
rect -3915 -1682 -3899 -1648
rect -4099 -1720 -3899 -1682
rect -3841 -1648 -3641 -1610
rect -3841 -1682 -3825 -1648
rect -3657 -1682 -3641 -1648
rect -3841 -1720 -3641 -1682
rect -3583 -1648 -3383 -1610
rect -3583 -1682 -3567 -1648
rect -3399 -1682 -3383 -1648
rect -3583 -1720 -3383 -1682
rect -3325 -1648 -3125 -1610
rect -3325 -1682 -3309 -1648
rect -3141 -1682 -3125 -1648
rect -3325 -1720 -3125 -1682
rect -3067 -1648 -2867 -1610
rect -3067 -1682 -3051 -1648
rect -2883 -1682 -2867 -1648
rect -3067 -1720 -2867 -1682
rect -2809 -1648 -2609 -1610
rect -2809 -1682 -2793 -1648
rect -2625 -1682 -2609 -1648
rect -2809 -1720 -2609 -1682
rect -2551 -1648 -2351 -1610
rect -2551 -1682 -2535 -1648
rect -2367 -1682 -2351 -1648
rect -2551 -1720 -2351 -1682
rect -2293 -1648 -2093 -1610
rect -2293 -1682 -2277 -1648
rect -2109 -1682 -2093 -1648
rect -2293 -1720 -2093 -1682
rect -2035 -1648 -1835 -1610
rect -2035 -1682 -2019 -1648
rect -1851 -1682 -1835 -1648
rect -2035 -1720 -1835 -1682
rect -1777 -1648 -1577 -1610
rect -1777 -1682 -1761 -1648
rect -1593 -1682 -1577 -1648
rect -1777 -1720 -1577 -1682
rect -1519 -1648 -1319 -1610
rect -1519 -1682 -1503 -1648
rect -1335 -1682 -1319 -1648
rect -1519 -1720 -1319 -1682
rect -1261 -1648 -1061 -1610
rect -1261 -1682 -1245 -1648
rect -1077 -1682 -1061 -1648
rect -1261 -1720 -1061 -1682
rect -1003 -1648 -803 -1610
rect -1003 -1682 -987 -1648
rect -819 -1682 -803 -1648
rect -1003 -1720 -803 -1682
rect -745 -1648 -545 -1610
rect -745 -1682 -729 -1648
rect -561 -1682 -545 -1648
rect -745 -1720 -545 -1682
rect -487 -1648 -287 -1610
rect -487 -1682 -471 -1648
rect -303 -1682 -287 -1648
rect -487 -1720 -287 -1682
rect -229 -1648 -29 -1610
rect -229 -1682 -213 -1648
rect -45 -1682 -29 -1648
rect -229 -1720 -29 -1682
rect 29 -1648 229 -1610
rect 29 -1682 45 -1648
rect 213 -1682 229 -1648
rect 29 -1720 229 -1682
rect 287 -1648 487 -1610
rect 287 -1682 303 -1648
rect 471 -1682 487 -1648
rect 287 -1720 487 -1682
rect 545 -1648 745 -1610
rect 545 -1682 561 -1648
rect 729 -1682 745 -1648
rect 545 -1720 745 -1682
rect 803 -1648 1003 -1610
rect 803 -1682 819 -1648
rect 987 -1682 1003 -1648
rect 803 -1720 1003 -1682
rect 1061 -1648 1261 -1610
rect 1061 -1682 1077 -1648
rect 1245 -1682 1261 -1648
rect 1061 -1720 1261 -1682
rect 1319 -1648 1519 -1610
rect 1319 -1682 1335 -1648
rect 1503 -1682 1519 -1648
rect 1319 -1720 1519 -1682
rect 1577 -1648 1777 -1610
rect 1577 -1682 1593 -1648
rect 1761 -1682 1777 -1648
rect 1577 -1720 1777 -1682
rect 1835 -1648 2035 -1610
rect 1835 -1682 1851 -1648
rect 2019 -1682 2035 -1648
rect 1835 -1720 2035 -1682
rect 2093 -1648 2293 -1610
rect 2093 -1682 2109 -1648
rect 2277 -1682 2293 -1648
rect 2093 -1720 2293 -1682
rect 2351 -1648 2551 -1610
rect 2351 -1682 2367 -1648
rect 2535 -1682 2551 -1648
rect 2351 -1720 2551 -1682
rect 2609 -1648 2809 -1610
rect 2609 -1682 2625 -1648
rect 2793 -1682 2809 -1648
rect 2609 -1720 2809 -1682
rect 2867 -1648 3067 -1610
rect 2867 -1682 2883 -1648
rect 3051 -1682 3067 -1648
rect 2867 -1720 3067 -1682
rect 3125 -1648 3325 -1610
rect 3125 -1682 3141 -1648
rect 3309 -1682 3325 -1648
rect 3125 -1720 3325 -1682
rect 3383 -1648 3583 -1610
rect 3383 -1682 3399 -1648
rect 3567 -1682 3583 -1648
rect 3383 -1720 3583 -1682
rect 3641 -1648 3841 -1610
rect 3641 -1682 3657 -1648
rect 3825 -1682 3841 -1648
rect 3641 -1720 3841 -1682
rect 3899 -1648 4099 -1610
rect 3899 -1682 3915 -1648
rect 4083 -1682 4099 -1648
rect 3899 -1720 4099 -1682
rect 4157 -1648 4357 -1610
rect 4157 -1682 4173 -1648
rect 4341 -1682 4357 -1648
rect 4157 -1720 4357 -1682
rect 4415 -1648 4615 -1610
rect 4415 -1682 4431 -1648
rect 4599 -1682 4615 -1648
rect 4415 -1720 4615 -1682
rect 4673 -1648 4873 -1610
rect 4673 -1682 4689 -1648
rect 4857 -1682 4873 -1648
rect 4673 -1720 4873 -1682
rect 4931 -1648 5131 -1610
rect 4931 -1682 4947 -1648
rect 5115 -1682 5131 -1648
rect 4931 -1720 5131 -1682
rect 5189 -1648 5389 -1610
rect 5189 -1682 5205 -1648
rect 5373 -1682 5389 -1648
rect 5189 -1720 5389 -1682
rect 5447 -1648 5647 -1610
rect 5447 -1682 5463 -1648
rect 5631 -1682 5647 -1648
rect 5447 -1720 5647 -1682
rect -5647 -2758 -5447 -2720
rect -5647 -2792 -5631 -2758
rect -5463 -2792 -5447 -2758
rect -5647 -2808 -5447 -2792
rect -5389 -2758 -5189 -2720
rect -5389 -2792 -5373 -2758
rect -5205 -2792 -5189 -2758
rect -5389 -2808 -5189 -2792
rect -5131 -2758 -4931 -2720
rect -5131 -2792 -5115 -2758
rect -4947 -2792 -4931 -2758
rect -5131 -2808 -4931 -2792
rect -4873 -2758 -4673 -2720
rect -4873 -2792 -4857 -2758
rect -4689 -2792 -4673 -2758
rect -4873 -2808 -4673 -2792
rect -4615 -2758 -4415 -2720
rect -4615 -2792 -4599 -2758
rect -4431 -2792 -4415 -2758
rect -4615 -2808 -4415 -2792
rect -4357 -2758 -4157 -2720
rect -4357 -2792 -4341 -2758
rect -4173 -2792 -4157 -2758
rect -4357 -2808 -4157 -2792
rect -4099 -2758 -3899 -2720
rect -4099 -2792 -4083 -2758
rect -3915 -2792 -3899 -2758
rect -4099 -2808 -3899 -2792
rect -3841 -2758 -3641 -2720
rect -3841 -2792 -3825 -2758
rect -3657 -2792 -3641 -2758
rect -3841 -2808 -3641 -2792
rect -3583 -2758 -3383 -2720
rect -3583 -2792 -3567 -2758
rect -3399 -2792 -3383 -2758
rect -3583 -2808 -3383 -2792
rect -3325 -2758 -3125 -2720
rect -3325 -2792 -3309 -2758
rect -3141 -2792 -3125 -2758
rect -3325 -2808 -3125 -2792
rect -3067 -2758 -2867 -2720
rect -3067 -2792 -3051 -2758
rect -2883 -2792 -2867 -2758
rect -3067 -2808 -2867 -2792
rect -2809 -2758 -2609 -2720
rect -2809 -2792 -2793 -2758
rect -2625 -2792 -2609 -2758
rect -2809 -2808 -2609 -2792
rect -2551 -2758 -2351 -2720
rect -2551 -2792 -2535 -2758
rect -2367 -2792 -2351 -2758
rect -2551 -2808 -2351 -2792
rect -2293 -2758 -2093 -2720
rect -2293 -2792 -2277 -2758
rect -2109 -2792 -2093 -2758
rect -2293 -2808 -2093 -2792
rect -2035 -2758 -1835 -2720
rect -2035 -2792 -2019 -2758
rect -1851 -2792 -1835 -2758
rect -2035 -2808 -1835 -2792
rect -1777 -2758 -1577 -2720
rect -1777 -2792 -1761 -2758
rect -1593 -2792 -1577 -2758
rect -1777 -2808 -1577 -2792
rect -1519 -2758 -1319 -2720
rect -1519 -2792 -1503 -2758
rect -1335 -2792 -1319 -2758
rect -1519 -2808 -1319 -2792
rect -1261 -2758 -1061 -2720
rect -1261 -2792 -1245 -2758
rect -1077 -2792 -1061 -2758
rect -1261 -2808 -1061 -2792
rect -1003 -2758 -803 -2720
rect -1003 -2792 -987 -2758
rect -819 -2792 -803 -2758
rect -1003 -2808 -803 -2792
rect -745 -2758 -545 -2720
rect -745 -2792 -729 -2758
rect -561 -2792 -545 -2758
rect -745 -2808 -545 -2792
rect -487 -2758 -287 -2720
rect -487 -2792 -471 -2758
rect -303 -2792 -287 -2758
rect -487 -2808 -287 -2792
rect -229 -2758 -29 -2720
rect -229 -2792 -213 -2758
rect -45 -2792 -29 -2758
rect -229 -2808 -29 -2792
rect 29 -2758 229 -2720
rect 29 -2792 45 -2758
rect 213 -2792 229 -2758
rect 29 -2808 229 -2792
rect 287 -2758 487 -2720
rect 287 -2792 303 -2758
rect 471 -2792 487 -2758
rect 287 -2808 487 -2792
rect 545 -2758 745 -2720
rect 545 -2792 561 -2758
rect 729 -2792 745 -2758
rect 545 -2808 745 -2792
rect 803 -2758 1003 -2720
rect 803 -2792 819 -2758
rect 987 -2792 1003 -2758
rect 803 -2808 1003 -2792
rect 1061 -2758 1261 -2720
rect 1061 -2792 1077 -2758
rect 1245 -2792 1261 -2758
rect 1061 -2808 1261 -2792
rect 1319 -2758 1519 -2720
rect 1319 -2792 1335 -2758
rect 1503 -2792 1519 -2758
rect 1319 -2808 1519 -2792
rect 1577 -2758 1777 -2720
rect 1577 -2792 1593 -2758
rect 1761 -2792 1777 -2758
rect 1577 -2808 1777 -2792
rect 1835 -2758 2035 -2720
rect 1835 -2792 1851 -2758
rect 2019 -2792 2035 -2758
rect 1835 -2808 2035 -2792
rect 2093 -2758 2293 -2720
rect 2093 -2792 2109 -2758
rect 2277 -2792 2293 -2758
rect 2093 -2808 2293 -2792
rect 2351 -2758 2551 -2720
rect 2351 -2792 2367 -2758
rect 2535 -2792 2551 -2758
rect 2351 -2808 2551 -2792
rect 2609 -2758 2809 -2720
rect 2609 -2792 2625 -2758
rect 2793 -2792 2809 -2758
rect 2609 -2808 2809 -2792
rect 2867 -2758 3067 -2720
rect 2867 -2792 2883 -2758
rect 3051 -2792 3067 -2758
rect 2867 -2808 3067 -2792
rect 3125 -2758 3325 -2720
rect 3125 -2792 3141 -2758
rect 3309 -2792 3325 -2758
rect 3125 -2808 3325 -2792
rect 3383 -2758 3583 -2720
rect 3383 -2792 3399 -2758
rect 3567 -2792 3583 -2758
rect 3383 -2808 3583 -2792
rect 3641 -2758 3841 -2720
rect 3641 -2792 3657 -2758
rect 3825 -2792 3841 -2758
rect 3641 -2808 3841 -2792
rect 3899 -2758 4099 -2720
rect 3899 -2792 3915 -2758
rect 4083 -2792 4099 -2758
rect 3899 -2808 4099 -2792
rect 4157 -2758 4357 -2720
rect 4157 -2792 4173 -2758
rect 4341 -2792 4357 -2758
rect 4157 -2808 4357 -2792
rect 4415 -2758 4615 -2720
rect 4415 -2792 4431 -2758
rect 4599 -2792 4615 -2758
rect 4415 -2808 4615 -2792
rect 4673 -2758 4873 -2720
rect 4673 -2792 4689 -2758
rect 4857 -2792 4873 -2758
rect 4673 -2808 4873 -2792
rect 4931 -2758 5131 -2720
rect 4931 -2792 4947 -2758
rect 5115 -2792 5131 -2758
rect 4931 -2808 5131 -2792
rect 5189 -2758 5389 -2720
rect 5189 -2792 5205 -2758
rect 5373 -2792 5389 -2758
rect 5189 -2808 5389 -2792
rect 5447 -2758 5647 -2720
rect 5447 -2792 5463 -2758
rect 5631 -2792 5647 -2758
rect 5447 -2808 5647 -2792
<< polycont >>
rect -5631 2758 -5463 2792
rect -5373 2758 -5205 2792
rect -5115 2758 -4947 2792
rect -4857 2758 -4689 2792
rect -4599 2758 -4431 2792
rect -4341 2758 -4173 2792
rect -4083 2758 -3915 2792
rect -3825 2758 -3657 2792
rect -3567 2758 -3399 2792
rect -3309 2758 -3141 2792
rect -3051 2758 -2883 2792
rect -2793 2758 -2625 2792
rect -2535 2758 -2367 2792
rect -2277 2758 -2109 2792
rect -2019 2758 -1851 2792
rect -1761 2758 -1593 2792
rect -1503 2758 -1335 2792
rect -1245 2758 -1077 2792
rect -987 2758 -819 2792
rect -729 2758 -561 2792
rect -471 2758 -303 2792
rect -213 2758 -45 2792
rect 45 2758 213 2792
rect 303 2758 471 2792
rect 561 2758 729 2792
rect 819 2758 987 2792
rect 1077 2758 1245 2792
rect 1335 2758 1503 2792
rect 1593 2758 1761 2792
rect 1851 2758 2019 2792
rect 2109 2758 2277 2792
rect 2367 2758 2535 2792
rect 2625 2758 2793 2792
rect 2883 2758 3051 2792
rect 3141 2758 3309 2792
rect 3399 2758 3567 2792
rect 3657 2758 3825 2792
rect 3915 2758 4083 2792
rect 4173 2758 4341 2792
rect 4431 2758 4599 2792
rect 4689 2758 4857 2792
rect 4947 2758 5115 2792
rect 5205 2758 5373 2792
rect 5463 2758 5631 2792
rect -5631 1648 -5463 1682
rect -5373 1648 -5205 1682
rect -5115 1648 -4947 1682
rect -4857 1648 -4689 1682
rect -4599 1648 -4431 1682
rect -4341 1648 -4173 1682
rect -4083 1648 -3915 1682
rect -3825 1648 -3657 1682
rect -3567 1648 -3399 1682
rect -3309 1648 -3141 1682
rect -3051 1648 -2883 1682
rect -2793 1648 -2625 1682
rect -2535 1648 -2367 1682
rect -2277 1648 -2109 1682
rect -2019 1648 -1851 1682
rect -1761 1648 -1593 1682
rect -1503 1648 -1335 1682
rect -1245 1648 -1077 1682
rect -987 1648 -819 1682
rect -729 1648 -561 1682
rect -471 1648 -303 1682
rect -213 1648 -45 1682
rect 45 1648 213 1682
rect 303 1648 471 1682
rect 561 1648 729 1682
rect 819 1648 987 1682
rect 1077 1648 1245 1682
rect 1335 1648 1503 1682
rect 1593 1648 1761 1682
rect 1851 1648 2019 1682
rect 2109 1648 2277 1682
rect 2367 1648 2535 1682
rect 2625 1648 2793 1682
rect 2883 1648 3051 1682
rect 3141 1648 3309 1682
rect 3399 1648 3567 1682
rect 3657 1648 3825 1682
rect 3915 1648 4083 1682
rect 4173 1648 4341 1682
rect 4431 1648 4599 1682
rect 4689 1648 4857 1682
rect 4947 1648 5115 1682
rect 5205 1648 5373 1682
rect 5463 1648 5631 1682
rect -5631 538 -5463 572
rect -5373 538 -5205 572
rect -5115 538 -4947 572
rect -4857 538 -4689 572
rect -4599 538 -4431 572
rect -4341 538 -4173 572
rect -4083 538 -3915 572
rect -3825 538 -3657 572
rect -3567 538 -3399 572
rect -3309 538 -3141 572
rect -3051 538 -2883 572
rect -2793 538 -2625 572
rect -2535 538 -2367 572
rect -2277 538 -2109 572
rect -2019 538 -1851 572
rect -1761 538 -1593 572
rect -1503 538 -1335 572
rect -1245 538 -1077 572
rect -987 538 -819 572
rect -729 538 -561 572
rect -471 538 -303 572
rect -213 538 -45 572
rect 45 538 213 572
rect 303 538 471 572
rect 561 538 729 572
rect 819 538 987 572
rect 1077 538 1245 572
rect 1335 538 1503 572
rect 1593 538 1761 572
rect 1851 538 2019 572
rect 2109 538 2277 572
rect 2367 538 2535 572
rect 2625 538 2793 572
rect 2883 538 3051 572
rect 3141 538 3309 572
rect 3399 538 3567 572
rect 3657 538 3825 572
rect 3915 538 4083 572
rect 4173 538 4341 572
rect 4431 538 4599 572
rect 4689 538 4857 572
rect 4947 538 5115 572
rect 5205 538 5373 572
rect 5463 538 5631 572
rect -5631 -572 -5463 -538
rect -5373 -572 -5205 -538
rect -5115 -572 -4947 -538
rect -4857 -572 -4689 -538
rect -4599 -572 -4431 -538
rect -4341 -572 -4173 -538
rect -4083 -572 -3915 -538
rect -3825 -572 -3657 -538
rect -3567 -572 -3399 -538
rect -3309 -572 -3141 -538
rect -3051 -572 -2883 -538
rect -2793 -572 -2625 -538
rect -2535 -572 -2367 -538
rect -2277 -572 -2109 -538
rect -2019 -572 -1851 -538
rect -1761 -572 -1593 -538
rect -1503 -572 -1335 -538
rect -1245 -572 -1077 -538
rect -987 -572 -819 -538
rect -729 -572 -561 -538
rect -471 -572 -303 -538
rect -213 -572 -45 -538
rect 45 -572 213 -538
rect 303 -572 471 -538
rect 561 -572 729 -538
rect 819 -572 987 -538
rect 1077 -572 1245 -538
rect 1335 -572 1503 -538
rect 1593 -572 1761 -538
rect 1851 -572 2019 -538
rect 2109 -572 2277 -538
rect 2367 -572 2535 -538
rect 2625 -572 2793 -538
rect 2883 -572 3051 -538
rect 3141 -572 3309 -538
rect 3399 -572 3567 -538
rect 3657 -572 3825 -538
rect 3915 -572 4083 -538
rect 4173 -572 4341 -538
rect 4431 -572 4599 -538
rect 4689 -572 4857 -538
rect 4947 -572 5115 -538
rect 5205 -572 5373 -538
rect 5463 -572 5631 -538
rect -5631 -1682 -5463 -1648
rect -5373 -1682 -5205 -1648
rect -5115 -1682 -4947 -1648
rect -4857 -1682 -4689 -1648
rect -4599 -1682 -4431 -1648
rect -4341 -1682 -4173 -1648
rect -4083 -1682 -3915 -1648
rect -3825 -1682 -3657 -1648
rect -3567 -1682 -3399 -1648
rect -3309 -1682 -3141 -1648
rect -3051 -1682 -2883 -1648
rect -2793 -1682 -2625 -1648
rect -2535 -1682 -2367 -1648
rect -2277 -1682 -2109 -1648
rect -2019 -1682 -1851 -1648
rect -1761 -1682 -1593 -1648
rect -1503 -1682 -1335 -1648
rect -1245 -1682 -1077 -1648
rect -987 -1682 -819 -1648
rect -729 -1682 -561 -1648
rect -471 -1682 -303 -1648
rect -213 -1682 -45 -1648
rect 45 -1682 213 -1648
rect 303 -1682 471 -1648
rect 561 -1682 729 -1648
rect 819 -1682 987 -1648
rect 1077 -1682 1245 -1648
rect 1335 -1682 1503 -1648
rect 1593 -1682 1761 -1648
rect 1851 -1682 2019 -1648
rect 2109 -1682 2277 -1648
rect 2367 -1682 2535 -1648
rect 2625 -1682 2793 -1648
rect 2883 -1682 3051 -1648
rect 3141 -1682 3309 -1648
rect 3399 -1682 3567 -1648
rect 3657 -1682 3825 -1648
rect 3915 -1682 4083 -1648
rect 4173 -1682 4341 -1648
rect 4431 -1682 4599 -1648
rect 4689 -1682 4857 -1648
rect 4947 -1682 5115 -1648
rect 5205 -1682 5373 -1648
rect 5463 -1682 5631 -1648
rect -5631 -2792 -5463 -2758
rect -5373 -2792 -5205 -2758
rect -5115 -2792 -4947 -2758
rect -4857 -2792 -4689 -2758
rect -4599 -2792 -4431 -2758
rect -4341 -2792 -4173 -2758
rect -4083 -2792 -3915 -2758
rect -3825 -2792 -3657 -2758
rect -3567 -2792 -3399 -2758
rect -3309 -2792 -3141 -2758
rect -3051 -2792 -2883 -2758
rect -2793 -2792 -2625 -2758
rect -2535 -2792 -2367 -2758
rect -2277 -2792 -2109 -2758
rect -2019 -2792 -1851 -2758
rect -1761 -2792 -1593 -2758
rect -1503 -2792 -1335 -2758
rect -1245 -2792 -1077 -2758
rect -987 -2792 -819 -2758
rect -729 -2792 -561 -2758
rect -471 -2792 -303 -2758
rect -213 -2792 -45 -2758
rect 45 -2792 213 -2758
rect 303 -2792 471 -2758
rect 561 -2792 729 -2758
rect 819 -2792 987 -2758
rect 1077 -2792 1245 -2758
rect 1335 -2792 1503 -2758
rect 1593 -2792 1761 -2758
rect 1851 -2792 2019 -2758
rect 2109 -2792 2277 -2758
rect 2367 -2792 2535 -2758
rect 2625 -2792 2793 -2758
rect 2883 -2792 3051 -2758
rect 3141 -2792 3309 -2758
rect 3399 -2792 3567 -2758
rect 3657 -2792 3825 -2758
rect 3915 -2792 4083 -2758
rect 4173 -2792 4341 -2758
rect 4431 -2792 4599 -2758
rect 4689 -2792 4857 -2758
rect 4947 -2792 5115 -2758
rect 5205 -2792 5373 -2758
rect 5463 -2792 5631 -2758
<< locali >>
rect -5827 2896 -5731 2930
rect 5731 2896 5827 2930
rect -5827 2834 -5793 2896
rect 5793 2834 5827 2896
rect -5647 2758 -5631 2792
rect -5463 2758 -5447 2792
rect -5389 2758 -5373 2792
rect -5205 2758 -5189 2792
rect -5131 2758 -5115 2792
rect -4947 2758 -4931 2792
rect -4873 2758 -4857 2792
rect -4689 2758 -4673 2792
rect -4615 2758 -4599 2792
rect -4431 2758 -4415 2792
rect -4357 2758 -4341 2792
rect -4173 2758 -4157 2792
rect -4099 2758 -4083 2792
rect -3915 2758 -3899 2792
rect -3841 2758 -3825 2792
rect -3657 2758 -3641 2792
rect -3583 2758 -3567 2792
rect -3399 2758 -3383 2792
rect -3325 2758 -3309 2792
rect -3141 2758 -3125 2792
rect -3067 2758 -3051 2792
rect -2883 2758 -2867 2792
rect -2809 2758 -2793 2792
rect -2625 2758 -2609 2792
rect -2551 2758 -2535 2792
rect -2367 2758 -2351 2792
rect -2293 2758 -2277 2792
rect -2109 2758 -2093 2792
rect -2035 2758 -2019 2792
rect -1851 2758 -1835 2792
rect -1777 2758 -1761 2792
rect -1593 2758 -1577 2792
rect -1519 2758 -1503 2792
rect -1335 2758 -1319 2792
rect -1261 2758 -1245 2792
rect -1077 2758 -1061 2792
rect -1003 2758 -987 2792
rect -819 2758 -803 2792
rect -745 2758 -729 2792
rect -561 2758 -545 2792
rect -487 2758 -471 2792
rect -303 2758 -287 2792
rect -229 2758 -213 2792
rect -45 2758 -29 2792
rect 29 2758 45 2792
rect 213 2758 229 2792
rect 287 2758 303 2792
rect 471 2758 487 2792
rect 545 2758 561 2792
rect 729 2758 745 2792
rect 803 2758 819 2792
rect 987 2758 1003 2792
rect 1061 2758 1077 2792
rect 1245 2758 1261 2792
rect 1319 2758 1335 2792
rect 1503 2758 1519 2792
rect 1577 2758 1593 2792
rect 1761 2758 1777 2792
rect 1835 2758 1851 2792
rect 2019 2758 2035 2792
rect 2093 2758 2109 2792
rect 2277 2758 2293 2792
rect 2351 2758 2367 2792
rect 2535 2758 2551 2792
rect 2609 2758 2625 2792
rect 2793 2758 2809 2792
rect 2867 2758 2883 2792
rect 3051 2758 3067 2792
rect 3125 2758 3141 2792
rect 3309 2758 3325 2792
rect 3383 2758 3399 2792
rect 3567 2758 3583 2792
rect 3641 2758 3657 2792
rect 3825 2758 3841 2792
rect 3899 2758 3915 2792
rect 4083 2758 4099 2792
rect 4157 2758 4173 2792
rect 4341 2758 4357 2792
rect 4415 2758 4431 2792
rect 4599 2758 4615 2792
rect 4673 2758 4689 2792
rect 4857 2758 4873 2792
rect 4931 2758 4947 2792
rect 5115 2758 5131 2792
rect 5189 2758 5205 2792
rect 5373 2758 5389 2792
rect 5447 2758 5463 2792
rect 5631 2758 5647 2792
rect -5693 2708 -5659 2724
rect -5693 1716 -5659 1732
rect -5435 2708 -5401 2724
rect -5435 1716 -5401 1732
rect -5177 2708 -5143 2724
rect -5177 1716 -5143 1732
rect -4919 2708 -4885 2724
rect -4919 1716 -4885 1732
rect -4661 2708 -4627 2724
rect -4661 1716 -4627 1732
rect -4403 2708 -4369 2724
rect -4403 1716 -4369 1732
rect -4145 2708 -4111 2724
rect -4145 1716 -4111 1732
rect -3887 2708 -3853 2724
rect -3887 1716 -3853 1732
rect -3629 2708 -3595 2724
rect -3629 1716 -3595 1732
rect -3371 2708 -3337 2724
rect -3371 1716 -3337 1732
rect -3113 2708 -3079 2724
rect -3113 1716 -3079 1732
rect -2855 2708 -2821 2724
rect -2855 1716 -2821 1732
rect -2597 2708 -2563 2724
rect -2597 1716 -2563 1732
rect -2339 2708 -2305 2724
rect -2339 1716 -2305 1732
rect -2081 2708 -2047 2724
rect -2081 1716 -2047 1732
rect -1823 2708 -1789 2724
rect -1823 1716 -1789 1732
rect -1565 2708 -1531 2724
rect -1565 1716 -1531 1732
rect -1307 2708 -1273 2724
rect -1307 1716 -1273 1732
rect -1049 2708 -1015 2724
rect -1049 1716 -1015 1732
rect -791 2708 -757 2724
rect -791 1716 -757 1732
rect -533 2708 -499 2724
rect -533 1716 -499 1732
rect -275 2708 -241 2724
rect -275 1716 -241 1732
rect -17 2708 17 2724
rect -17 1716 17 1732
rect 241 2708 275 2724
rect 241 1716 275 1732
rect 499 2708 533 2724
rect 499 1716 533 1732
rect 757 2708 791 2724
rect 757 1716 791 1732
rect 1015 2708 1049 2724
rect 1015 1716 1049 1732
rect 1273 2708 1307 2724
rect 1273 1716 1307 1732
rect 1531 2708 1565 2724
rect 1531 1716 1565 1732
rect 1789 2708 1823 2724
rect 1789 1716 1823 1732
rect 2047 2708 2081 2724
rect 2047 1716 2081 1732
rect 2305 2708 2339 2724
rect 2305 1716 2339 1732
rect 2563 2708 2597 2724
rect 2563 1716 2597 1732
rect 2821 2708 2855 2724
rect 2821 1716 2855 1732
rect 3079 2708 3113 2724
rect 3079 1716 3113 1732
rect 3337 2708 3371 2724
rect 3337 1716 3371 1732
rect 3595 2708 3629 2724
rect 3595 1716 3629 1732
rect 3853 2708 3887 2724
rect 3853 1716 3887 1732
rect 4111 2708 4145 2724
rect 4111 1716 4145 1732
rect 4369 2708 4403 2724
rect 4369 1716 4403 1732
rect 4627 2708 4661 2724
rect 4627 1716 4661 1732
rect 4885 2708 4919 2724
rect 4885 1716 4919 1732
rect 5143 2708 5177 2724
rect 5143 1716 5177 1732
rect 5401 2708 5435 2724
rect 5401 1716 5435 1732
rect 5659 2708 5693 2724
rect 5659 1716 5693 1732
rect -5647 1648 -5631 1682
rect -5463 1648 -5447 1682
rect -5389 1648 -5373 1682
rect -5205 1648 -5189 1682
rect -5131 1648 -5115 1682
rect -4947 1648 -4931 1682
rect -4873 1648 -4857 1682
rect -4689 1648 -4673 1682
rect -4615 1648 -4599 1682
rect -4431 1648 -4415 1682
rect -4357 1648 -4341 1682
rect -4173 1648 -4157 1682
rect -4099 1648 -4083 1682
rect -3915 1648 -3899 1682
rect -3841 1648 -3825 1682
rect -3657 1648 -3641 1682
rect -3583 1648 -3567 1682
rect -3399 1648 -3383 1682
rect -3325 1648 -3309 1682
rect -3141 1648 -3125 1682
rect -3067 1648 -3051 1682
rect -2883 1648 -2867 1682
rect -2809 1648 -2793 1682
rect -2625 1648 -2609 1682
rect -2551 1648 -2535 1682
rect -2367 1648 -2351 1682
rect -2293 1648 -2277 1682
rect -2109 1648 -2093 1682
rect -2035 1648 -2019 1682
rect -1851 1648 -1835 1682
rect -1777 1648 -1761 1682
rect -1593 1648 -1577 1682
rect -1519 1648 -1503 1682
rect -1335 1648 -1319 1682
rect -1261 1648 -1245 1682
rect -1077 1648 -1061 1682
rect -1003 1648 -987 1682
rect -819 1648 -803 1682
rect -745 1648 -729 1682
rect -561 1648 -545 1682
rect -487 1648 -471 1682
rect -303 1648 -287 1682
rect -229 1648 -213 1682
rect -45 1648 -29 1682
rect 29 1648 45 1682
rect 213 1648 229 1682
rect 287 1648 303 1682
rect 471 1648 487 1682
rect 545 1648 561 1682
rect 729 1648 745 1682
rect 803 1648 819 1682
rect 987 1648 1003 1682
rect 1061 1648 1077 1682
rect 1245 1648 1261 1682
rect 1319 1648 1335 1682
rect 1503 1648 1519 1682
rect 1577 1648 1593 1682
rect 1761 1648 1777 1682
rect 1835 1648 1851 1682
rect 2019 1648 2035 1682
rect 2093 1648 2109 1682
rect 2277 1648 2293 1682
rect 2351 1648 2367 1682
rect 2535 1648 2551 1682
rect 2609 1648 2625 1682
rect 2793 1648 2809 1682
rect 2867 1648 2883 1682
rect 3051 1648 3067 1682
rect 3125 1648 3141 1682
rect 3309 1648 3325 1682
rect 3383 1648 3399 1682
rect 3567 1648 3583 1682
rect 3641 1648 3657 1682
rect 3825 1648 3841 1682
rect 3899 1648 3915 1682
rect 4083 1648 4099 1682
rect 4157 1648 4173 1682
rect 4341 1648 4357 1682
rect 4415 1648 4431 1682
rect 4599 1648 4615 1682
rect 4673 1648 4689 1682
rect 4857 1648 4873 1682
rect 4931 1648 4947 1682
rect 5115 1648 5131 1682
rect 5189 1648 5205 1682
rect 5373 1648 5389 1682
rect 5447 1648 5463 1682
rect 5631 1648 5647 1682
rect -5693 1598 -5659 1614
rect -5693 606 -5659 622
rect -5435 1598 -5401 1614
rect -5435 606 -5401 622
rect -5177 1598 -5143 1614
rect -5177 606 -5143 622
rect -4919 1598 -4885 1614
rect -4919 606 -4885 622
rect -4661 1598 -4627 1614
rect -4661 606 -4627 622
rect -4403 1598 -4369 1614
rect -4403 606 -4369 622
rect -4145 1598 -4111 1614
rect -4145 606 -4111 622
rect -3887 1598 -3853 1614
rect -3887 606 -3853 622
rect -3629 1598 -3595 1614
rect -3629 606 -3595 622
rect -3371 1598 -3337 1614
rect -3371 606 -3337 622
rect -3113 1598 -3079 1614
rect -3113 606 -3079 622
rect -2855 1598 -2821 1614
rect -2855 606 -2821 622
rect -2597 1598 -2563 1614
rect -2597 606 -2563 622
rect -2339 1598 -2305 1614
rect -2339 606 -2305 622
rect -2081 1598 -2047 1614
rect -2081 606 -2047 622
rect -1823 1598 -1789 1614
rect -1823 606 -1789 622
rect -1565 1598 -1531 1614
rect -1565 606 -1531 622
rect -1307 1598 -1273 1614
rect -1307 606 -1273 622
rect -1049 1598 -1015 1614
rect -1049 606 -1015 622
rect -791 1598 -757 1614
rect -791 606 -757 622
rect -533 1598 -499 1614
rect -533 606 -499 622
rect -275 1598 -241 1614
rect -275 606 -241 622
rect -17 1598 17 1614
rect -17 606 17 622
rect 241 1598 275 1614
rect 241 606 275 622
rect 499 1598 533 1614
rect 499 606 533 622
rect 757 1598 791 1614
rect 757 606 791 622
rect 1015 1598 1049 1614
rect 1015 606 1049 622
rect 1273 1598 1307 1614
rect 1273 606 1307 622
rect 1531 1598 1565 1614
rect 1531 606 1565 622
rect 1789 1598 1823 1614
rect 1789 606 1823 622
rect 2047 1598 2081 1614
rect 2047 606 2081 622
rect 2305 1598 2339 1614
rect 2305 606 2339 622
rect 2563 1598 2597 1614
rect 2563 606 2597 622
rect 2821 1598 2855 1614
rect 2821 606 2855 622
rect 3079 1598 3113 1614
rect 3079 606 3113 622
rect 3337 1598 3371 1614
rect 3337 606 3371 622
rect 3595 1598 3629 1614
rect 3595 606 3629 622
rect 3853 1598 3887 1614
rect 3853 606 3887 622
rect 4111 1598 4145 1614
rect 4111 606 4145 622
rect 4369 1598 4403 1614
rect 4369 606 4403 622
rect 4627 1598 4661 1614
rect 4627 606 4661 622
rect 4885 1598 4919 1614
rect 4885 606 4919 622
rect 5143 1598 5177 1614
rect 5143 606 5177 622
rect 5401 1598 5435 1614
rect 5401 606 5435 622
rect 5659 1598 5693 1614
rect 5659 606 5693 622
rect -5647 538 -5631 572
rect -5463 538 -5447 572
rect -5389 538 -5373 572
rect -5205 538 -5189 572
rect -5131 538 -5115 572
rect -4947 538 -4931 572
rect -4873 538 -4857 572
rect -4689 538 -4673 572
rect -4615 538 -4599 572
rect -4431 538 -4415 572
rect -4357 538 -4341 572
rect -4173 538 -4157 572
rect -4099 538 -4083 572
rect -3915 538 -3899 572
rect -3841 538 -3825 572
rect -3657 538 -3641 572
rect -3583 538 -3567 572
rect -3399 538 -3383 572
rect -3325 538 -3309 572
rect -3141 538 -3125 572
rect -3067 538 -3051 572
rect -2883 538 -2867 572
rect -2809 538 -2793 572
rect -2625 538 -2609 572
rect -2551 538 -2535 572
rect -2367 538 -2351 572
rect -2293 538 -2277 572
rect -2109 538 -2093 572
rect -2035 538 -2019 572
rect -1851 538 -1835 572
rect -1777 538 -1761 572
rect -1593 538 -1577 572
rect -1519 538 -1503 572
rect -1335 538 -1319 572
rect -1261 538 -1245 572
rect -1077 538 -1061 572
rect -1003 538 -987 572
rect -819 538 -803 572
rect -745 538 -729 572
rect -561 538 -545 572
rect -487 538 -471 572
rect -303 538 -287 572
rect -229 538 -213 572
rect -45 538 -29 572
rect 29 538 45 572
rect 213 538 229 572
rect 287 538 303 572
rect 471 538 487 572
rect 545 538 561 572
rect 729 538 745 572
rect 803 538 819 572
rect 987 538 1003 572
rect 1061 538 1077 572
rect 1245 538 1261 572
rect 1319 538 1335 572
rect 1503 538 1519 572
rect 1577 538 1593 572
rect 1761 538 1777 572
rect 1835 538 1851 572
rect 2019 538 2035 572
rect 2093 538 2109 572
rect 2277 538 2293 572
rect 2351 538 2367 572
rect 2535 538 2551 572
rect 2609 538 2625 572
rect 2793 538 2809 572
rect 2867 538 2883 572
rect 3051 538 3067 572
rect 3125 538 3141 572
rect 3309 538 3325 572
rect 3383 538 3399 572
rect 3567 538 3583 572
rect 3641 538 3657 572
rect 3825 538 3841 572
rect 3899 538 3915 572
rect 4083 538 4099 572
rect 4157 538 4173 572
rect 4341 538 4357 572
rect 4415 538 4431 572
rect 4599 538 4615 572
rect 4673 538 4689 572
rect 4857 538 4873 572
rect 4931 538 4947 572
rect 5115 538 5131 572
rect 5189 538 5205 572
rect 5373 538 5389 572
rect 5447 538 5463 572
rect 5631 538 5647 572
rect -5693 488 -5659 504
rect -5693 -504 -5659 -488
rect -5435 488 -5401 504
rect -5435 -504 -5401 -488
rect -5177 488 -5143 504
rect -5177 -504 -5143 -488
rect -4919 488 -4885 504
rect -4919 -504 -4885 -488
rect -4661 488 -4627 504
rect -4661 -504 -4627 -488
rect -4403 488 -4369 504
rect -4403 -504 -4369 -488
rect -4145 488 -4111 504
rect -4145 -504 -4111 -488
rect -3887 488 -3853 504
rect -3887 -504 -3853 -488
rect -3629 488 -3595 504
rect -3629 -504 -3595 -488
rect -3371 488 -3337 504
rect -3371 -504 -3337 -488
rect -3113 488 -3079 504
rect -3113 -504 -3079 -488
rect -2855 488 -2821 504
rect -2855 -504 -2821 -488
rect -2597 488 -2563 504
rect -2597 -504 -2563 -488
rect -2339 488 -2305 504
rect -2339 -504 -2305 -488
rect -2081 488 -2047 504
rect -2081 -504 -2047 -488
rect -1823 488 -1789 504
rect -1823 -504 -1789 -488
rect -1565 488 -1531 504
rect -1565 -504 -1531 -488
rect -1307 488 -1273 504
rect -1307 -504 -1273 -488
rect -1049 488 -1015 504
rect -1049 -504 -1015 -488
rect -791 488 -757 504
rect -791 -504 -757 -488
rect -533 488 -499 504
rect -533 -504 -499 -488
rect -275 488 -241 504
rect -275 -504 -241 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 241 488 275 504
rect 241 -504 275 -488
rect 499 488 533 504
rect 499 -504 533 -488
rect 757 488 791 504
rect 757 -504 791 -488
rect 1015 488 1049 504
rect 1015 -504 1049 -488
rect 1273 488 1307 504
rect 1273 -504 1307 -488
rect 1531 488 1565 504
rect 1531 -504 1565 -488
rect 1789 488 1823 504
rect 1789 -504 1823 -488
rect 2047 488 2081 504
rect 2047 -504 2081 -488
rect 2305 488 2339 504
rect 2305 -504 2339 -488
rect 2563 488 2597 504
rect 2563 -504 2597 -488
rect 2821 488 2855 504
rect 2821 -504 2855 -488
rect 3079 488 3113 504
rect 3079 -504 3113 -488
rect 3337 488 3371 504
rect 3337 -504 3371 -488
rect 3595 488 3629 504
rect 3595 -504 3629 -488
rect 3853 488 3887 504
rect 3853 -504 3887 -488
rect 4111 488 4145 504
rect 4111 -504 4145 -488
rect 4369 488 4403 504
rect 4369 -504 4403 -488
rect 4627 488 4661 504
rect 4627 -504 4661 -488
rect 4885 488 4919 504
rect 4885 -504 4919 -488
rect 5143 488 5177 504
rect 5143 -504 5177 -488
rect 5401 488 5435 504
rect 5401 -504 5435 -488
rect 5659 488 5693 504
rect 5659 -504 5693 -488
rect -5647 -572 -5631 -538
rect -5463 -572 -5447 -538
rect -5389 -572 -5373 -538
rect -5205 -572 -5189 -538
rect -5131 -572 -5115 -538
rect -4947 -572 -4931 -538
rect -4873 -572 -4857 -538
rect -4689 -572 -4673 -538
rect -4615 -572 -4599 -538
rect -4431 -572 -4415 -538
rect -4357 -572 -4341 -538
rect -4173 -572 -4157 -538
rect -4099 -572 -4083 -538
rect -3915 -572 -3899 -538
rect -3841 -572 -3825 -538
rect -3657 -572 -3641 -538
rect -3583 -572 -3567 -538
rect -3399 -572 -3383 -538
rect -3325 -572 -3309 -538
rect -3141 -572 -3125 -538
rect -3067 -572 -3051 -538
rect -2883 -572 -2867 -538
rect -2809 -572 -2793 -538
rect -2625 -572 -2609 -538
rect -2551 -572 -2535 -538
rect -2367 -572 -2351 -538
rect -2293 -572 -2277 -538
rect -2109 -572 -2093 -538
rect -2035 -572 -2019 -538
rect -1851 -572 -1835 -538
rect -1777 -572 -1761 -538
rect -1593 -572 -1577 -538
rect -1519 -572 -1503 -538
rect -1335 -572 -1319 -538
rect -1261 -572 -1245 -538
rect -1077 -572 -1061 -538
rect -1003 -572 -987 -538
rect -819 -572 -803 -538
rect -745 -572 -729 -538
rect -561 -572 -545 -538
rect -487 -572 -471 -538
rect -303 -572 -287 -538
rect -229 -572 -213 -538
rect -45 -572 -29 -538
rect 29 -572 45 -538
rect 213 -572 229 -538
rect 287 -572 303 -538
rect 471 -572 487 -538
rect 545 -572 561 -538
rect 729 -572 745 -538
rect 803 -572 819 -538
rect 987 -572 1003 -538
rect 1061 -572 1077 -538
rect 1245 -572 1261 -538
rect 1319 -572 1335 -538
rect 1503 -572 1519 -538
rect 1577 -572 1593 -538
rect 1761 -572 1777 -538
rect 1835 -572 1851 -538
rect 2019 -572 2035 -538
rect 2093 -572 2109 -538
rect 2277 -572 2293 -538
rect 2351 -572 2367 -538
rect 2535 -572 2551 -538
rect 2609 -572 2625 -538
rect 2793 -572 2809 -538
rect 2867 -572 2883 -538
rect 3051 -572 3067 -538
rect 3125 -572 3141 -538
rect 3309 -572 3325 -538
rect 3383 -572 3399 -538
rect 3567 -572 3583 -538
rect 3641 -572 3657 -538
rect 3825 -572 3841 -538
rect 3899 -572 3915 -538
rect 4083 -572 4099 -538
rect 4157 -572 4173 -538
rect 4341 -572 4357 -538
rect 4415 -572 4431 -538
rect 4599 -572 4615 -538
rect 4673 -572 4689 -538
rect 4857 -572 4873 -538
rect 4931 -572 4947 -538
rect 5115 -572 5131 -538
rect 5189 -572 5205 -538
rect 5373 -572 5389 -538
rect 5447 -572 5463 -538
rect 5631 -572 5647 -538
rect -5693 -622 -5659 -606
rect -5693 -1614 -5659 -1598
rect -5435 -622 -5401 -606
rect -5435 -1614 -5401 -1598
rect -5177 -622 -5143 -606
rect -5177 -1614 -5143 -1598
rect -4919 -622 -4885 -606
rect -4919 -1614 -4885 -1598
rect -4661 -622 -4627 -606
rect -4661 -1614 -4627 -1598
rect -4403 -622 -4369 -606
rect -4403 -1614 -4369 -1598
rect -4145 -622 -4111 -606
rect -4145 -1614 -4111 -1598
rect -3887 -622 -3853 -606
rect -3887 -1614 -3853 -1598
rect -3629 -622 -3595 -606
rect -3629 -1614 -3595 -1598
rect -3371 -622 -3337 -606
rect -3371 -1614 -3337 -1598
rect -3113 -622 -3079 -606
rect -3113 -1614 -3079 -1598
rect -2855 -622 -2821 -606
rect -2855 -1614 -2821 -1598
rect -2597 -622 -2563 -606
rect -2597 -1614 -2563 -1598
rect -2339 -622 -2305 -606
rect -2339 -1614 -2305 -1598
rect -2081 -622 -2047 -606
rect -2081 -1614 -2047 -1598
rect -1823 -622 -1789 -606
rect -1823 -1614 -1789 -1598
rect -1565 -622 -1531 -606
rect -1565 -1614 -1531 -1598
rect -1307 -622 -1273 -606
rect -1307 -1614 -1273 -1598
rect -1049 -622 -1015 -606
rect -1049 -1614 -1015 -1598
rect -791 -622 -757 -606
rect -791 -1614 -757 -1598
rect -533 -622 -499 -606
rect -533 -1614 -499 -1598
rect -275 -622 -241 -606
rect -275 -1614 -241 -1598
rect -17 -622 17 -606
rect -17 -1614 17 -1598
rect 241 -622 275 -606
rect 241 -1614 275 -1598
rect 499 -622 533 -606
rect 499 -1614 533 -1598
rect 757 -622 791 -606
rect 757 -1614 791 -1598
rect 1015 -622 1049 -606
rect 1015 -1614 1049 -1598
rect 1273 -622 1307 -606
rect 1273 -1614 1307 -1598
rect 1531 -622 1565 -606
rect 1531 -1614 1565 -1598
rect 1789 -622 1823 -606
rect 1789 -1614 1823 -1598
rect 2047 -622 2081 -606
rect 2047 -1614 2081 -1598
rect 2305 -622 2339 -606
rect 2305 -1614 2339 -1598
rect 2563 -622 2597 -606
rect 2563 -1614 2597 -1598
rect 2821 -622 2855 -606
rect 2821 -1614 2855 -1598
rect 3079 -622 3113 -606
rect 3079 -1614 3113 -1598
rect 3337 -622 3371 -606
rect 3337 -1614 3371 -1598
rect 3595 -622 3629 -606
rect 3595 -1614 3629 -1598
rect 3853 -622 3887 -606
rect 3853 -1614 3887 -1598
rect 4111 -622 4145 -606
rect 4111 -1614 4145 -1598
rect 4369 -622 4403 -606
rect 4369 -1614 4403 -1598
rect 4627 -622 4661 -606
rect 4627 -1614 4661 -1598
rect 4885 -622 4919 -606
rect 4885 -1614 4919 -1598
rect 5143 -622 5177 -606
rect 5143 -1614 5177 -1598
rect 5401 -622 5435 -606
rect 5401 -1614 5435 -1598
rect 5659 -622 5693 -606
rect 5659 -1614 5693 -1598
rect -5647 -1682 -5631 -1648
rect -5463 -1682 -5447 -1648
rect -5389 -1682 -5373 -1648
rect -5205 -1682 -5189 -1648
rect -5131 -1682 -5115 -1648
rect -4947 -1682 -4931 -1648
rect -4873 -1682 -4857 -1648
rect -4689 -1682 -4673 -1648
rect -4615 -1682 -4599 -1648
rect -4431 -1682 -4415 -1648
rect -4357 -1682 -4341 -1648
rect -4173 -1682 -4157 -1648
rect -4099 -1682 -4083 -1648
rect -3915 -1682 -3899 -1648
rect -3841 -1682 -3825 -1648
rect -3657 -1682 -3641 -1648
rect -3583 -1682 -3567 -1648
rect -3399 -1682 -3383 -1648
rect -3325 -1682 -3309 -1648
rect -3141 -1682 -3125 -1648
rect -3067 -1682 -3051 -1648
rect -2883 -1682 -2867 -1648
rect -2809 -1682 -2793 -1648
rect -2625 -1682 -2609 -1648
rect -2551 -1682 -2535 -1648
rect -2367 -1682 -2351 -1648
rect -2293 -1682 -2277 -1648
rect -2109 -1682 -2093 -1648
rect -2035 -1682 -2019 -1648
rect -1851 -1682 -1835 -1648
rect -1777 -1682 -1761 -1648
rect -1593 -1682 -1577 -1648
rect -1519 -1682 -1503 -1648
rect -1335 -1682 -1319 -1648
rect -1261 -1682 -1245 -1648
rect -1077 -1682 -1061 -1648
rect -1003 -1682 -987 -1648
rect -819 -1682 -803 -1648
rect -745 -1682 -729 -1648
rect -561 -1682 -545 -1648
rect -487 -1682 -471 -1648
rect -303 -1682 -287 -1648
rect -229 -1682 -213 -1648
rect -45 -1682 -29 -1648
rect 29 -1682 45 -1648
rect 213 -1682 229 -1648
rect 287 -1682 303 -1648
rect 471 -1682 487 -1648
rect 545 -1682 561 -1648
rect 729 -1682 745 -1648
rect 803 -1682 819 -1648
rect 987 -1682 1003 -1648
rect 1061 -1682 1077 -1648
rect 1245 -1682 1261 -1648
rect 1319 -1682 1335 -1648
rect 1503 -1682 1519 -1648
rect 1577 -1682 1593 -1648
rect 1761 -1682 1777 -1648
rect 1835 -1682 1851 -1648
rect 2019 -1682 2035 -1648
rect 2093 -1682 2109 -1648
rect 2277 -1682 2293 -1648
rect 2351 -1682 2367 -1648
rect 2535 -1682 2551 -1648
rect 2609 -1682 2625 -1648
rect 2793 -1682 2809 -1648
rect 2867 -1682 2883 -1648
rect 3051 -1682 3067 -1648
rect 3125 -1682 3141 -1648
rect 3309 -1682 3325 -1648
rect 3383 -1682 3399 -1648
rect 3567 -1682 3583 -1648
rect 3641 -1682 3657 -1648
rect 3825 -1682 3841 -1648
rect 3899 -1682 3915 -1648
rect 4083 -1682 4099 -1648
rect 4157 -1682 4173 -1648
rect 4341 -1682 4357 -1648
rect 4415 -1682 4431 -1648
rect 4599 -1682 4615 -1648
rect 4673 -1682 4689 -1648
rect 4857 -1682 4873 -1648
rect 4931 -1682 4947 -1648
rect 5115 -1682 5131 -1648
rect 5189 -1682 5205 -1648
rect 5373 -1682 5389 -1648
rect 5447 -1682 5463 -1648
rect 5631 -1682 5647 -1648
rect -5693 -1732 -5659 -1716
rect -5693 -2724 -5659 -2708
rect -5435 -1732 -5401 -1716
rect -5435 -2724 -5401 -2708
rect -5177 -1732 -5143 -1716
rect -5177 -2724 -5143 -2708
rect -4919 -1732 -4885 -1716
rect -4919 -2724 -4885 -2708
rect -4661 -1732 -4627 -1716
rect -4661 -2724 -4627 -2708
rect -4403 -1732 -4369 -1716
rect -4403 -2724 -4369 -2708
rect -4145 -1732 -4111 -1716
rect -4145 -2724 -4111 -2708
rect -3887 -1732 -3853 -1716
rect -3887 -2724 -3853 -2708
rect -3629 -1732 -3595 -1716
rect -3629 -2724 -3595 -2708
rect -3371 -1732 -3337 -1716
rect -3371 -2724 -3337 -2708
rect -3113 -1732 -3079 -1716
rect -3113 -2724 -3079 -2708
rect -2855 -1732 -2821 -1716
rect -2855 -2724 -2821 -2708
rect -2597 -1732 -2563 -1716
rect -2597 -2724 -2563 -2708
rect -2339 -1732 -2305 -1716
rect -2339 -2724 -2305 -2708
rect -2081 -1732 -2047 -1716
rect -2081 -2724 -2047 -2708
rect -1823 -1732 -1789 -1716
rect -1823 -2724 -1789 -2708
rect -1565 -1732 -1531 -1716
rect -1565 -2724 -1531 -2708
rect -1307 -1732 -1273 -1716
rect -1307 -2724 -1273 -2708
rect -1049 -1732 -1015 -1716
rect -1049 -2724 -1015 -2708
rect -791 -1732 -757 -1716
rect -791 -2724 -757 -2708
rect -533 -1732 -499 -1716
rect -533 -2724 -499 -2708
rect -275 -1732 -241 -1716
rect -275 -2724 -241 -2708
rect -17 -1732 17 -1716
rect -17 -2724 17 -2708
rect 241 -1732 275 -1716
rect 241 -2724 275 -2708
rect 499 -1732 533 -1716
rect 499 -2724 533 -2708
rect 757 -1732 791 -1716
rect 757 -2724 791 -2708
rect 1015 -1732 1049 -1716
rect 1015 -2724 1049 -2708
rect 1273 -1732 1307 -1716
rect 1273 -2724 1307 -2708
rect 1531 -1732 1565 -1716
rect 1531 -2724 1565 -2708
rect 1789 -1732 1823 -1716
rect 1789 -2724 1823 -2708
rect 2047 -1732 2081 -1716
rect 2047 -2724 2081 -2708
rect 2305 -1732 2339 -1716
rect 2305 -2724 2339 -2708
rect 2563 -1732 2597 -1716
rect 2563 -2724 2597 -2708
rect 2821 -1732 2855 -1716
rect 2821 -2724 2855 -2708
rect 3079 -1732 3113 -1716
rect 3079 -2724 3113 -2708
rect 3337 -1732 3371 -1716
rect 3337 -2724 3371 -2708
rect 3595 -1732 3629 -1716
rect 3595 -2724 3629 -2708
rect 3853 -1732 3887 -1716
rect 3853 -2724 3887 -2708
rect 4111 -1732 4145 -1716
rect 4111 -2724 4145 -2708
rect 4369 -1732 4403 -1716
rect 4369 -2724 4403 -2708
rect 4627 -1732 4661 -1716
rect 4627 -2724 4661 -2708
rect 4885 -1732 4919 -1716
rect 4885 -2724 4919 -2708
rect 5143 -1732 5177 -1716
rect 5143 -2724 5177 -2708
rect 5401 -1732 5435 -1716
rect 5401 -2724 5435 -2708
rect 5659 -1732 5693 -1716
rect 5659 -2724 5693 -2708
rect -5647 -2792 -5631 -2758
rect -5463 -2792 -5447 -2758
rect -5389 -2792 -5373 -2758
rect -5205 -2792 -5189 -2758
rect -5131 -2792 -5115 -2758
rect -4947 -2792 -4931 -2758
rect -4873 -2792 -4857 -2758
rect -4689 -2792 -4673 -2758
rect -4615 -2792 -4599 -2758
rect -4431 -2792 -4415 -2758
rect -4357 -2792 -4341 -2758
rect -4173 -2792 -4157 -2758
rect -4099 -2792 -4083 -2758
rect -3915 -2792 -3899 -2758
rect -3841 -2792 -3825 -2758
rect -3657 -2792 -3641 -2758
rect -3583 -2792 -3567 -2758
rect -3399 -2792 -3383 -2758
rect -3325 -2792 -3309 -2758
rect -3141 -2792 -3125 -2758
rect -3067 -2792 -3051 -2758
rect -2883 -2792 -2867 -2758
rect -2809 -2792 -2793 -2758
rect -2625 -2792 -2609 -2758
rect -2551 -2792 -2535 -2758
rect -2367 -2792 -2351 -2758
rect -2293 -2792 -2277 -2758
rect -2109 -2792 -2093 -2758
rect -2035 -2792 -2019 -2758
rect -1851 -2792 -1835 -2758
rect -1777 -2792 -1761 -2758
rect -1593 -2792 -1577 -2758
rect -1519 -2792 -1503 -2758
rect -1335 -2792 -1319 -2758
rect -1261 -2792 -1245 -2758
rect -1077 -2792 -1061 -2758
rect -1003 -2792 -987 -2758
rect -819 -2792 -803 -2758
rect -745 -2792 -729 -2758
rect -561 -2792 -545 -2758
rect -487 -2792 -471 -2758
rect -303 -2792 -287 -2758
rect -229 -2792 -213 -2758
rect -45 -2792 -29 -2758
rect 29 -2792 45 -2758
rect 213 -2792 229 -2758
rect 287 -2792 303 -2758
rect 471 -2792 487 -2758
rect 545 -2792 561 -2758
rect 729 -2792 745 -2758
rect 803 -2792 819 -2758
rect 987 -2792 1003 -2758
rect 1061 -2792 1077 -2758
rect 1245 -2792 1261 -2758
rect 1319 -2792 1335 -2758
rect 1503 -2792 1519 -2758
rect 1577 -2792 1593 -2758
rect 1761 -2792 1777 -2758
rect 1835 -2792 1851 -2758
rect 2019 -2792 2035 -2758
rect 2093 -2792 2109 -2758
rect 2277 -2792 2293 -2758
rect 2351 -2792 2367 -2758
rect 2535 -2792 2551 -2758
rect 2609 -2792 2625 -2758
rect 2793 -2792 2809 -2758
rect 2867 -2792 2883 -2758
rect 3051 -2792 3067 -2758
rect 3125 -2792 3141 -2758
rect 3309 -2792 3325 -2758
rect 3383 -2792 3399 -2758
rect 3567 -2792 3583 -2758
rect 3641 -2792 3657 -2758
rect 3825 -2792 3841 -2758
rect 3899 -2792 3915 -2758
rect 4083 -2792 4099 -2758
rect 4157 -2792 4173 -2758
rect 4341 -2792 4357 -2758
rect 4415 -2792 4431 -2758
rect 4599 -2792 4615 -2758
rect 4673 -2792 4689 -2758
rect 4857 -2792 4873 -2758
rect 4931 -2792 4947 -2758
rect 5115 -2792 5131 -2758
rect 5189 -2792 5205 -2758
rect 5373 -2792 5389 -2758
rect 5447 -2792 5463 -2758
rect 5631 -2792 5647 -2758
rect -5827 -2896 -5793 -2834
rect 5793 -2896 5827 -2834
rect -5827 -2930 -5731 -2896
rect 5731 -2930 5827 -2896
<< viali >>
rect -5631 2758 -5463 2792
rect -5373 2758 -5205 2792
rect -5115 2758 -4947 2792
rect -4857 2758 -4689 2792
rect -4599 2758 -4431 2792
rect -4341 2758 -4173 2792
rect -4083 2758 -3915 2792
rect -3825 2758 -3657 2792
rect -3567 2758 -3399 2792
rect -3309 2758 -3141 2792
rect -3051 2758 -2883 2792
rect -2793 2758 -2625 2792
rect -2535 2758 -2367 2792
rect -2277 2758 -2109 2792
rect -2019 2758 -1851 2792
rect -1761 2758 -1593 2792
rect -1503 2758 -1335 2792
rect -1245 2758 -1077 2792
rect -987 2758 -819 2792
rect -729 2758 -561 2792
rect -471 2758 -303 2792
rect -213 2758 -45 2792
rect 45 2758 213 2792
rect 303 2758 471 2792
rect 561 2758 729 2792
rect 819 2758 987 2792
rect 1077 2758 1245 2792
rect 1335 2758 1503 2792
rect 1593 2758 1761 2792
rect 1851 2758 2019 2792
rect 2109 2758 2277 2792
rect 2367 2758 2535 2792
rect 2625 2758 2793 2792
rect 2883 2758 3051 2792
rect 3141 2758 3309 2792
rect 3399 2758 3567 2792
rect 3657 2758 3825 2792
rect 3915 2758 4083 2792
rect 4173 2758 4341 2792
rect 4431 2758 4599 2792
rect 4689 2758 4857 2792
rect 4947 2758 5115 2792
rect 5205 2758 5373 2792
rect 5463 2758 5631 2792
rect -5693 1732 -5659 2708
rect -5435 1732 -5401 2708
rect -5177 1732 -5143 2708
rect -4919 1732 -4885 2708
rect -4661 1732 -4627 2708
rect -4403 1732 -4369 2708
rect -4145 1732 -4111 2708
rect -3887 1732 -3853 2708
rect -3629 1732 -3595 2708
rect -3371 1732 -3337 2708
rect -3113 1732 -3079 2708
rect -2855 1732 -2821 2708
rect -2597 1732 -2563 2708
rect -2339 1732 -2305 2708
rect -2081 1732 -2047 2708
rect -1823 1732 -1789 2708
rect -1565 1732 -1531 2708
rect -1307 1732 -1273 2708
rect -1049 1732 -1015 2708
rect -791 1732 -757 2708
rect -533 1732 -499 2708
rect -275 1732 -241 2708
rect -17 1732 17 2708
rect 241 1732 275 2708
rect 499 1732 533 2708
rect 757 1732 791 2708
rect 1015 1732 1049 2708
rect 1273 1732 1307 2708
rect 1531 1732 1565 2708
rect 1789 1732 1823 2708
rect 2047 1732 2081 2708
rect 2305 1732 2339 2708
rect 2563 1732 2597 2708
rect 2821 1732 2855 2708
rect 3079 1732 3113 2708
rect 3337 1732 3371 2708
rect 3595 1732 3629 2708
rect 3853 1732 3887 2708
rect 4111 1732 4145 2708
rect 4369 1732 4403 2708
rect 4627 1732 4661 2708
rect 4885 1732 4919 2708
rect 5143 1732 5177 2708
rect 5401 1732 5435 2708
rect 5659 1732 5693 2708
rect -5631 1648 -5463 1682
rect -5373 1648 -5205 1682
rect -5115 1648 -4947 1682
rect -4857 1648 -4689 1682
rect -4599 1648 -4431 1682
rect -4341 1648 -4173 1682
rect -4083 1648 -3915 1682
rect -3825 1648 -3657 1682
rect -3567 1648 -3399 1682
rect -3309 1648 -3141 1682
rect -3051 1648 -2883 1682
rect -2793 1648 -2625 1682
rect -2535 1648 -2367 1682
rect -2277 1648 -2109 1682
rect -2019 1648 -1851 1682
rect -1761 1648 -1593 1682
rect -1503 1648 -1335 1682
rect -1245 1648 -1077 1682
rect -987 1648 -819 1682
rect -729 1648 -561 1682
rect -471 1648 -303 1682
rect -213 1648 -45 1682
rect 45 1648 213 1682
rect 303 1648 471 1682
rect 561 1648 729 1682
rect 819 1648 987 1682
rect 1077 1648 1245 1682
rect 1335 1648 1503 1682
rect 1593 1648 1761 1682
rect 1851 1648 2019 1682
rect 2109 1648 2277 1682
rect 2367 1648 2535 1682
rect 2625 1648 2793 1682
rect 2883 1648 3051 1682
rect 3141 1648 3309 1682
rect 3399 1648 3567 1682
rect 3657 1648 3825 1682
rect 3915 1648 4083 1682
rect 4173 1648 4341 1682
rect 4431 1648 4599 1682
rect 4689 1648 4857 1682
rect 4947 1648 5115 1682
rect 5205 1648 5373 1682
rect 5463 1648 5631 1682
rect -5693 622 -5659 1598
rect -5435 622 -5401 1598
rect -5177 622 -5143 1598
rect -4919 622 -4885 1598
rect -4661 622 -4627 1598
rect -4403 622 -4369 1598
rect -4145 622 -4111 1598
rect -3887 622 -3853 1598
rect -3629 622 -3595 1598
rect -3371 622 -3337 1598
rect -3113 622 -3079 1598
rect -2855 622 -2821 1598
rect -2597 622 -2563 1598
rect -2339 622 -2305 1598
rect -2081 622 -2047 1598
rect -1823 622 -1789 1598
rect -1565 622 -1531 1598
rect -1307 622 -1273 1598
rect -1049 622 -1015 1598
rect -791 622 -757 1598
rect -533 622 -499 1598
rect -275 622 -241 1598
rect -17 622 17 1598
rect 241 622 275 1598
rect 499 622 533 1598
rect 757 622 791 1598
rect 1015 622 1049 1598
rect 1273 622 1307 1598
rect 1531 622 1565 1598
rect 1789 622 1823 1598
rect 2047 622 2081 1598
rect 2305 622 2339 1598
rect 2563 622 2597 1598
rect 2821 622 2855 1598
rect 3079 622 3113 1598
rect 3337 622 3371 1598
rect 3595 622 3629 1598
rect 3853 622 3887 1598
rect 4111 622 4145 1598
rect 4369 622 4403 1598
rect 4627 622 4661 1598
rect 4885 622 4919 1598
rect 5143 622 5177 1598
rect 5401 622 5435 1598
rect 5659 622 5693 1598
rect -5631 538 -5463 572
rect -5373 538 -5205 572
rect -5115 538 -4947 572
rect -4857 538 -4689 572
rect -4599 538 -4431 572
rect -4341 538 -4173 572
rect -4083 538 -3915 572
rect -3825 538 -3657 572
rect -3567 538 -3399 572
rect -3309 538 -3141 572
rect -3051 538 -2883 572
rect -2793 538 -2625 572
rect -2535 538 -2367 572
rect -2277 538 -2109 572
rect -2019 538 -1851 572
rect -1761 538 -1593 572
rect -1503 538 -1335 572
rect -1245 538 -1077 572
rect -987 538 -819 572
rect -729 538 -561 572
rect -471 538 -303 572
rect -213 538 -45 572
rect 45 538 213 572
rect 303 538 471 572
rect 561 538 729 572
rect 819 538 987 572
rect 1077 538 1245 572
rect 1335 538 1503 572
rect 1593 538 1761 572
rect 1851 538 2019 572
rect 2109 538 2277 572
rect 2367 538 2535 572
rect 2625 538 2793 572
rect 2883 538 3051 572
rect 3141 538 3309 572
rect 3399 538 3567 572
rect 3657 538 3825 572
rect 3915 538 4083 572
rect 4173 538 4341 572
rect 4431 538 4599 572
rect 4689 538 4857 572
rect 4947 538 5115 572
rect 5205 538 5373 572
rect 5463 538 5631 572
rect -5693 -488 -5659 488
rect -5435 -488 -5401 488
rect -5177 -488 -5143 488
rect -4919 -488 -4885 488
rect -4661 -488 -4627 488
rect -4403 -488 -4369 488
rect -4145 -488 -4111 488
rect -3887 -488 -3853 488
rect -3629 -488 -3595 488
rect -3371 -488 -3337 488
rect -3113 -488 -3079 488
rect -2855 -488 -2821 488
rect -2597 -488 -2563 488
rect -2339 -488 -2305 488
rect -2081 -488 -2047 488
rect -1823 -488 -1789 488
rect -1565 -488 -1531 488
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
rect 1531 -488 1565 488
rect 1789 -488 1823 488
rect 2047 -488 2081 488
rect 2305 -488 2339 488
rect 2563 -488 2597 488
rect 2821 -488 2855 488
rect 3079 -488 3113 488
rect 3337 -488 3371 488
rect 3595 -488 3629 488
rect 3853 -488 3887 488
rect 4111 -488 4145 488
rect 4369 -488 4403 488
rect 4627 -488 4661 488
rect 4885 -488 4919 488
rect 5143 -488 5177 488
rect 5401 -488 5435 488
rect 5659 -488 5693 488
rect -5631 -572 -5463 -538
rect -5373 -572 -5205 -538
rect -5115 -572 -4947 -538
rect -4857 -572 -4689 -538
rect -4599 -572 -4431 -538
rect -4341 -572 -4173 -538
rect -4083 -572 -3915 -538
rect -3825 -572 -3657 -538
rect -3567 -572 -3399 -538
rect -3309 -572 -3141 -538
rect -3051 -572 -2883 -538
rect -2793 -572 -2625 -538
rect -2535 -572 -2367 -538
rect -2277 -572 -2109 -538
rect -2019 -572 -1851 -538
rect -1761 -572 -1593 -538
rect -1503 -572 -1335 -538
rect -1245 -572 -1077 -538
rect -987 -572 -819 -538
rect -729 -572 -561 -538
rect -471 -572 -303 -538
rect -213 -572 -45 -538
rect 45 -572 213 -538
rect 303 -572 471 -538
rect 561 -572 729 -538
rect 819 -572 987 -538
rect 1077 -572 1245 -538
rect 1335 -572 1503 -538
rect 1593 -572 1761 -538
rect 1851 -572 2019 -538
rect 2109 -572 2277 -538
rect 2367 -572 2535 -538
rect 2625 -572 2793 -538
rect 2883 -572 3051 -538
rect 3141 -572 3309 -538
rect 3399 -572 3567 -538
rect 3657 -572 3825 -538
rect 3915 -572 4083 -538
rect 4173 -572 4341 -538
rect 4431 -572 4599 -538
rect 4689 -572 4857 -538
rect 4947 -572 5115 -538
rect 5205 -572 5373 -538
rect 5463 -572 5631 -538
rect -5693 -1598 -5659 -622
rect -5435 -1598 -5401 -622
rect -5177 -1598 -5143 -622
rect -4919 -1598 -4885 -622
rect -4661 -1598 -4627 -622
rect -4403 -1598 -4369 -622
rect -4145 -1598 -4111 -622
rect -3887 -1598 -3853 -622
rect -3629 -1598 -3595 -622
rect -3371 -1598 -3337 -622
rect -3113 -1598 -3079 -622
rect -2855 -1598 -2821 -622
rect -2597 -1598 -2563 -622
rect -2339 -1598 -2305 -622
rect -2081 -1598 -2047 -622
rect -1823 -1598 -1789 -622
rect -1565 -1598 -1531 -622
rect -1307 -1598 -1273 -622
rect -1049 -1598 -1015 -622
rect -791 -1598 -757 -622
rect -533 -1598 -499 -622
rect -275 -1598 -241 -622
rect -17 -1598 17 -622
rect 241 -1598 275 -622
rect 499 -1598 533 -622
rect 757 -1598 791 -622
rect 1015 -1598 1049 -622
rect 1273 -1598 1307 -622
rect 1531 -1598 1565 -622
rect 1789 -1598 1823 -622
rect 2047 -1598 2081 -622
rect 2305 -1598 2339 -622
rect 2563 -1598 2597 -622
rect 2821 -1598 2855 -622
rect 3079 -1598 3113 -622
rect 3337 -1598 3371 -622
rect 3595 -1598 3629 -622
rect 3853 -1598 3887 -622
rect 4111 -1598 4145 -622
rect 4369 -1598 4403 -622
rect 4627 -1598 4661 -622
rect 4885 -1598 4919 -622
rect 5143 -1598 5177 -622
rect 5401 -1598 5435 -622
rect 5659 -1598 5693 -622
rect -5631 -1682 -5463 -1648
rect -5373 -1682 -5205 -1648
rect -5115 -1682 -4947 -1648
rect -4857 -1682 -4689 -1648
rect -4599 -1682 -4431 -1648
rect -4341 -1682 -4173 -1648
rect -4083 -1682 -3915 -1648
rect -3825 -1682 -3657 -1648
rect -3567 -1682 -3399 -1648
rect -3309 -1682 -3141 -1648
rect -3051 -1682 -2883 -1648
rect -2793 -1682 -2625 -1648
rect -2535 -1682 -2367 -1648
rect -2277 -1682 -2109 -1648
rect -2019 -1682 -1851 -1648
rect -1761 -1682 -1593 -1648
rect -1503 -1682 -1335 -1648
rect -1245 -1682 -1077 -1648
rect -987 -1682 -819 -1648
rect -729 -1682 -561 -1648
rect -471 -1682 -303 -1648
rect -213 -1682 -45 -1648
rect 45 -1682 213 -1648
rect 303 -1682 471 -1648
rect 561 -1682 729 -1648
rect 819 -1682 987 -1648
rect 1077 -1682 1245 -1648
rect 1335 -1682 1503 -1648
rect 1593 -1682 1761 -1648
rect 1851 -1682 2019 -1648
rect 2109 -1682 2277 -1648
rect 2367 -1682 2535 -1648
rect 2625 -1682 2793 -1648
rect 2883 -1682 3051 -1648
rect 3141 -1682 3309 -1648
rect 3399 -1682 3567 -1648
rect 3657 -1682 3825 -1648
rect 3915 -1682 4083 -1648
rect 4173 -1682 4341 -1648
rect 4431 -1682 4599 -1648
rect 4689 -1682 4857 -1648
rect 4947 -1682 5115 -1648
rect 5205 -1682 5373 -1648
rect 5463 -1682 5631 -1648
rect -5693 -2708 -5659 -1732
rect -5435 -2708 -5401 -1732
rect -5177 -2708 -5143 -1732
rect -4919 -2708 -4885 -1732
rect -4661 -2708 -4627 -1732
rect -4403 -2708 -4369 -1732
rect -4145 -2708 -4111 -1732
rect -3887 -2708 -3853 -1732
rect -3629 -2708 -3595 -1732
rect -3371 -2708 -3337 -1732
rect -3113 -2708 -3079 -1732
rect -2855 -2708 -2821 -1732
rect -2597 -2708 -2563 -1732
rect -2339 -2708 -2305 -1732
rect -2081 -2708 -2047 -1732
rect -1823 -2708 -1789 -1732
rect -1565 -2708 -1531 -1732
rect -1307 -2708 -1273 -1732
rect -1049 -2708 -1015 -1732
rect -791 -2708 -757 -1732
rect -533 -2708 -499 -1732
rect -275 -2708 -241 -1732
rect -17 -2708 17 -1732
rect 241 -2708 275 -1732
rect 499 -2708 533 -1732
rect 757 -2708 791 -1732
rect 1015 -2708 1049 -1732
rect 1273 -2708 1307 -1732
rect 1531 -2708 1565 -1732
rect 1789 -2708 1823 -1732
rect 2047 -2708 2081 -1732
rect 2305 -2708 2339 -1732
rect 2563 -2708 2597 -1732
rect 2821 -2708 2855 -1732
rect 3079 -2708 3113 -1732
rect 3337 -2708 3371 -1732
rect 3595 -2708 3629 -1732
rect 3853 -2708 3887 -1732
rect 4111 -2708 4145 -1732
rect 4369 -2708 4403 -1732
rect 4627 -2708 4661 -1732
rect 4885 -2708 4919 -1732
rect 5143 -2708 5177 -1732
rect 5401 -2708 5435 -1732
rect 5659 -2708 5693 -1732
rect -5631 -2792 -5463 -2758
rect -5373 -2792 -5205 -2758
rect -5115 -2792 -4947 -2758
rect -4857 -2792 -4689 -2758
rect -4599 -2792 -4431 -2758
rect -4341 -2792 -4173 -2758
rect -4083 -2792 -3915 -2758
rect -3825 -2792 -3657 -2758
rect -3567 -2792 -3399 -2758
rect -3309 -2792 -3141 -2758
rect -3051 -2792 -2883 -2758
rect -2793 -2792 -2625 -2758
rect -2535 -2792 -2367 -2758
rect -2277 -2792 -2109 -2758
rect -2019 -2792 -1851 -2758
rect -1761 -2792 -1593 -2758
rect -1503 -2792 -1335 -2758
rect -1245 -2792 -1077 -2758
rect -987 -2792 -819 -2758
rect -729 -2792 -561 -2758
rect -471 -2792 -303 -2758
rect -213 -2792 -45 -2758
rect 45 -2792 213 -2758
rect 303 -2792 471 -2758
rect 561 -2792 729 -2758
rect 819 -2792 987 -2758
rect 1077 -2792 1245 -2758
rect 1335 -2792 1503 -2758
rect 1593 -2792 1761 -2758
rect 1851 -2792 2019 -2758
rect 2109 -2792 2277 -2758
rect 2367 -2792 2535 -2758
rect 2625 -2792 2793 -2758
rect 2883 -2792 3051 -2758
rect 3141 -2792 3309 -2758
rect 3399 -2792 3567 -2758
rect 3657 -2792 3825 -2758
rect 3915 -2792 4083 -2758
rect 4173 -2792 4341 -2758
rect 4431 -2792 4599 -2758
rect 4689 -2792 4857 -2758
rect 4947 -2792 5115 -2758
rect 5205 -2792 5373 -2758
rect 5463 -2792 5631 -2758
<< metal1 >>
rect -5643 2792 -5451 2798
rect -5643 2758 -5631 2792
rect -5463 2758 -5451 2792
rect -5643 2752 -5451 2758
rect -5385 2792 -5193 2798
rect -5385 2758 -5373 2792
rect -5205 2758 -5193 2792
rect -5385 2752 -5193 2758
rect -5127 2792 -4935 2798
rect -5127 2758 -5115 2792
rect -4947 2758 -4935 2792
rect -5127 2752 -4935 2758
rect -4869 2792 -4677 2798
rect -4869 2758 -4857 2792
rect -4689 2758 -4677 2792
rect -4869 2752 -4677 2758
rect -4611 2792 -4419 2798
rect -4611 2758 -4599 2792
rect -4431 2758 -4419 2792
rect -4611 2752 -4419 2758
rect -4353 2792 -4161 2798
rect -4353 2758 -4341 2792
rect -4173 2758 -4161 2792
rect -4353 2752 -4161 2758
rect -4095 2792 -3903 2798
rect -4095 2758 -4083 2792
rect -3915 2758 -3903 2792
rect -4095 2752 -3903 2758
rect -3837 2792 -3645 2798
rect -3837 2758 -3825 2792
rect -3657 2758 -3645 2792
rect -3837 2752 -3645 2758
rect -3579 2792 -3387 2798
rect -3579 2758 -3567 2792
rect -3399 2758 -3387 2792
rect -3579 2752 -3387 2758
rect -3321 2792 -3129 2798
rect -3321 2758 -3309 2792
rect -3141 2758 -3129 2792
rect -3321 2752 -3129 2758
rect -3063 2792 -2871 2798
rect -3063 2758 -3051 2792
rect -2883 2758 -2871 2792
rect -3063 2752 -2871 2758
rect -2805 2792 -2613 2798
rect -2805 2758 -2793 2792
rect -2625 2758 -2613 2792
rect -2805 2752 -2613 2758
rect -2547 2792 -2355 2798
rect -2547 2758 -2535 2792
rect -2367 2758 -2355 2792
rect -2547 2752 -2355 2758
rect -2289 2792 -2097 2798
rect -2289 2758 -2277 2792
rect -2109 2758 -2097 2792
rect -2289 2752 -2097 2758
rect -2031 2792 -1839 2798
rect -2031 2758 -2019 2792
rect -1851 2758 -1839 2792
rect -2031 2752 -1839 2758
rect -1773 2792 -1581 2798
rect -1773 2758 -1761 2792
rect -1593 2758 -1581 2792
rect -1773 2752 -1581 2758
rect -1515 2792 -1323 2798
rect -1515 2758 -1503 2792
rect -1335 2758 -1323 2792
rect -1515 2752 -1323 2758
rect -1257 2792 -1065 2798
rect -1257 2758 -1245 2792
rect -1077 2758 -1065 2792
rect -1257 2752 -1065 2758
rect -999 2792 -807 2798
rect -999 2758 -987 2792
rect -819 2758 -807 2792
rect -999 2752 -807 2758
rect -741 2792 -549 2798
rect -741 2758 -729 2792
rect -561 2758 -549 2792
rect -741 2752 -549 2758
rect -483 2792 -291 2798
rect -483 2758 -471 2792
rect -303 2758 -291 2792
rect -483 2752 -291 2758
rect -225 2792 -33 2798
rect -225 2758 -213 2792
rect -45 2758 -33 2792
rect -225 2752 -33 2758
rect 33 2792 225 2798
rect 33 2758 45 2792
rect 213 2758 225 2792
rect 33 2752 225 2758
rect 291 2792 483 2798
rect 291 2758 303 2792
rect 471 2758 483 2792
rect 291 2752 483 2758
rect 549 2792 741 2798
rect 549 2758 561 2792
rect 729 2758 741 2792
rect 549 2752 741 2758
rect 807 2792 999 2798
rect 807 2758 819 2792
rect 987 2758 999 2792
rect 807 2752 999 2758
rect 1065 2792 1257 2798
rect 1065 2758 1077 2792
rect 1245 2758 1257 2792
rect 1065 2752 1257 2758
rect 1323 2792 1515 2798
rect 1323 2758 1335 2792
rect 1503 2758 1515 2792
rect 1323 2752 1515 2758
rect 1581 2792 1773 2798
rect 1581 2758 1593 2792
rect 1761 2758 1773 2792
rect 1581 2752 1773 2758
rect 1839 2792 2031 2798
rect 1839 2758 1851 2792
rect 2019 2758 2031 2792
rect 1839 2752 2031 2758
rect 2097 2792 2289 2798
rect 2097 2758 2109 2792
rect 2277 2758 2289 2792
rect 2097 2752 2289 2758
rect 2355 2792 2547 2798
rect 2355 2758 2367 2792
rect 2535 2758 2547 2792
rect 2355 2752 2547 2758
rect 2613 2792 2805 2798
rect 2613 2758 2625 2792
rect 2793 2758 2805 2792
rect 2613 2752 2805 2758
rect 2871 2792 3063 2798
rect 2871 2758 2883 2792
rect 3051 2758 3063 2792
rect 2871 2752 3063 2758
rect 3129 2792 3321 2798
rect 3129 2758 3141 2792
rect 3309 2758 3321 2792
rect 3129 2752 3321 2758
rect 3387 2792 3579 2798
rect 3387 2758 3399 2792
rect 3567 2758 3579 2792
rect 3387 2752 3579 2758
rect 3645 2792 3837 2798
rect 3645 2758 3657 2792
rect 3825 2758 3837 2792
rect 3645 2752 3837 2758
rect 3903 2792 4095 2798
rect 3903 2758 3915 2792
rect 4083 2758 4095 2792
rect 3903 2752 4095 2758
rect 4161 2792 4353 2798
rect 4161 2758 4173 2792
rect 4341 2758 4353 2792
rect 4161 2752 4353 2758
rect 4419 2792 4611 2798
rect 4419 2758 4431 2792
rect 4599 2758 4611 2792
rect 4419 2752 4611 2758
rect 4677 2792 4869 2798
rect 4677 2758 4689 2792
rect 4857 2758 4869 2792
rect 4677 2752 4869 2758
rect 4935 2792 5127 2798
rect 4935 2758 4947 2792
rect 5115 2758 5127 2792
rect 4935 2752 5127 2758
rect 5193 2792 5385 2798
rect 5193 2758 5205 2792
rect 5373 2758 5385 2792
rect 5193 2752 5385 2758
rect 5451 2792 5643 2798
rect 5451 2758 5463 2792
rect 5631 2758 5643 2792
rect 5451 2752 5643 2758
rect -5699 2708 -5653 2720
rect -5699 1732 -5693 2708
rect -5659 1732 -5653 2708
rect -5699 1720 -5653 1732
rect -5441 2708 -5395 2720
rect -5441 1732 -5435 2708
rect -5401 1732 -5395 2708
rect -5441 1720 -5395 1732
rect -5183 2708 -5137 2720
rect -5183 1732 -5177 2708
rect -5143 1732 -5137 2708
rect -5183 1720 -5137 1732
rect -4925 2708 -4879 2720
rect -4925 1732 -4919 2708
rect -4885 1732 -4879 2708
rect -4925 1720 -4879 1732
rect -4667 2708 -4621 2720
rect -4667 1732 -4661 2708
rect -4627 1732 -4621 2708
rect -4667 1720 -4621 1732
rect -4409 2708 -4363 2720
rect -4409 1732 -4403 2708
rect -4369 1732 -4363 2708
rect -4409 1720 -4363 1732
rect -4151 2708 -4105 2720
rect -4151 1732 -4145 2708
rect -4111 1732 -4105 2708
rect -4151 1720 -4105 1732
rect -3893 2708 -3847 2720
rect -3893 1732 -3887 2708
rect -3853 1732 -3847 2708
rect -3893 1720 -3847 1732
rect -3635 2708 -3589 2720
rect -3635 1732 -3629 2708
rect -3595 1732 -3589 2708
rect -3635 1720 -3589 1732
rect -3377 2708 -3331 2720
rect -3377 1732 -3371 2708
rect -3337 1732 -3331 2708
rect -3377 1720 -3331 1732
rect -3119 2708 -3073 2720
rect -3119 1732 -3113 2708
rect -3079 1732 -3073 2708
rect -3119 1720 -3073 1732
rect -2861 2708 -2815 2720
rect -2861 1732 -2855 2708
rect -2821 1732 -2815 2708
rect -2861 1720 -2815 1732
rect -2603 2708 -2557 2720
rect -2603 1732 -2597 2708
rect -2563 1732 -2557 2708
rect -2603 1720 -2557 1732
rect -2345 2708 -2299 2720
rect -2345 1732 -2339 2708
rect -2305 1732 -2299 2708
rect -2345 1720 -2299 1732
rect -2087 2708 -2041 2720
rect -2087 1732 -2081 2708
rect -2047 1732 -2041 2708
rect -2087 1720 -2041 1732
rect -1829 2708 -1783 2720
rect -1829 1732 -1823 2708
rect -1789 1732 -1783 2708
rect -1829 1720 -1783 1732
rect -1571 2708 -1525 2720
rect -1571 1732 -1565 2708
rect -1531 1732 -1525 2708
rect -1571 1720 -1525 1732
rect -1313 2708 -1267 2720
rect -1313 1732 -1307 2708
rect -1273 1732 -1267 2708
rect -1313 1720 -1267 1732
rect -1055 2708 -1009 2720
rect -1055 1732 -1049 2708
rect -1015 1732 -1009 2708
rect -1055 1720 -1009 1732
rect -797 2708 -751 2720
rect -797 1732 -791 2708
rect -757 1732 -751 2708
rect -797 1720 -751 1732
rect -539 2708 -493 2720
rect -539 1732 -533 2708
rect -499 1732 -493 2708
rect -539 1720 -493 1732
rect -281 2708 -235 2720
rect -281 1732 -275 2708
rect -241 1732 -235 2708
rect -281 1720 -235 1732
rect -23 2708 23 2720
rect -23 1732 -17 2708
rect 17 1732 23 2708
rect -23 1720 23 1732
rect 235 2708 281 2720
rect 235 1732 241 2708
rect 275 1732 281 2708
rect 235 1720 281 1732
rect 493 2708 539 2720
rect 493 1732 499 2708
rect 533 1732 539 2708
rect 493 1720 539 1732
rect 751 2708 797 2720
rect 751 1732 757 2708
rect 791 1732 797 2708
rect 751 1720 797 1732
rect 1009 2708 1055 2720
rect 1009 1732 1015 2708
rect 1049 1732 1055 2708
rect 1009 1720 1055 1732
rect 1267 2708 1313 2720
rect 1267 1732 1273 2708
rect 1307 1732 1313 2708
rect 1267 1720 1313 1732
rect 1525 2708 1571 2720
rect 1525 1732 1531 2708
rect 1565 1732 1571 2708
rect 1525 1720 1571 1732
rect 1783 2708 1829 2720
rect 1783 1732 1789 2708
rect 1823 1732 1829 2708
rect 1783 1720 1829 1732
rect 2041 2708 2087 2720
rect 2041 1732 2047 2708
rect 2081 1732 2087 2708
rect 2041 1720 2087 1732
rect 2299 2708 2345 2720
rect 2299 1732 2305 2708
rect 2339 1732 2345 2708
rect 2299 1720 2345 1732
rect 2557 2708 2603 2720
rect 2557 1732 2563 2708
rect 2597 1732 2603 2708
rect 2557 1720 2603 1732
rect 2815 2708 2861 2720
rect 2815 1732 2821 2708
rect 2855 1732 2861 2708
rect 2815 1720 2861 1732
rect 3073 2708 3119 2720
rect 3073 1732 3079 2708
rect 3113 1732 3119 2708
rect 3073 1720 3119 1732
rect 3331 2708 3377 2720
rect 3331 1732 3337 2708
rect 3371 1732 3377 2708
rect 3331 1720 3377 1732
rect 3589 2708 3635 2720
rect 3589 1732 3595 2708
rect 3629 1732 3635 2708
rect 3589 1720 3635 1732
rect 3847 2708 3893 2720
rect 3847 1732 3853 2708
rect 3887 1732 3893 2708
rect 3847 1720 3893 1732
rect 4105 2708 4151 2720
rect 4105 1732 4111 2708
rect 4145 1732 4151 2708
rect 4105 1720 4151 1732
rect 4363 2708 4409 2720
rect 4363 1732 4369 2708
rect 4403 1732 4409 2708
rect 4363 1720 4409 1732
rect 4621 2708 4667 2720
rect 4621 1732 4627 2708
rect 4661 1732 4667 2708
rect 4621 1720 4667 1732
rect 4879 2708 4925 2720
rect 4879 1732 4885 2708
rect 4919 1732 4925 2708
rect 4879 1720 4925 1732
rect 5137 2708 5183 2720
rect 5137 1732 5143 2708
rect 5177 1732 5183 2708
rect 5137 1720 5183 1732
rect 5395 2708 5441 2720
rect 5395 1732 5401 2708
rect 5435 1732 5441 2708
rect 5395 1720 5441 1732
rect 5653 2708 5699 2720
rect 5653 1732 5659 2708
rect 5693 1732 5699 2708
rect 5653 1720 5699 1732
rect -5643 1682 -5451 1688
rect -5643 1648 -5631 1682
rect -5463 1648 -5451 1682
rect -5643 1642 -5451 1648
rect -5385 1682 -5193 1688
rect -5385 1648 -5373 1682
rect -5205 1648 -5193 1682
rect -5385 1642 -5193 1648
rect -5127 1682 -4935 1688
rect -5127 1648 -5115 1682
rect -4947 1648 -4935 1682
rect -5127 1642 -4935 1648
rect -4869 1682 -4677 1688
rect -4869 1648 -4857 1682
rect -4689 1648 -4677 1682
rect -4869 1642 -4677 1648
rect -4611 1682 -4419 1688
rect -4611 1648 -4599 1682
rect -4431 1648 -4419 1682
rect -4611 1642 -4419 1648
rect -4353 1682 -4161 1688
rect -4353 1648 -4341 1682
rect -4173 1648 -4161 1682
rect -4353 1642 -4161 1648
rect -4095 1682 -3903 1688
rect -4095 1648 -4083 1682
rect -3915 1648 -3903 1682
rect -4095 1642 -3903 1648
rect -3837 1682 -3645 1688
rect -3837 1648 -3825 1682
rect -3657 1648 -3645 1682
rect -3837 1642 -3645 1648
rect -3579 1682 -3387 1688
rect -3579 1648 -3567 1682
rect -3399 1648 -3387 1682
rect -3579 1642 -3387 1648
rect -3321 1682 -3129 1688
rect -3321 1648 -3309 1682
rect -3141 1648 -3129 1682
rect -3321 1642 -3129 1648
rect -3063 1682 -2871 1688
rect -3063 1648 -3051 1682
rect -2883 1648 -2871 1682
rect -3063 1642 -2871 1648
rect -2805 1682 -2613 1688
rect -2805 1648 -2793 1682
rect -2625 1648 -2613 1682
rect -2805 1642 -2613 1648
rect -2547 1682 -2355 1688
rect -2547 1648 -2535 1682
rect -2367 1648 -2355 1682
rect -2547 1642 -2355 1648
rect -2289 1682 -2097 1688
rect -2289 1648 -2277 1682
rect -2109 1648 -2097 1682
rect -2289 1642 -2097 1648
rect -2031 1682 -1839 1688
rect -2031 1648 -2019 1682
rect -1851 1648 -1839 1682
rect -2031 1642 -1839 1648
rect -1773 1682 -1581 1688
rect -1773 1648 -1761 1682
rect -1593 1648 -1581 1682
rect -1773 1642 -1581 1648
rect -1515 1682 -1323 1688
rect -1515 1648 -1503 1682
rect -1335 1648 -1323 1682
rect -1515 1642 -1323 1648
rect -1257 1682 -1065 1688
rect -1257 1648 -1245 1682
rect -1077 1648 -1065 1682
rect -1257 1642 -1065 1648
rect -999 1682 -807 1688
rect -999 1648 -987 1682
rect -819 1648 -807 1682
rect -999 1642 -807 1648
rect -741 1682 -549 1688
rect -741 1648 -729 1682
rect -561 1648 -549 1682
rect -741 1642 -549 1648
rect -483 1682 -291 1688
rect -483 1648 -471 1682
rect -303 1648 -291 1682
rect -483 1642 -291 1648
rect -225 1682 -33 1688
rect -225 1648 -213 1682
rect -45 1648 -33 1682
rect -225 1642 -33 1648
rect 33 1682 225 1688
rect 33 1648 45 1682
rect 213 1648 225 1682
rect 33 1642 225 1648
rect 291 1682 483 1688
rect 291 1648 303 1682
rect 471 1648 483 1682
rect 291 1642 483 1648
rect 549 1682 741 1688
rect 549 1648 561 1682
rect 729 1648 741 1682
rect 549 1642 741 1648
rect 807 1682 999 1688
rect 807 1648 819 1682
rect 987 1648 999 1682
rect 807 1642 999 1648
rect 1065 1682 1257 1688
rect 1065 1648 1077 1682
rect 1245 1648 1257 1682
rect 1065 1642 1257 1648
rect 1323 1682 1515 1688
rect 1323 1648 1335 1682
rect 1503 1648 1515 1682
rect 1323 1642 1515 1648
rect 1581 1682 1773 1688
rect 1581 1648 1593 1682
rect 1761 1648 1773 1682
rect 1581 1642 1773 1648
rect 1839 1682 2031 1688
rect 1839 1648 1851 1682
rect 2019 1648 2031 1682
rect 1839 1642 2031 1648
rect 2097 1682 2289 1688
rect 2097 1648 2109 1682
rect 2277 1648 2289 1682
rect 2097 1642 2289 1648
rect 2355 1682 2547 1688
rect 2355 1648 2367 1682
rect 2535 1648 2547 1682
rect 2355 1642 2547 1648
rect 2613 1682 2805 1688
rect 2613 1648 2625 1682
rect 2793 1648 2805 1682
rect 2613 1642 2805 1648
rect 2871 1682 3063 1688
rect 2871 1648 2883 1682
rect 3051 1648 3063 1682
rect 2871 1642 3063 1648
rect 3129 1682 3321 1688
rect 3129 1648 3141 1682
rect 3309 1648 3321 1682
rect 3129 1642 3321 1648
rect 3387 1682 3579 1688
rect 3387 1648 3399 1682
rect 3567 1648 3579 1682
rect 3387 1642 3579 1648
rect 3645 1682 3837 1688
rect 3645 1648 3657 1682
rect 3825 1648 3837 1682
rect 3645 1642 3837 1648
rect 3903 1682 4095 1688
rect 3903 1648 3915 1682
rect 4083 1648 4095 1682
rect 3903 1642 4095 1648
rect 4161 1682 4353 1688
rect 4161 1648 4173 1682
rect 4341 1648 4353 1682
rect 4161 1642 4353 1648
rect 4419 1682 4611 1688
rect 4419 1648 4431 1682
rect 4599 1648 4611 1682
rect 4419 1642 4611 1648
rect 4677 1682 4869 1688
rect 4677 1648 4689 1682
rect 4857 1648 4869 1682
rect 4677 1642 4869 1648
rect 4935 1682 5127 1688
rect 4935 1648 4947 1682
rect 5115 1648 5127 1682
rect 4935 1642 5127 1648
rect 5193 1682 5385 1688
rect 5193 1648 5205 1682
rect 5373 1648 5385 1682
rect 5193 1642 5385 1648
rect 5451 1682 5643 1688
rect 5451 1648 5463 1682
rect 5631 1648 5643 1682
rect 5451 1642 5643 1648
rect -5699 1598 -5653 1610
rect -5699 622 -5693 1598
rect -5659 622 -5653 1598
rect -5699 610 -5653 622
rect -5441 1598 -5395 1610
rect -5441 622 -5435 1598
rect -5401 622 -5395 1598
rect -5441 610 -5395 622
rect -5183 1598 -5137 1610
rect -5183 622 -5177 1598
rect -5143 622 -5137 1598
rect -5183 610 -5137 622
rect -4925 1598 -4879 1610
rect -4925 622 -4919 1598
rect -4885 622 -4879 1598
rect -4925 610 -4879 622
rect -4667 1598 -4621 1610
rect -4667 622 -4661 1598
rect -4627 622 -4621 1598
rect -4667 610 -4621 622
rect -4409 1598 -4363 1610
rect -4409 622 -4403 1598
rect -4369 622 -4363 1598
rect -4409 610 -4363 622
rect -4151 1598 -4105 1610
rect -4151 622 -4145 1598
rect -4111 622 -4105 1598
rect -4151 610 -4105 622
rect -3893 1598 -3847 1610
rect -3893 622 -3887 1598
rect -3853 622 -3847 1598
rect -3893 610 -3847 622
rect -3635 1598 -3589 1610
rect -3635 622 -3629 1598
rect -3595 622 -3589 1598
rect -3635 610 -3589 622
rect -3377 1598 -3331 1610
rect -3377 622 -3371 1598
rect -3337 622 -3331 1598
rect -3377 610 -3331 622
rect -3119 1598 -3073 1610
rect -3119 622 -3113 1598
rect -3079 622 -3073 1598
rect -3119 610 -3073 622
rect -2861 1598 -2815 1610
rect -2861 622 -2855 1598
rect -2821 622 -2815 1598
rect -2861 610 -2815 622
rect -2603 1598 -2557 1610
rect -2603 622 -2597 1598
rect -2563 622 -2557 1598
rect -2603 610 -2557 622
rect -2345 1598 -2299 1610
rect -2345 622 -2339 1598
rect -2305 622 -2299 1598
rect -2345 610 -2299 622
rect -2087 1598 -2041 1610
rect -2087 622 -2081 1598
rect -2047 622 -2041 1598
rect -2087 610 -2041 622
rect -1829 1598 -1783 1610
rect -1829 622 -1823 1598
rect -1789 622 -1783 1598
rect -1829 610 -1783 622
rect -1571 1598 -1525 1610
rect -1571 622 -1565 1598
rect -1531 622 -1525 1598
rect -1571 610 -1525 622
rect -1313 1598 -1267 1610
rect -1313 622 -1307 1598
rect -1273 622 -1267 1598
rect -1313 610 -1267 622
rect -1055 1598 -1009 1610
rect -1055 622 -1049 1598
rect -1015 622 -1009 1598
rect -1055 610 -1009 622
rect -797 1598 -751 1610
rect -797 622 -791 1598
rect -757 622 -751 1598
rect -797 610 -751 622
rect -539 1598 -493 1610
rect -539 622 -533 1598
rect -499 622 -493 1598
rect -539 610 -493 622
rect -281 1598 -235 1610
rect -281 622 -275 1598
rect -241 622 -235 1598
rect -281 610 -235 622
rect -23 1598 23 1610
rect -23 622 -17 1598
rect 17 622 23 1598
rect -23 610 23 622
rect 235 1598 281 1610
rect 235 622 241 1598
rect 275 622 281 1598
rect 235 610 281 622
rect 493 1598 539 1610
rect 493 622 499 1598
rect 533 622 539 1598
rect 493 610 539 622
rect 751 1598 797 1610
rect 751 622 757 1598
rect 791 622 797 1598
rect 751 610 797 622
rect 1009 1598 1055 1610
rect 1009 622 1015 1598
rect 1049 622 1055 1598
rect 1009 610 1055 622
rect 1267 1598 1313 1610
rect 1267 622 1273 1598
rect 1307 622 1313 1598
rect 1267 610 1313 622
rect 1525 1598 1571 1610
rect 1525 622 1531 1598
rect 1565 622 1571 1598
rect 1525 610 1571 622
rect 1783 1598 1829 1610
rect 1783 622 1789 1598
rect 1823 622 1829 1598
rect 1783 610 1829 622
rect 2041 1598 2087 1610
rect 2041 622 2047 1598
rect 2081 622 2087 1598
rect 2041 610 2087 622
rect 2299 1598 2345 1610
rect 2299 622 2305 1598
rect 2339 622 2345 1598
rect 2299 610 2345 622
rect 2557 1598 2603 1610
rect 2557 622 2563 1598
rect 2597 622 2603 1598
rect 2557 610 2603 622
rect 2815 1598 2861 1610
rect 2815 622 2821 1598
rect 2855 622 2861 1598
rect 2815 610 2861 622
rect 3073 1598 3119 1610
rect 3073 622 3079 1598
rect 3113 622 3119 1598
rect 3073 610 3119 622
rect 3331 1598 3377 1610
rect 3331 622 3337 1598
rect 3371 622 3377 1598
rect 3331 610 3377 622
rect 3589 1598 3635 1610
rect 3589 622 3595 1598
rect 3629 622 3635 1598
rect 3589 610 3635 622
rect 3847 1598 3893 1610
rect 3847 622 3853 1598
rect 3887 622 3893 1598
rect 3847 610 3893 622
rect 4105 1598 4151 1610
rect 4105 622 4111 1598
rect 4145 622 4151 1598
rect 4105 610 4151 622
rect 4363 1598 4409 1610
rect 4363 622 4369 1598
rect 4403 622 4409 1598
rect 4363 610 4409 622
rect 4621 1598 4667 1610
rect 4621 622 4627 1598
rect 4661 622 4667 1598
rect 4621 610 4667 622
rect 4879 1598 4925 1610
rect 4879 622 4885 1598
rect 4919 622 4925 1598
rect 4879 610 4925 622
rect 5137 1598 5183 1610
rect 5137 622 5143 1598
rect 5177 622 5183 1598
rect 5137 610 5183 622
rect 5395 1598 5441 1610
rect 5395 622 5401 1598
rect 5435 622 5441 1598
rect 5395 610 5441 622
rect 5653 1598 5699 1610
rect 5653 622 5659 1598
rect 5693 622 5699 1598
rect 5653 610 5699 622
rect -5643 572 -5451 578
rect -5643 538 -5631 572
rect -5463 538 -5451 572
rect -5643 532 -5451 538
rect -5385 572 -5193 578
rect -5385 538 -5373 572
rect -5205 538 -5193 572
rect -5385 532 -5193 538
rect -5127 572 -4935 578
rect -5127 538 -5115 572
rect -4947 538 -4935 572
rect -5127 532 -4935 538
rect -4869 572 -4677 578
rect -4869 538 -4857 572
rect -4689 538 -4677 572
rect -4869 532 -4677 538
rect -4611 572 -4419 578
rect -4611 538 -4599 572
rect -4431 538 -4419 572
rect -4611 532 -4419 538
rect -4353 572 -4161 578
rect -4353 538 -4341 572
rect -4173 538 -4161 572
rect -4353 532 -4161 538
rect -4095 572 -3903 578
rect -4095 538 -4083 572
rect -3915 538 -3903 572
rect -4095 532 -3903 538
rect -3837 572 -3645 578
rect -3837 538 -3825 572
rect -3657 538 -3645 572
rect -3837 532 -3645 538
rect -3579 572 -3387 578
rect -3579 538 -3567 572
rect -3399 538 -3387 572
rect -3579 532 -3387 538
rect -3321 572 -3129 578
rect -3321 538 -3309 572
rect -3141 538 -3129 572
rect -3321 532 -3129 538
rect -3063 572 -2871 578
rect -3063 538 -3051 572
rect -2883 538 -2871 572
rect -3063 532 -2871 538
rect -2805 572 -2613 578
rect -2805 538 -2793 572
rect -2625 538 -2613 572
rect -2805 532 -2613 538
rect -2547 572 -2355 578
rect -2547 538 -2535 572
rect -2367 538 -2355 572
rect -2547 532 -2355 538
rect -2289 572 -2097 578
rect -2289 538 -2277 572
rect -2109 538 -2097 572
rect -2289 532 -2097 538
rect -2031 572 -1839 578
rect -2031 538 -2019 572
rect -1851 538 -1839 572
rect -2031 532 -1839 538
rect -1773 572 -1581 578
rect -1773 538 -1761 572
rect -1593 538 -1581 572
rect -1773 532 -1581 538
rect -1515 572 -1323 578
rect -1515 538 -1503 572
rect -1335 538 -1323 572
rect -1515 532 -1323 538
rect -1257 572 -1065 578
rect -1257 538 -1245 572
rect -1077 538 -1065 572
rect -1257 532 -1065 538
rect -999 572 -807 578
rect -999 538 -987 572
rect -819 538 -807 572
rect -999 532 -807 538
rect -741 572 -549 578
rect -741 538 -729 572
rect -561 538 -549 572
rect -741 532 -549 538
rect -483 572 -291 578
rect -483 538 -471 572
rect -303 538 -291 572
rect -483 532 -291 538
rect -225 572 -33 578
rect -225 538 -213 572
rect -45 538 -33 572
rect -225 532 -33 538
rect 33 572 225 578
rect 33 538 45 572
rect 213 538 225 572
rect 33 532 225 538
rect 291 572 483 578
rect 291 538 303 572
rect 471 538 483 572
rect 291 532 483 538
rect 549 572 741 578
rect 549 538 561 572
rect 729 538 741 572
rect 549 532 741 538
rect 807 572 999 578
rect 807 538 819 572
rect 987 538 999 572
rect 807 532 999 538
rect 1065 572 1257 578
rect 1065 538 1077 572
rect 1245 538 1257 572
rect 1065 532 1257 538
rect 1323 572 1515 578
rect 1323 538 1335 572
rect 1503 538 1515 572
rect 1323 532 1515 538
rect 1581 572 1773 578
rect 1581 538 1593 572
rect 1761 538 1773 572
rect 1581 532 1773 538
rect 1839 572 2031 578
rect 1839 538 1851 572
rect 2019 538 2031 572
rect 1839 532 2031 538
rect 2097 572 2289 578
rect 2097 538 2109 572
rect 2277 538 2289 572
rect 2097 532 2289 538
rect 2355 572 2547 578
rect 2355 538 2367 572
rect 2535 538 2547 572
rect 2355 532 2547 538
rect 2613 572 2805 578
rect 2613 538 2625 572
rect 2793 538 2805 572
rect 2613 532 2805 538
rect 2871 572 3063 578
rect 2871 538 2883 572
rect 3051 538 3063 572
rect 2871 532 3063 538
rect 3129 572 3321 578
rect 3129 538 3141 572
rect 3309 538 3321 572
rect 3129 532 3321 538
rect 3387 572 3579 578
rect 3387 538 3399 572
rect 3567 538 3579 572
rect 3387 532 3579 538
rect 3645 572 3837 578
rect 3645 538 3657 572
rect 3825 538 3837 572
rect 3645 532 3837 538
rect 3903 572 4095 578
rect 3903 538 3915 572
rect 4083 538 4095 572
rect 3903 532 4095 538
rect 4161 572 4353 578
rect 4161 538 4173 572
rect 4341 538 4353 572
rect 4161 532 4353 538
rect 4419 572 4611 578
rect 4419 538 4431 572
rect 4599 538 4611 572
rect 4419 532 4611 538
rect 4677 572 4869 578
rect 4677 538 4689 572
rect 4857 538 4869 572
rect 4677 532 4869 538
rect 4935 572 5127 578
rect 4935 538 4947 572
rect 5115 538 5127 572
rect 4935 532 5127 538
rect 5193 572 5385 578
rect 5193 538 5205 572
rect 5373 538 5385 572
rect 5193 532 5385 538
rect 5451 572 5643 578
rect 5451 538 5463 572
rect 5631 538 5643 572
rect 5451 532 5643 538
rect -5699 488 -5653 500
rect -5699 -488 -5693 488
rect -5659 -488 -5653 488
rect -5699 -500 -5653 -488
rect -5441 488 -5395 500
rect -5441 -488 -5435 488
rect -5401 -488 -5395 488
rect -5441 -500 -5395 -488
rect -5183 488 -5137 500
rect -5183 -488 -5177 488
rect -5143 -488 -5137 488
rect -5183 -500 -5137 -488
rect -4925 488 -4879 500
rect -4925 -488 -4919 488
rect -4885 -488 -4879 488
rect -4925 -500 -4879 -488
rect -4667 488 -4621 500
rect -4667 -488 -4661 488
rect -4627 -488 -4621 488
rect -4667 -500 -4621 -488
rect -4409 488 -4363 500
rect -4409 -488 -4403 488
rect -4369 -488 -4363 488
rect -4409 -500 -4363 -488
rect -4151 488 -4105 500
rect -4151 -488 -4145 488
rect -4111 -488 -4105 488
rect -4151 -500 -4105 -488
rect -3893 488 -3847 500
rect -3893 -488 -3887 488
rect -3853 -488 -3847 488
rect -3893 -500 -3847 -488
rect -3635 488 -3589 500
rect -3635 -488 -3629 488
rect -3595 -488 -3589 488
rect -3635 -500 -3589 -488
rect -3377 488 -3331 500
rect -3377 -488 -3371 488
rect -3337 -488 -3331 488
rect -3377 -500 -3331 -488
rect -3119 488 -3073 500
rect -3119 -488 -3113 488
rect -3079 -488 -3073 488
rect -3119 -500 -3073 -488
rect -2861 488 -2815 500
rect -2861 -488 -2855 488
rect -2821 -488 -2815 488
rect -2861 -500 -2815 -488
rect -2603 488 -2557 500
rect -2603 -488 -2597 488
rect -2563 -488 -2557 488
rect -2603 -500 -2557 -488
rect -2345 488 -2299 500
rect -2345 -488 -2339 488
rect -2305 -488 -2299 488
rect -2345 -500 -2299 -488
rect -2087 488 -2041 500
rect -2087 -488 -2081 488
rect -2047 -488 -2041 488
rect -2087 -500 -2041 -488
rect -1829 488 -1783 500
rect -1829 -488 -1823 488
rect -1789 -488 -1783 488
rect -1829 -500 -1783 -488
rect -1571 488 -1525 500
rect -1571 -488 -1565 488
rect -1531 -488 -1525 488
rect -1571 -500 -1525 -488
rect -1313 488 -1267 500
rect -1313 -488 -1307 488
rect -1273 -488 -1267 488
rect -1313 -500 -1267 -488
rect -1055 488 -1009 500
rect -1055 -488 -1049 488
rect -1015 -488 -1009 488
rect -1055 -500 -1009 -488
rect -797 488 -751 500
rect -797 -488 -791 488
rect -757 -488 -751 488
rect -797 -500 -751 -488
rect -539 488 -493 500
rect -539 -488 -533 488
rect -499 -488 -493 488
rect -539 -500 -493 -488
rect -281 488 -235 500
rect -281 -488 -275 488
rect -241 -488 -235 488
rect -281 -500 -235 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 235 488 281 500
rect 235 -488 241 488
rect 275 -488 281 488
rect 235 -500 281 -488
rect 493 488 539 500
rect 493 -488 499 488
rect 533 -488 539 488
rect 493 -500 539 -488
rect 751 488 797 500
rect 751 -488 757 488
rect 791 -488 797 488
rect 751 -500 797 -488
rect 1009 488 1055 500
rect 1009 -488 1015 488
rect 1049 -488 1055 488
rect 1009 -500 1055 -488
rect 1267 488 1313 500
rect 1267 -488 1273 488
rect 1307 -488 1313 488
rect 1267 -500 1313 -488
rect 1525 488 1571 500
rect 1525 -488 1531 488
rect 1565 -488 1571 488
rect 1525 -500 1571 -488
rect 1783 488 1829 500
rect 1783 -488 1789 488
rect 1823 -488 1829 488
rect 1783 -500 1829 -488
rect 2041 488 2087 500
rect 2041 -488 2047 488
rect 2081 -488 2087 488
rect 2041 -500 2087 -488
rect 2299 488 2345 500
rect 2299 -488 2305 488
rect 2339 -488 2345 488
rect 2299 -500 2345 -488
rect 2557 488 2603 500
rect 2557 -488 2563 488
rect 2597 -488 2603 488
rect 2557 -500 2603 -488
rect 2815 488 2861 500
rect 2815 -488 2821 488
rect 2855 -488 2861 488
rect 2815 -500 2861 -488
rect 3073 488 3119 500
rect 3073 -488 3079 488
rect 3113 -488 3119 488
rect 3073 -500 3119 -488
rect 3331 488 3377 500
rect 3331 -488 3337 488
rect 3371 -488 3377 488
rect 3331 -500 3377 -488
rect 3589 488 3635 500
rect 3589 -488 3595 488
rect 3629 -488 3635 488
rect 3589 -500 3635 -488
rect 3847 488 3893 500
rect 3847 -488 3853 488
rect 3887 -488 3893 488
rect 3847 -500 3893 -488
rect 4105 488 4151 500
rect 4105 -488 4111 488
rect 4145 -488 4151 488
rect 4105 -500 4151 -488
rect 4363 488 4409 500
rect 4363 -488 4369 488
rect 4403 -488 4409 488
rect 4363 -500 4409 -488
rect 4621 488 4667 500
rect 4621 -488 4627 488
rect 4661 -488 4667 488
rect 4621 -500 4667 -488
rect 4879 488 4925 500
rect 4879 -488 4885 488
rect 4919 -488 4925 488
rect 4879 -500 4925 -488
rect 5137 488 5183 500
rect 5137 -488 5143 488
rect 5177 -488 5183 488
rect 5137 -500 5183 -488
rect 5395 488 5441 500
rect 5395 -488 5401 488
rect 5435 -488 5441 488
rect 5395 -500 5441 -488
rect 5653 488 5699 500
rect 5653 -488 5659 488
rect 5693 -488 5699 488
rect 5653 -500 5699 -488
rect -5643 -538 -5451 -532
rect -5643 -572 -5631 -538
rect -5463 -572 -5451 -538
rect -5643 -578 -5451 -572
rect -5385 -538 -5193 -532
rect -5385 -572 -5373 -538
rect -5205 -572 -5193 -538
rect -5385 -578 -5193 -572
rect -5127 -538 -4935 -532
rect -5127 -572 -5115 -538
rect -4947 -572 -4935 -538
rect -5127 -578 -4935 -572
rect -4869 -538 -4677 -532
rect -4869 -572 -4857 -538
rect -4689 -572 -4677 -538
rect -4869 -578 -4677 -572
rect -4611 -538 -4419 -532
rect -4611 -572 -4599 -538
rect -4431 -572 -4419 -538
rect -4611 -578 -4419 -572
rect -4353 -538 -4161 -532
rect -4353 -572 -4341 -538
rect -4173 -572 -4161 -538
rect -4353 -578 -4161 -572
rect -4095 -538 -3903 -532
rect -4095 -572 -4083 -538
rect -3915 -572 -3903 -538
rect -4095 -578 -3903 -572
rect -3837 -538 -3645 -532
rect -3837 -572 -3825 -538
rect -3657 -572 -3645 -538
rect -3837 -578 -3645 -572
rect -3579 -538 -3387 -532
rect -3579 -572 -3567 -538
rect -3399 -572 -3387 -538
rect -3579 -578 -3387 -572
rect -3321 -538 -3129 -532
rect -3321 -572 -3309 -538
rect -3141 -572 -3129 -538
rect -3321 -578 -3129 -572
rect -3063 -538 -2871 -532
rect -3063 -572 -3051 -538
rect -2883 -572 -2871 -538
rect -3063 -578 -2871 -572
rect -2805 -538 -2613 -532
rect -2805 -572 -2793 -538
rect -2625 -572 -2613 -538
rect -2805 -578 -2613 -572
rect -2547 -538 -2355 -532
rect -2547 -572 -2535 -538
rect -2367 -572 -2355 -538
rect -2547 -578 -2355 -572
rect -2289 -538 -2097 -532
rect -2289 -572 -2277 -538
rect -2109 -572 -2097 -538
rect -2289 -578 -2097 -572
rect -2031 -538 -1839 -532
rect -2031 -572 -2019 -538
rect -1851 -572 -1839 -538
rect -2031 -578 -1839 -572
rect -1773 -538 -1581 -532
rect -1773 -572 -1761 -538
rect -1593 -572 -1581 -538
rect -1773 -578 -1581 -572
rect -1515 -538 -1323 -532
rect -1515 -572 -1503 -538
rect -1335 -572 -1323 -538
rect -1515 -578 -1323 -572
rect -1257 -538 -1065 -532
rect -1257 -572 -1245 -538
rect -1077 -572 -1065 -538
rect -1257 -578 -1065 -572
rect -999 -538 -807 -532
rect -999 -572 -987 -538
rect -819 -572 -807 -538
rect -999 -578 -807 -572
rect -741 -538 -549 -532
rect -741 -572 -729 -538
rect -561 -572 -549 -538
rect -741 -578 -549 -572
rect -483 -538 -291 -532
rect -483 -572 -471 -538
rect -303 -572 -291 -538
rect -483 -578 -291 -572
rect -225 -538 -33 -532
rect -225 -572 -213 -538
rect -45 -572 -33 -538
rect -225 -578 -33 -572
rect 33 -538 225 -532
rect 33 -572 45 -538
rect 213 -572 225 -538
rect 33 -578 225 -572
rect 291 -538 483 -532
rect 291 -572 303 -538
rect 471 -572 483 -538
rect 291 -578 483 -572
rect 549 -538 741 -532
rect 549 -572 561 -538
rect 729 -572 741 -538
rect 549 -578 741 -572
rect 807 -538 999 -532
rect 807 -572 819 -538
rect 987 -572 999 -538
rect 807 -578 999 -572
rect 1065 -538 1257 -532
rect 1065 -572 1077 -538
rect 1245 -572 1257 -538
rect 1065 -578 1257 -572
rect 1323 -538 1515 -532
rect 1323 -572 1335 -538
rect 1503 -572 1515 -538
rect 1323 -578 1515 -572
rect 1581 -538 1773 -532
rect 1581 -572 1593 -538
rect 1761 -572 1773 -538
rect 1581 -578 1773 -572
rect 1839 -538 2031 -532
rect 1839 -572 1851 -538
rect 2019 -572 2031 -538
rect 1839 -578 2031 -572
rect 2097 -538 2289 -532
rect 2097 -572 2109 -538
rect 2277 -572 2289 -538
rect 2097 -578 2289 -572
rect 2355 -538 2547 -532
rect 2355 -572 2367 -538
rect 2535 -572 2547 -538
rect 2355 -578 2547 -572
rect 2613 -538 2805 -532
rect 2613 -572 2625 -538
rect 2793 -572 2805 -538
rect 2613 -578 2805 -572
rect 2871 -538 3063 -532
rect 2871 -572 2883 -538
rect 3051 -572 3063 -538
rect 2871 -578 3063 -572
rect 3129 -538 3321 -532
rect 3129 -572 3141 -538
rect 3309 -572 3321 -538
rect 3129 -578 3321 -572
rect 3387 -538 3579 -532
rect 3387 -572 3399 -538
rect 3567 -572 3579 -538
rect 3387 -578 3579 -572
rect 3645 -538 3837 -532
rect 3645 -572 3657 -538
rect 3825 -572 3837 -538
rect 3645 -578 3837 -572
rect 3903 -538 4095 -532
rect 3903 -572 3915 -538
rect 4083 -572 4095 -538
rect 3903 -578 4095 -572
rect 4161 -538 4353 -532
rect 4161 -572 4173 -538
rect 4341 -572 4353 -538
rect 4161 -578 4353 -572
rect 4419 -538 4611 -532
rect 4419 -572 4431 -538
rect 4599 -572 4611 -538
rect 4419 -578 4611 -572
rect 4677 -538 4869 -532
rect 4677 -572 4689 -538
rect 4857 -572 4869 -538
rect 4677 -578 4869 -572
rect 4935 -538 5127 -532
rect 4935 -572 4947 -538
rect 5115 -572 5127 -538
rect 4935 -578 5127 -572
rect 5193 -538 5385 -532
rect 5193 -572 5205 -538
rect 5373 -572 5385 -538
rect 5193 -578 5385 -572
rect 5451 -538 5643 -532
rect 5451 -572 5463 -538
rect 5631 -572 5643 -538
rect 5451 -578 5643 -572
rect -5699 -622 -5653 -610
rect -5699 -1598 -5693 -622
rect -5659 -1598 -5653 -622
rect -5699 -1610 -5653 -1598
rect -5441 -622 -5395 -610
rect -5441 -1598 -5435 -622
rect -5401 -1598 -5395 -622
rect -5441 -1610 -5395 -1598
rect -5183 -622 -5137 -610
rect -5183 -1598 -5177 -622
rect -5143 -1598 -5137 -622
rect -5183 -1610 -5137 -1598
rect -4925 -622 -4879 -610
rect -4925 -1598 -4919 -622
rect -4885 -1598 -4879 -622
rect -4925 -1610 -4879 -1598
rect -4667 -622 -4621 -610
rect -4667 -1598 -4661 -622
rect -4627 -1598 -4621 -622
rect -4667 -1610 -4621 -1598
rect -4409 -622 -4363 -610
rect -4409 -1598 -4403 -622
rect -4369 -1598 -4363 -622
rect -4409 -1610 -4363 -1598
rect -4151 -622 -4105 -610
rect -4151 -1598 -4145 -622
rect -4111 -1598 -4105 -622
rect -4151 -1610 -4105 -1598
rect -3893 -622 -3847 -610
rect -3893 -1598 -3887 -622
rect -3853 -1598 -3847 -622
rect -3893 -1610 -3847 -1598
rect -3635 -622 -3589 -610
rect -3635 -1598 -3629 -622
rect -3595 -1598 -3589 -622
rect -3635 -1610 -3589 -1598
rect -3377 -622 -3331 -610
rect -3377 -1598 -3371 -622
rect -3337 -1598 -3331 -622
rect -3377 -1610 -3331 -1598
rect -3119 -622 -3073 -610
rect -3119 -1598 -3113 -622
rect -3079 -1598 -3073 -622
rect -3119 -1610 -3073 -1598
rect -2861 -622 -2815 -610
rect -2861 -1598 -2855 -622
rect -2821 -1598 -2815 -622
rect -2861 -1610 -2815 -1598
rect -2603 -622 -2557 -610
rect -2603 -1598 -2597 -622
rect -2563 -1598 -2557 -622
rect -2603 -1610 -2557 -1598
rect -2345 -622 -2299 -610
rect -2345 -1598 -2339 -622
rect -2305 -1598 -2299 -622
rect -2345 -1610 -2299 -1598
rect -2087 -622 -2041 -610
rect -2087 -1598 -2081 -622
rect -2047 -1598 -2041 -622
rect -2087 -1610 -2041 -1598
rect -1829 -622 -1783 -610
rect -1829 -1598 -1823 -622
rect -1789 -1598 -1783 -622
rect -1829 -1610 -1783 -1598
rect -1571 -622 -1525 -610
rect -1571 -1598 -1565 -622
rect -1531 -1598 -1525 -622
rect -1571 -1610 -1525 -1598
rect -1313 -622 -1267 -610
rect -1313 -1598 -1307 -622
rect -1273 -1598 -1267 -622
rect -1313 -1610 -1267 -1598
rect -1055 -622 -1009 -610
rect -1055 -1598 -1049 -622
rect -1015 -1598 -1009 -622
rect -1055 -1610 -1009 -1598
rect -797 -622 -751 -610
rect -797 -1598 -791 -622
rect -757 -1598 -751 -622
rect -797 -1610 -751 -1598
rect -539 -622 -493 -610
rect -539 -1598 -533 -622
rect -499 -1598 -493 -622
rect -539 -1610 -493 -1598
rect -281 -622 -235 -610
rect -281 -1598 -275 -622
rect -241 -1598 -235 -622
rect -281 -1610 -235 -1598
rect -23 -622 23 -610
rect -23 -1598 -17 -622
rect 17 -1598 23 -622
rect -23 -1610 23 -1598
rect 235 -622 281 -610
rect 235 -1598 241 -622
rect 275 -1598 281 -622
rect 235 -1610 281 -1598
rect 493 -622 539 -610
rect 493 -1598 499 -622
rect 533 -1598 539 -622
rect 493 -1610 539 -1598
rect 751 -622 797 -610
rect 751 -1598 757 -622
rect 791 -1598 797 -622
rect 751 -1610 797 -1598
rect 1009 -622 1055 -610
rect 1009 -1598 1015 -622
rect 1049 -1598 1055 -622
rect 1009 -1610 1055 -1598
rect 1267 -622 1313 -610
rect 1267 -1598 1273 -622
rect 1307 -1598 1313 -622
rect 1267 -1610 1313 -1598
rect 1525 -622 1571 -610
rect 1525 -1598 1531 -622
rect 1565 -1598 1571 -622
rect 1525 -1610 1571 -1598
rect 1783 -622 1829 -610
rect 1783 -1598 1789 -622
rect 1823 -1598 1829 -622
rect 1783 -1610 1829 -1598
rect 2041 -622 2087 -610
rect 2041 -1598 2047 -622
rect 2081 -1598 2087 -622
rect 2041 -1610 2087 -1598
rect 2299 -622 2345 -610
rect 2299 -1598 2305 -622
rect 2339 -1598 2345 -622
rect 2299 -1610 2345 -1598
rect 2557 -622 2603 -610
rect 2557 -1598 2563 -622
rect 2597 -1598 2603 -622
rect 2557 -1610 2603 -1598
rect 2815 -622 2861 -610
rect 2815 -1598 2821 -622
rect 2855 -1598 2861 -622
rect 2815 -1610 2861 -1598
rect 3073 -622 3119 -610
rect 3073 -1598 3079 -622
rect 3113 -1598 3119 -622
rect 3073 -1610 3119 -1598
rect 3331 -622 3377 -610
rect 3331 -1598 3337 -622
rect 3371 -1598 3377 -622
rect 3331 -1610 3377 -1598
rect 3589 -622 3635 -610
rect 3589 -1598 3595 -622
rect 3629 -1598 3635 -622
rect 3589 -1610 3635 -1598
rect 3847 -622 3893 -610
rect 3847 -1598 3853 -622
rect 3887 -1598 3893 -622
rect 3847 -1610 3893 -1598
rect 4105 -622 4151 -610
rect 4105 -1598 4111 -622
rect 4145 -1598 4151 -622
rect 4105 -1610 4151 -1598
rect 4363 -622 4409 -610
rect 4363 -1598 4369 -622
rect 4403 -1598 4409 -622
rect 4363 -1610 4409 -1598
rect 4621 -622 4667 -610
rect 4621 -1598 4627 -622
rect 4661 -1598 4667 -622
rect 4621 -1610 4667 -1598
rect 4879 -622 4925 -610
rect 4879 -1598 4885 -622
rect 4919 -1598 4925 -622
rect 4879 -1610 4925 -1598
rect 5137 -622 5183 -610
rect 5137 -1598 5143 -622
rect 5177 -1598 5183 -622
rect 5137 -1610 5183 -1598
rect 5395 -622 5441 -610
rect 5395 -1598 5401 -622
rect 5435 -1598 5441 -622
rect 5395 -1610 5441 -1598
rect 5653 -622 5699 -610
rect 5653 -1598 5659 -622
rect 5693 -1598 5699 -622
rect 5653 -1610 5699 -1598
rect -5643 -1648 -5451 -1642
rect -5643 -1682 -5631 -1648
rect -5463 -1682 -5451 -1648
rect -5643 -1688 -5451 -1682
rect -5385 -1648 -5193 -1642
rect -5385 -1682 -5373 -1648
rect -5205 -1682 -5193 -1648
rect -5385 -1688 -5193 -1682
rect -5127 -1648 -4935 -1642
rect -5127 -1682 -5115 -1648
rect -4947 -1682 -4935 -1648
rect -5127 -1688 -4935 -1682
rect -4869 -1648 -4677 -1642
rect -4869 -1682 -4857 -1648
rect -4689 -1682 -4677 -1648
rect -4869 -1688 -4677 -1682
rect -4611 -1648 -4419 -1642
rect -4611 -1682 -4599 -1648
rect -4431 -1682 -4419 -1648
rect -4611 -1688 -4419 -1682
rect -4353 -1648 -4161 -1642
rect -4353 -1682 -4341 -1648
rect -4173 -1682 -4161 -1648
rect -4353 -1688 -4161 -1682
rect -4095 -1648 -3903 -1642
rect -4095 -1682 -4083 -1648
rect -3915 -1682 -3903 -1648
rect -4095 -1688 -3903 -1682
rect -3837 -1648 -3645 -1642
rect -3837 -1682 -3825 -1648
rect -3657 -1682 -3645 -1648
rect -3837 -1688 -3645 -1682
rect -3579 -1648 -3387 -1642
rect -3579 -1682 -3567 -1648
rect -3399 -1682 -3387 -1648
rect -3579 -1688 -3387 -1682
rect -3321 -1648 -3129 -1642
rect -3321 -1682 -3309 -1648
rect -3141 -1682 -3129 -1648
rect -3321 -1688 -3129 -1682
rect -3063 -1648 -2871 -1642
rect -3063 -1682 -3051 -1648
rect -2883 -1682 -2871 -1648
rect -3063 -1688 -2871 -1682
rect -2805 -1648 -2613 -1642
rect -2805 -1682 -2793 -1648
rect -2625 -1682 -2613 -1648
rect -2805 -1688 -2613 -1682
rect -2547 -1648 -2355 -1642
rect -2547 -1682 -2535 -1648
rect -2367 -1682 -2355 -1648
rect -2547 -1688 -2355 -1682
rect -2289 -1648 -2097 -1642
rect -2289 -1682 -2277 -1648
rect -2109 -1682 -2097 -1648
rect -2289 -1688 -2097 -1682
rect -2031 -1648 -1839 -1642
rect -2031 -1682 -2019 -1648
rect -1851 -1682 -1839 -1648
rect -2031 -1688 -1839 -1682
rect -1773 -1648 -1581 -1642
rect -1773 -1682 -1761 -1648
rect -1593 -1682 -1581 -1648
rect -1773 -1688 -1581 -1682
rect -1515 -1648 -1323 -1642
rect -1515 -1682 -1503 -1648
rect -1335 -1682 -1323 -1648
rect -1515 -1688 -1323 -1682
rect -1257 -1648 -1065 -1642
rect -1257 -1682 -1245 -1648
rect -1077 -1682 -1065 -1648
rect -1257 -1688 -1065 -1682
rect -999 -1648 -807 -1642
rect -999 -1682 -987 -1648
rect -819 -1682 -807 -1648
rect -999 -1688 -807 -1682
rect -741 -1648 -549 -1642
rect -741 -1682 -729 -1648
rect -561 -1682 -549 -1648
rect -741 -1688 -549 -1682
rect -483 -1648 -291 -1642
rect -483 -1682 -471 -1648
rect -303 -1682 -291 -1648
rect -483 -1688 -291 -1682
rect -225 -1648 -33 -1642
rect -225 -1682 -213 -1648
rect -45 -1682 -33 -1648
rect -225 -1688 -33 -1682
rect 33 -1648 225 -1642
rect 33 -1682 45 -1648
rect 213 -1682 225 -1648
rect 33 -1688 225 -1682
rect 291 -1648 483 -1642
rect 291 -1682 303 -1648
rect 471 -1682 483 -1648
rect 291 -1688 483 -1682
rect 549 -1648 741 -1642
rect 549 -1682 561 -1648
rect 729 -1682 741 -1648
rect 549 -1688 741 -1682
rect 807 -1648 999 -1642
rect 807 -1682 819 -1648
rect 987 -1682 999 -1648
rect 807 -1688 999 -1682
rect 1065 -1648 1257 -1642
rect 1065 -1682 1077 -1648
rect 1245 -1682 1257 -1648
rect 1065 -1688 1257 -1682
rect 1323 -1648 1515 -1642
rect 1323 -1682 1335 -1648
rect 1503 -1682 1515 -1648
rect 1323 -1688 1515 -1682
rect 1581 -1648 1773 -1642
rect 1581 -1682 1593 -1648
rect 1761 -1682 1773 -1648
rect 1581 -1688 1773 -1682
rect 1839 -1648 2031 -1642
rect 1839 -1682 1851 -1648
rect 2019 -1682 2031 -1648
rect 1839 -1688 2031 -1682
rect 2097 -1648 2289 -1642
rect 2097 -1682 2109 -1648
rect 2277 -1682 2289 -1648
rect 2097 -1688 2289 -1682
rect 2355 -1648 2547 -1642
rect 2355 -1682 2367 -1648
rect 2535 -1682 2547 -1648
rect 2355 -1688 2547 -1682
rect 2613 -1648 2805 -1642
rect 2613 -1682 2625 -1648
rect 2793 -1682 2805 -1648
rect 2613 -1688 2805 -1682
rect 2871 -1648 3063 -1642
rect 2871 -1682 2883 -1648
rect 3051 -1682 3063 -1648
rect 2871 -1688 3063 -1682
rect 3129 -1648 3321 -1642
rect 3129 -1682 3141 -1648
rect 3309 -1682 3321 -1648
rect 3129 -1688 3321 -1682
rect 3387 -1648 3579 -1642
rect 3387 -1682 3399 -1648
rect 3567 -1682 3579 -1648
rect 3387 -1688 3579 -1682
rect 3645 -1648 3837 -1642
rect 3645 -1682 3657 -1648
rect 3825 -1682 3837 -1648
rect 3645 -1688 3837 -1682
rect 3903 -1648 4095 -1642
rect 3903 -1682 3915 -1648
rect 4083 -1682 4095 -1648
rect 3903 -1688 4095 -1682
rect 4161 -1648 4353 -1642
rect 4161 -1682 4173 -1648
rect 4341 -1682 4353 -1648
rect 4161 -1688 4353 -1682
rect 4419 -1648 4611 -1642
rect 4419 -1682 4431 -1648
rect 4599 -1682 4611 -1648
rect 4419 -1688 4611 -1682
rect 4677 -1648 4869 -1642
rect 4677 -1682 4689 -1648
rect 4857 -1682 4869 -1648
rect 4677 -1688 4869 -1682
rect 4935 -1648 5127 -1642
rect 4935 -1682 4947 -1648
rect 5115 -1682 5127 -1648
rect 4935 -1688 5127 -1682
rect 5193 -1648 5385 -1642
rect 5193 -1682 5205 -1648
rect 5373 -1682 5385 -1648
rect 5193 -1688 5385 -1682
rect 5451 -1648 5643 -1642
rect 5451 -1682 5463 -1648
rect 5631 -1682 5643 -1648
rect 5451 -1688 5643 -1682
rect -5699 -1732 -5653 -1720
rect -5699 -2708 -5693 -1732
rect -5659 -2708 -5653 -1732
rect -5699 -2720 -5653 -2708
rect -5441 -1732 -5395 -1720
rect -5441 -2708 -5435 -1732
rect -5401 -2708 -5395 -1732
rect -5441 -2720 -5395 -2708
rect -5183 -1732 -5137 -1720
rect -5183 -2708 -5177 -1732
rect -5143 -2708 -5137 -1732
rect -5183 -2720 -5137 -2708
rect -4925 -1732 -4879 -1720
rect -4925 -2708 -4919 -1732
rect -4885 -2708 -4879 -1732
rect -4925 -2720 -4879 -2708
rect -4667 -1732 -4621 -1720
rect -4667 -2708 -4661 -1732
rect -4627 -2708 -4621 -1732
rect -4667 -2720 -4621 -2708
rect -4409 -1732 -4363 -1720
rect -4409 -2708 -4403 -1732
rect -4369 -2708 -4363 -1732
rect -4409 -2720 -4363 -2708
rect -4151 -1732 -4105 -1720
rect -4151 -2708 -4145 -1732
rect -4111 -2708 -4105 -1732
rect -4151 -2720 -4105 -2708
rect -3893 -1732 -3847 -1720
rect -3893 -2708 -3887 -1732
rect -3853 -2708 -3847 -1732
rect -3893 -2720 -3847 -2708
rect -3635 -1732 -3589 -1720
rect -3635 -2708 -3629 -1732
rect -3595 -2708 -3589 -1732
rect -3635 -2720 -3589 -2708
rect -3377 -1732 -3331 -1720
rect -3377 -2708 -3371 -1732
rect -3337 -2708 -3331 -1732
rect -3377 -2720 -3331 -2708
rect -3119 -1732 -3073 -1720
rect -3119 -2708 -3113 -1732
rect -3079 -2708 -3073 -1732
rect -3119 -2720 -3073 -2708
rect -2861 -1732 -2815 -1720
rect -2861 -2708 -2855 -1732
rect -2821 -2708 -2815 -1732
rect -2861 -2720 -2815 -2708
rect -2603 -1732 -2557 -1720
rect -2603 -2708 -2597 -1732
rect -2563 -2708 -2557 -1732
rect -2603 -2720 -2557 -2708
rect -2345 -1732 -2299 -1720
rect -2345 -2708 -2339 -1732
rect -2305 -2708 -2299 -1732
rect -2345 -2720 -2299 -2708
rect -2087 -1732 -2041 -1720
rect -2087 -2708 -2081 -1732
rect -2047 -2708 -2041 -1732
rect -2087 -2720 -2041 -2708
rect -1829 -1732 -1783 -1720
rect -1829 -2708 -1823 -1732
rect -1789 -2708 -1783 -1732
rect -1829 -2720 -1783 -2708
rect -1571 -1732 -1525 -1720
rect -1571 -2708 -1565 -1732
rect -1531 -2708 -1525 -1732
rect -1571 -2720 -1525 -2708
rect -1313 -1732 -1267 -1720
rect -1313 -2708 -1307 -1732
rect -1273 -2708 -1267 -1732
rect -1313 -2720 -1267 -2708
rect -1055 -1732 -1009 -1720
rect -1055 -2708 -1049 -1732
rect -1015 -2708 -1009 -1732
rect -1055 -2720 -1009 -2708
rect -797 -1732 -751 -1720
rect -797 -2708 -791 -1732
rect -757 -2708 -751 -1732
rect -797 -2720 -751 -2708
rect -539 -1732 -493 -1720
rect -539 -2708 -533 -1732
rect -499 -2708 -493 -1732
rect -539 -2720 -493 -2708
rect -281 -1732 -235 -1720
rect -281 -2708 -275 -1732
rect -241 -2708 -235 -1732
rect -281 -2720 -235 -2708
rect -23 -1732 23 -1720
rect -23 -2708 -17 -1732
rect 17 -2708 23 -1732
rect -23 -2720 23 -2708
rect 235 -1732 281 -1720
rect 235 -2708 241 -1732
rect 275 -2708 281 -1732
rect 235 -2720 281 -2708
rect 493 -1732 539 -1720
rect 493 -2708 499 -1732
rect 533 -2708 539 -1732
rect 493 -2720 539 -2708
rect 751 -1732 797 -1720
rect 751 -2708 757 -1732
rect 791 -2708 797 -1732
rect 751 -2720 797 -2708
rect 1009 -1732 1055 -1720
rect 1009 -2708 1015 -1732
rect 1049 -2708 1055 -1732
rect 1009 -2720 1055 -2708
rect 1267 -1732 1313 -1720
rect 1267 -2708 1273 -1732
rect 1307 -2708 1313 -1732
rect 1267 -2720 1313 -2708
rect 1525 -1732 1571 -1720
rect 1525 -2708 1531 -1732
rect 1565 -2708 1571 -1732
rect 1525 -2720 1571 -2708
rect 1783 -1732 1829 -1720
rect 1783 -2708 1789 -1732
rect 1823 -2708 1829 -1732
rect 1783 -2720 1829 -2708
rect 2041 -1732 2087 -1720
rect 2041 -2708 2047 -1732
rect 2081 -2708 2087 -1732
rect 2041 -2720 2087 -2708
rect 2299 -1732 2345 -1720
rect 2299 -2708 2305 -1732
rect 2339 -2708 2345 -1732
rect 2299 -2720 2345 -2708
rect 2557 -1732 2603 -1720
rect 2557 -2708 2563 -1732
rect 2597 -2708 2603 -1732
rect 2557 -2720 2603 -2708
rect 2815 -1732 2861 -1720
rect 2815 -2708 2821 -1732
rect 2855 -2708 2861 -1732
rect 2815 -2720 2861 -2708
rect 3073 -1732 3119 -1720
rect 3073 -2708 3079 -1732
rect 3113 -2708 3119 -1732
rect 3073 -2720 3119 -2708
rect 3331 -1732 3377 -1720
rect 3331 -2708 3337 -1732
rect 3371 -2708 3377 -1732
rect 3331 -2720 3377 -2708
rect 3589 -1732 3635 -1720
rect 3589 -2708 3595 -1732
rect 3629 -2708 3635 -1732
rect 3589 -2720 3635 -2708
rect 3847 -1732 3893 -1720
rect 3847 -2708 3853 -1732
rect 3887 -2708 3893 -1732
rect 3847 -2720 3893 -2708
rect 4105 -1732 4151 -1720
rect 4105 -2708 4111 -1732
rect 4145 -2708 4151 -1732
rect 4105 -2720 4151 -2708
rect 4363 -1732 4409 -1720
rect 4363 -2708 4369 -1732
rect 4403 -2708 4409 -1732
rect 4363 -2720 4409 -2708
rect 4621 -1732 4667 -1720
rect 4621 -2708 4627 -1732
rect 4661 -2708 4667 -1732
rect 4621 -2720 4667 -2708
rect 4879 -1732 4925 -1720
rect 4879 -2708 4885 -1732
rect 4919 -2708 4925 -1732
rect 4879 -2720 4925 -2708
rect 5137 -1732 5183 -1720
rect 5137 -2708 5143 -1732
rect 5177 -2708 5183 -1732
rect 5137 -2720 5183 -2708
rect 5395 -1732 5441 -1720
rect 5395 -2708 5401 -1732
rect 5435 -2708 5441 -1732
rect 5395 -2720 5441 -2708
rect 5653 -1732 5699 -1720
rect 5653 -2708 5659 -1732
rect 5693 -2708 5699 -1732
rect 5653 -2720 5699 -2708
rect -5643 -2758 -5451 -2752
rect -5643 -2792 -5631 -2758
rect -5463 -2792 -5451 -2758
rect -5643 -2798 -5451 -2792
rect -5385 -2758 -5193 -2752
rect -5385 -2792 -5373 -2758
rect -5205 -2792 -5193 -2758
rect -5385 -2798 -5193 -2792
rect -5127 -2758 -4935 -2752
rect -5127 -2792 -5115 -2758
rect -4947 -2792 -4935 -2758
rect -5127 -2798 -4935 -2792
rect -4869 -2758 -4677 -2752
rect -4869 -2792 -4857 -2758
rect -4689 -2792 -4677 -2758
rect -4869 -2798 -4677 -2792
rect -4611 -2758 -4419 -2752
rect -4611 -2792 -4599 -2758
rect -4431 -2792 -4419 -2758
rect -4611 -2798 -4419 -2792
rect -4353 -2758 -4161 -2752
rect -4353 -2792 -4341 -2758
rect -4173 -2792 -4161 -2758
rect -4353 -2798 -4161 -2792
rect -4095 -2758 -3903 -2752
rect -4095 -2792 -4083 -2758
rect -3915 -2792 -3903 -2758
rect -4095 -2798 -3903 -2792
rect -3837 -2758 -3645 -2752
rect -3837 -2792 -3825 -2758
rect -3657 -2792 -3645 -2758
rect -3837 -2798 -3645 -2792
rect -3579 -2758 -3387 -2752
rect -3579 -2792 -3567 -2758
rect -3399 -2792 -3387 -2758
rect -3579 -2798 -3387 -2792
rect -3321 -2758 -3129 -2752
rect -3321 -2792 -3309 -2758
rect -3141 -2792 -3129 -2758
rect -3321 -2798 -3129 -2792
rect -3063 -2758 -2871 -2752
rect -3063 -2792 -3051 -2758
rect -2883 -2792 -2871 -2758
rect -3063 -2798 -2871 -2792
rect -2805 -2758 -2613 -2752
rect -2805 -2792 -2793 -2758
rect -2625 -2792 -2613 -2758
rect -2805 -2798 -2613 -2792
rect -2547 -2758 -2355 -2752
rect -2547 -2792 -2535 -2758
rect -2367 -2792 -2355 -2758
rect -2547 -2798 -2355 -2792
rect -2289 -2758 -2097 -2752
rect -2289 -2792 -2277 -2758
rect -2109 -2792 -2097 -2758
rect -2289 -2798 -2097 -2792
rect -2031 -2758 -1839 -2752
rect -2031 -2792 -2019 -2758
rect -1851 -2792 -1839 -2758
rect -2031 -2798 -1839 -2792
rect -1773 -2758 -1581 -2752
rect -1773 -2792 -1761 -2758
rect -1593 -2792 -1581 -2758
rect -1773 -2798 -1581 -2792
rect -1515 -2758 -1323 -2752
rect -1515 -2792 -1503 -2758
rect -1335 -2792 -1323 -2758
rect -1515 -2798 -1323 -2792
rect -1257 -2758 -1065 -2752
rect -1257 -2792 -1245 -2758
rect -1077 -2792 -1065 -2758
rect -1257 -2798 -1065 -2792
rect -999 -2758 -807 -2752
rect -999 -2792 -987 -2758
rect -819 -2792 -807 -2758
rect -999 -2798 -807 -2792
rect -741 -2758 -549 -2752
rect -741 -2792 -729 -2758
rect -561 -2792 -549 -2758
rect -741 -2798 -549 -2792
rect -483 -2758 -291 -2752
rect -483 -2792 -471 -2758
rect -303 -2792 -291 -2758
rect -483 -2798 -291 -2792
rect -225 -2758 -33 -2752
rect -225 -2792 -213 -2758
rect -45 -2792 -33 -2758
rect -225 -2798 -33 -2792
rect 33 -2758 225 -2752
rect 33 -2792 45 -2758
rect 213 -2792 225 -2758
rect 33 -2798 225 -2792
rect 291 -2758 483 -2752
rect 291 -2792 303 -2758
rect 471 -2792 483 -2758
rect 291 -2798 483 -2792
rect 549 -2758 741 -2752
rect 549 -2792 561 -2758
rect 729 -2792 741 -2758
rect 549 -2798 741 -2792
rect 807 -2758 999 -2752
rect 807 -2792 819 -2758
rect 987 -2792 999 -2758
rect 807 -2798 999 -2792
rect 1065 -2758 1257 -2752
rect 1065 -2792 1077 -2758
rect 1245 -2792 1257 -2758
rect 1065 -2798 1257 -2792
rect 1323 -2758 1515 -2752
rect 1323 -2792 1335 -2758
rect 1503 -2792 1515 -2758
rect 1323 -2798 1515 -2792
rect 1581 -2758 1773 -2752
rect 1581 -2792 1593 -2758
rect 1761 -2792 1773 -2758
rect 1581 -2798 1773 -2792
rect 1839 -2758 2031 -2752
rect 1839 -2792 1851 -2758
rect 2019 -2792 2031 -2758
rect 1839 -2798 2031 -2792
rect 2097 -2758 2289 -2752
rect 2097 -2792 2109 -2758
rect 2277 -2792 2289 -2758
rect 2097 -2798 2289 -2792
rect 2355 -2758 2547 -2752
rect 2355 -2792 2367 -2758
rect 2535 -2792 2547 -2758
rect 2355 -2798 2547 -2792
rect 2613 -2758 2805 -2752
rect 2613 -2792 2625 -2758
rect 2793 -2792 2805 -2758
rect 2613 -2798 2805 -2792
rect 2871 -2758 3063 -2752
rect 2871 -2792 2883 -2758
rect 3051 -2792 3063 -2758
rect 2871 -2798 3063 -2792
rect 3129 -2758 3321 -2752
rect 3129 -2792 3141 -2758
rect 3309 -2792 3321 -2758
rect 3129 -2798 3321 -2792
rect 3387 -2758 3579 -2752
rect 3387 -2792 3399 -2758
rect 3567 -2792 3579 -2758
rect 3387 -2798 3579 -2792
rect 3645 -2758 3837 -2752
rect 3645 -2792 3657 -2758
rect 3825 -2792 3837 -2758
rect 3645 -2798 3837 -2792
rect 3903 -2758 4095 -2752
rect 3903 -2792 3915 -2758
rect 4083 -2792 4095 -2758
rect 3903 -2798 4095 -2792
rect 4161 -2758 4353 -2752
rect 4161 -2792 4173 -2758
rect 4341 -2792 4353 -2758
rect 4161 -2798 4353 -2792
rect 4419 -2758 4611 -2752
rect 4419 -2792 4431 -2758
rect 4599 -2792 4611 -2758
rect 4419 -2798 4611 -2792
rect 4677 -2758 4869 -2752
rect 4677 -2792 4689 -2758
rect 4857 -2792 4869 -2758
rect 4677 -2798 4869 -2792
rect 4935 -2758 5127 -2752
rect 4935 -2792 4947 -2758
rect 5115 -2792 5127 -2758
rect 4935 -2798 5127 -2792
rect 5193 -2758 5385 -2752
rect 5193 -2792 5205 -2758
rect 5373 -2792 5385 -2758
rect 5193 -2798 5385 -2792
rect 5451 -2758 5643 -2752
rect 5451 -2792 5463 -2758
rect 5631 -2792 5643 -2758
rect 5451 -2798 5643 -2792
<< properties >>
string FIXED_BBOX -5810 -2913 5810 2913
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 1.0 m 5 nf 44 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
