magic
tech sky130A
magscale 1 2
timestamp 1730992408
<< dnwell >>
rect 14128 -7904 19768 -7862
rect 22482 -7904 29106 -7862
rect 14128 -35804 29106 -7904
rect 14128 -36806 29108 -35804
rect 14132 -36862 29108 -36806
rect 14132 -36866 21822 -36862
<< locali >>
rect 14880 -8006 19731 -7992
rect 14880 -8042 14988 -8006
rect 19650 -8042 19731 -8006
rect 14880 -8054 19731 -8042
rect 14880 -8130 14942 -8054
rect 14880 -12422 14894 -8130
rect 14932 -12422 14942 -8130
rect 14880 -12442 14942 -12422
rect 19669 -8134 19731 -8054
rect 19669 -13042 19682 -8134
rect 19716 -13034 19731 -8134
rect 19716 -13042 19936 -13034
rect 19669 -13075 19936 -13042
rect 19670 -13076 19936 -13075
rect 15434 -18237 24321 -18236
rect 15433 -18250 24321 -18237
rect 15433 -18256 15984 -18250
rect 15433 -22834 15450 -18256
rect 15502 -18300 15984 -18256
rect 24202 -18260 24321 -18250
rect 24202 -18300 24254 -18260
rect 15502 -18318 24254 -18300
rect 15502 -22775 15515 -18318
rect 24239 -22775 24254 -18318
rect 15502 -22794 24254 -22775
rect 15502 -22834 16104 -22794
rect 15433 -22840 16104 -22834
rect 23956 -22828 24254 -22794
rect 24304 -22828 24321 -18260
rect 23956 -22840 24321 -22828
rect 15433 -22857 24321 -22840
rect 15426 -27926 24362 -27910
rect 15426 -27946 16050 -27926
rect 15426 -32362 15458 -27946
rect 15520 -27992 16050 -27946
rect 24232 -27992 24362 -27926
rect 15520 -28010 24362 -27992
rect 15520 -32362 15526 -28010
rect 15426 -32490 15526 -32362
rect 24262 -28032 24362 -28010
rect 24262 -32490 24280 -28032
rect 24346 -32490 24362 -28032
rect 15426 -32496 24362 -32490
rect 15426 -32572 16192 -32496
rect 23938 -32572 24362 -32496
rect 15426 -32590 24362 -32572
<< viali >>
rect 14988 -8042 19650 -8006
rect 14894 -12422 14932 -8130
rect 19682 -13042 19716 -8134
rect 15450 -22834 15502 -18256
rect 15984 -18300 24202 -18250
rect 16104 -22840 23956 -22794
rect 24254 -22828 24304 -18260
rect 15458 -32362 15520 -27946
rect 16050 -27992 24232 -27926
rect 24280 -32490 24346 -28032
rect 16192 -32572 23938 -32496
<< metal1 >>
rect 14880 -8002 19731 -7992
rect 14880 -8058 14956 -8002
rect 19662 -8058 19731 -8002
rect 14880 -8076 19731 -8058
rect 14880 -8130 14942 -8076
rect 14880 -12422 14894 -8130
rect 14932 -12422 14942 -8130
rect 19669 -8134 19731 -8076
rect 26526 -8124 26726 -7924
rect 15030 -8586 15266 -8154
rect 15362 -8586 15598 -8154
rect 15694 -8586 15930 -8154
rect 16026 -8586 16262 -8154
rect 16358 -8586 16594 -8154
rect 16690 -8586 16926 -8154
rect 17022 -8586 17258 -8154
rect 17354 -8586 17590 -8154
rect 17686 -8586 17922 -8154
rect 18018 -8586 18254 -8154
rect 18350 -8586 18586 -8154
rect 18682 -8586 18918 -8154
rect 19014 -8586 19250 -8154
rect 19346 -8586 19582 -8154
rect 14880 -12442 14942 -12422
rect 14672 -12522 15100 -12514
rect 14672 -12938 14682 -12522
rect 14874 -12938 15100 -12522
rect 14672 -12946 15100 -12938
rect 15196 -12946 15434 -12514
rect 15528 -12946 15766 -12514
rect 15860 -12946 16098 -12514
rect 16192 -12946 16430 -12514
rect 16524 -12946 16762 -12514
rect 16856 -12946 17094 -12514
rect 17188 -13326 17258 -12916
rect 14682 -13406 17258 -13326
rect 14566 -13948 14642 -13939
rect 14566 -17574 14642 -14146
rect 14682 -17392 14758 -13406
rect 17354 -13486 17424 -12896
rect 17520 -12946 17758 -12514
rect 17852 -12946 18090 -12514
rect 18184 -12946 18422 -12514
rect 18516 -12946 18754 -12514
rect 18848 -12946 19086 -12514
rect 19180 -12946 19418 -12514
rect 14954 -13566 17424 -13486
rect 14954 -13948 15034 -13566
rect 19512 -13925 19582 -12890
rect 19669 -13042 19682 -8134
rect 19716 -13034 19731 -8134
rect 19716 -13042 19936 -13034
rect 19669 -13075 19936 -13042
rect 19670 -13076 19936 -13075
rect 19511 -13991 25752 -13925
rect 14954 -14156 15034 -14146
rect 25686 -14682 25752 -13991
rect 25481 -14748 25752 -14682
rect 21738 -17392 21940 -17316
rect 14682 -17400 15584 -17392
rect 14682 -17496 14692 -17400
rect 15572 -17496 15584 -17400
rect 14682 -17502 15584 -17496
rect 14566 -17582 15064 -17574
rect 14566 -17680 14574 -17582
rect 15050 -17680 15064 -17582
rect 14566 -17690 15064 -17680
rect 15103 -23667 15165 -17502
rect 21738 -17528 21940 -17502
rect 15224 -17582 15584 -17572
rect 15224 -17684 15236 -17582
rect 15572 -17684 15584 -17582
rect 15224 -17692 15584 -17684
rect 14554 -23729 15165 -23667
rect 15238 -22904 15330 -17692
rect 15390 -17756 15686 -17746
rect 15390 -17842 15402 -17756
rect 15676 -17842 15686 -17756
rect 15390 -17854 15686 -17842
rect 15766 -17758 16062 -17746
rect 15766 -17844 15778 -17758
rect 16052 -17844 16062 -17758
rect 15766 -17854 16062 -17844
rect 22302 -17756 22502 -17316
rect 26526 -17701 26592 -17249
rect 15430 -18250 15516 -18236
rect 15430 -18372 15434 -18250
rect 15510 -18372 15516 -18250
rect 15430 -22834 15450 -18372
rect 15502 -22834 15516 -18372
rect 15606 -18844 15676 -17854
rect 15772 -18842 15842 -17854
rect 22302 -17878 22502 -17844
rect 15930 -18242 24321 -18236
rect 15930 -18306 15954 -18242
rect 24266 -18260 24321 -18242
rect 15930 -18318 24254 -18306
rect 15936 -18840 16172 -18408
rect 16268 -18840 16504 -18408
rect 16600 -18840 16836 -18408
rect 16932 -18840 17168 -18408
rect 17264 -18840 17500 -18408
rect 17596 -18840 17832 -18408
rect 17928 -18840 18164 -18408
rect 18260 -18840 18496 -18408
rect 18592 -18840 18828 -18408
rect 18924 -18840 19160 -18408
rect 19256 -18840 19492 -18408
rect 19588 -18840 19824 -18408
rect 19920 -18840 20156 -18408
rect 20252 -18840 20488 -18408
rect 20584 -18840 20820 -18408
rect 20916 -18840 21152 -18408
rect 21248 -18840 21484 -18408
rect 21580 -18840 21816 -18408
rect 21912 -18840 22148 -18408
rect 22244 -18840 22480 -18408
rect 22576 -18840 22812 -18408
rect 22908 -18840 23144 -18408
rect 23240 -18840 23476 -18408
rect 23572 -18840 23808 -18408
rect 23904 -18840 24140 -18408
rect 15770 -22260 15842 -22258
rect 15606 -22692 15842 -22260
rect 15430 -22858 15516 -22834
rect 15938 -22904 16012 -22258
rect 16102 -22690 16338 -22258
rect 16434 -22690 16670 -22258
rect 16766 -22690 17002 -22258
rect 17098 -22690 17334 -22258
rect 17430 -22690 17666 -22258
rect 17762 -22690 17998 -22258
rect 18094 -22690 18330 -22258
rect 18426 -22690 18662 -22258
rect 18758 -22690 18994 -22258
rect 19090 -22690 19326 -22258
rect 19422 -22690 19658 -22258
rect 19754 -22690 19990 -22258
rect 20086 -22690 20322 -22258
rect 20418 -22690 20654 -22258
rect 20750 -22690 20986 -22258
rect 21082 -22690 21318 -22258
rect 21414 -22690 21650 -22258
rect 21746 -22690 21982 -22258
rect 22078 -22690 22314 -22258
rect 22410 -22690 22646 -22258
rect 22742 -22690 22978 -22258
rect 23074 -22690 23310 -22258
rect 23406 -22690 23642 -22258
rect 23738 -22690 23974 -22258
rect 16076 -22794 23988 -22774
rect 16076 -22840 16104 -22794
rect 23956 -22840 23988 -22794
rect 16076 -22860 23988 -22840
rect 15238 -23036 16012 -22904
rect 14554 -27132 14616 -23729
rect 15238 -23793 15330 -23036
rect 24070 -23678 24140 -22258
rect 24239 -22828 24254 -18318
rect 24304 -22828 24321 -18260
rect 24239 -22857 24321 -22828
rect 24070 -23692 25747 -23678
rect 24070 -23748 25748 -23692
rect 14672 -23863 15330 -23793
rect 14354 -27142 14618 -27132
rect 14354 -27204 14366 -27142
rect 14606 -27204 14618 -27142
rect 14354 -27212 14618 -27204
rect 14672 -27285 14738 -23863
rect 25677 -24434 25748 -23748
rect 25438 -24490 25748 -24434
rect 15616 -27138 15876 -27132
rect 15616 -27206 15628 -27138
rect 15862 -27206 15876 -27138
rect 15616 -27214 15876 -27206
rect 22294 -27190 22494 -27064
rect 14672 -27351 15353 -27285
rect 14672 -27352 14738 -27351
rect 15287 -32486 15353 -27351
rect 15452 -27494 15712 -27488
rect 15452 -27562 15466 -27494
rect 15700 -27562 15712 -27494
rect 15452 -27570 15712 -27562
rect 15424 -27946 15542 -27910
rect 15424 -32362 15458 -27946
rect 15520 -32362 15542 -27946
rect 15634 -28132 15704 -27570
rect 15802 -28558 15870 -27214
rect 22294 -27292 22494 -27286
rect 26518 -27407 26584 -26999
rect 16000 -27916 24362 -27910
rect 16000 -27926 16082 -27916
rect 24200 -27926 24362 -27916
rect 16000 -27992 16050 -27926
rect 24232 -27992 24362 -27926
rect 16000 -28004 16082 -27992
rect 24200 -28004 24362 -27992
rect 16000 -28010 24362 -28004
rect 24262 -28032 24362 -28010
rect 15966 -28558 16202 -28126
rect 16298 -28558 16534 -28126
rect 16630 -28558 16866 -28126
rect 16962 -28558 17198 -28126
rect 17294 -28558 17530 -28126
rect 17626 -28558 17862 -28126
rect 17958 -28558 18194 -28126
rect 18290 -28558 18526 -28126
rect 18622 -28558 18858 -28126
rect 18954 -28558 19190 -28126
rect 19286 -28558 19522 -28126
rect 19618 -28558 19854 -28126
rect 19950 -28558 20186 -28126
rect 20282 -28558 20518 -28126
rect 20614 -28558 20850 -28126
rect 20946 -28558 21182 -28126
rect 21278 -28558 21514 -28126
rect 21610 -28558 21846 -28126
rect 21942 -28558 22178 -28126
rect 22274 -28558 22510 -28126
rect 22606 -28558 22842 -28126
rect 22938 -28558 23174 -28126
rect 23270 -28558 23506 -28126
rect 23602 -28558 23838 -28126
rect 23934 -28558 24170 -28126
rect 15424 -32400 15542 -32362
rect 15634 -32408 15870 -31976
rect 15966 -32486 16038 -31974
rect 16132 -32408 16368 -31976
rect 16464 -32408 16700 -31976
rect 16796 -32408 17032 -31976
rect 17128 -32408 17364 -31976
rect 17460 -32408 17696 -31976
rect 17792 -32408 18028 -31976
rect 18124 -32408 18360 -31976
rect 18456 -32408 18692 -31976
rect 18788 -32408 19024 -31976
rect 19120 -32408 19356 -31976
rect 19452 -32408 19688 -31976
rect 19784 -32408 20020 -31976
rect 20116 -32408 20352 -31976
rect 20448 -32408 20684 -31976
rect 20780 -32408 21016 -31976
rect 21112 -32408 21348 -31976
rect 21444 -32408 21680 -31976
rect 21776 -32408 22012 -31976
rect 22108 -32408 22344 -31976
rect 22440 -32408 22676 -31976
rect 22772 -32408 23008 -31976
rect 23104 -32408 23340 -31976
rect 23436 -32408 23672 -31976
rect 23768 -32408 24004 -31976
rect 15287 -32549 16038 -32486
rect 15288 -32580 16038 -32549
rect 16156 -32496 23994 -32484
rect 16156 -32572 16192 -32496
rect 23938 -32572 23994 -32496
rect 16156 -32594 23994 -32572
rect 24096 -33380 24174 -31970
rect 24262 -32490 24280 -28032
rect 24346 -32490 24362 -28032
rect 24262 -32534 24362 -32490
rect 24096 -33459 25728 -33380
rect 25649 -34154 25728 -33459
rect 25444 -34210 25728 -34154
rect 22294 -36876 22494 -36784
rect 22286 -36978 22294 -36876
rect 22494 -36978 22502 -36876
<< via1 >>
rect 14956 -8006 19662 -8002
rect 14956 -8042 14988 -8006
rect 14988 -8042 19650 -8006
rect 19650 -8042 19662 -8006
rect 14956 -8058 19662 -8042
rect 14682 -12938 14874 -12522
rect 14566 -14146 14642 -13948
rect 14954 -14146 15034 -13948
rect 14692 -17496 15572 -17400
rect 21738 -17502 21940 -17392
rect 14574 -17680 15050 -17582
rect 15236 -17684 15572 -17582
rect 15402 -17842 15676 -17756
rect 15778 -17844 16052 -17758
rect 22302 -17844 22502 -17756
rect 15434 -18256 15510 -18250
rect 15434 -18372 15450 -18256
rect 15450 -18372 15502 -18256
rect 15502 -18372 15510 -18256
rect 15954 -18250 24266 -18242
rect 15954 -18300 15984 -18250
rect 15984 -18300 24202 -18250
rect 24202 -18260 24266 -18250
rect 24202 -18300 24254 -18260
rect 15954 -18306 24254 -18300
rect 24254 -18306 24266 -18260
rect 14366 -27204 14606 -27142
rect 18718 -24482 19240 -24426
rect 15628 -27206 15862 -27138
rect 15466 -27562 15700 -27494
rect 22294 -27286 22494 -27190
rect 16082 -27926 24200 -27916
rect 16082 -27992 24200 -27926
rect 16082 -28004 24200 -27992
rect 18734 -34202 19360 -34146
rect 22294 -36978 22494 -36876
<< metal2 >>
rect 14864 -8002 19938 -7970
rect 14864 -8058 14956 -8002
rect 19662 -8058 19938 -8002
rect 14864 -8106 19938 -8058
rect 14672 -12522 14884 -12514
rect 14672 -12938 14682 -12522
rect 14874 -12938 14884 -12522
rect 14672 -12946 14884 -12938
rect 14509 -14146 14566 -13948
rect 14642 -14146 14954 -13948
rect 15034 -14146 15041 -13948
rect 14649 -17400 21738 -17392
rect 14649 -17496 14692 -17400
rect 15572 -17496 21738 -17400
rect 14649 -17502 21738 -17496
rect 21940 -17502 21966 -17392
rect 28948 -17500 29148 -17426
rect 14514 -17580 15064 -17574
rect 15224 -17580 15584 -17572
rect 23918 -17580 29148 -17500
rect 14514 -17582 29148 -17580
rect 14514 -17680 14574 -17582
rect 15050 -17680 15236 -17582
rect 14514 -17690 15064 -17680
rect 15224 -17684 15236 -17680
rect 15572 -17600 29148 -17582
rect 15572 -17680 24030 -17600
rect 28948 -17626 29148 -17600
rect 15572 -17684 15584 -17680
rect 15224 -17692 15584 -17684
rect 14656 -17752 14878 -17750
rect 15390 -17752 15686 -17746
rect 14656 -17756 15686 -17752
rect 14656 -17758 15402 -17756
rect 14656 -17994 14674 -17758
rect 14868 -17840 15402 -17758
rect 14868 -17994 14878 -17840
rect 15390 -17842 15402 -17840
rect 15676 -17842 15686 -17756
rect 15390 -17854 15686 -17842
rect 15766 -17756 16062 -17746
rect 15766 -17758 22302 -17756
rect 15766 -17844 15778 -17758
rect 16052 -17844 22302 -17758
rect 22502 -17844 22536 -17756
rect 15766 -17854 16062 -17844
rect 14656 -18002 14878 -17994
rect 15398 -18242 24516 -18004
rect 15398 -18250 15954 -18242
rect 15398 -18372 15434 -18250
rect 15510 -18306 15954 -18250
rect 24266 -18306 24516 -18242
rect 15510 -18372 24516 -18306
rect 15398 -18398 24516 -18372
rect 16594 -24190 19240 -23976
rect 18718 -24426 19240 -24190
rect 18718 -24488 19240 -24482
rect 14354 -27138 15876 -27132
rect 14354 -27142 15628 -27138
rect 14354 -27204 14366 -27142
rect 14606 -27204 15628 -27142
rect 14354 -27206 15628 -27204
rect 15862 -27206 15876 -27138
rect 28890 -27190 29090 -27150
rect 14354 -27212 15876 -27206
rect 15616 -27214 15876 -27212
rect 22286 -27286 22294 -27190
rect 22494 -27286 29090 -27190
rect 28890 -27350 29090 -27286
rect 14656 -27466 14886 -27452
rect 14656 -27608 14676 -27466
rect 14868 -27488 14886 -27466
rect 14868 -27494 15714 -27488
rect 14868 -27562 15466 -27494
rect 15700 -27562 15714 -27494
rect 14868 -27570 15714 -27562
rect 14868 -27608 14886 -27570
rect 14656 -27618 14886 -27608
rect 16032 -27916 24510 -27418
rect 16032 -28004 16082 -27916
rect 24200 -28004 24510 -27916
rect 16032 -28118 24510 -28004
rect 16600 -33910 19360 -33722
rect 18734 -34146 19360 -33910
rect 18734 -34210 19360 -34202
rect 28882 -36876 29082 -36844
rect 22286 -36978 22294 -36876
rect 22494 -36978 29082 -36876
rect 22294 -37004 29082 -36978
rect 28882 -37044 29082 -37004
<< via2 >>
rect 14682 -12938 14874 -12522
rect 14674 -17994 14868 -17758
rect 14676 -27608 14868 -27466
<< metal3 >>
rect 14672 -8786 14884 -7866
rect 28626 -8204 28826 -8004
rect 26794 -9158 26994 -8958
rect 26734 -17692 27004 -16094
rect 28458 -17696 28958 -17320
rect 14664 -17758 14876 -17752
rect 14664 -17994 14674 -17758
rect 14868 -17994 14876 -17758
rect 14664 -18524 14876 -17994
rect 26726 -27410 26996 -25842
rect 28458 -27418 28958 -27068
rect 14664 -27466 14876 -27458
rect 14664 -27608 14676 -27466
rect 14868 -27608 14876 -27466
rect 14664 -28248 14876 -27608
<< comment >>
rect 17292 -13064 17322 -8044
use sky130_fd_pr__res_xhigh_po_0p35_QHQRGL  sky130_fd_pr__res_xhigh_po_0p35_QHQRGL_0 paramcells
timestamp 1730992408
transform 1 0 17306 0 1 -10550
box -2442 -2562 2442 2562
use sky130_fd_pr__res_xhigh_po_0p35_TVN32V  sky130_fd_pr__res_xhigh_po_0p35_TVN32V_0 paramcells
timestamp 1730992408
transform 1 0 19874 0 1 -20551
box -4434 -2307 4434 2307
use sky130_fd_pr__res_xhigh_po_0p35_TVN32V  sky130_fd_pr__res_xhigh_po_0p35_TVN32V_1
timestamp 1730992408
transform 1 0 19902 0 1 -30267
box -4434 -2307 4434 2307
use Input_Stage_OA1  x1
timestamp 1730992408
transform 1 0 14036 0 1 -35700
box 628 -1154 15010 8321
use Input_Stage_OA1  x2
timestamp 1730992408
transform 1 0 14036 0 1 -25980
box 628 -1154 15010 8321
use Input_Stage_OA2  x3
timestamp 1730992408
transform 1 0 14044 0 1 -16232
box 628 -1154 15010 8321
<< labels >>
flabel metal2 28882 -37044 29082 -36844 0 FreeSans 256 90 0 0 VINN
port 3 nsew
flabel metal2 28890 -27350 29090 -27150 0 FreeSans 256 90 0 0 VINP
port 1 nsew
flabel metal2 28948 -17626 29148 -17426 0 FreeSans 256 90 0 0 CM
port 4 nsew
flabel metal3 14678 -8072 14878 -7872 0 FreeSans 256 90 0 0 VOUT1
port 2 nsew
flabel metal1 26526 -8124 26726 -7924 0 FreeSans 256 0 0 0 VBIAS
port 6 nsew
flabel metal3 26794 -9158 26994 -8958 0 FreeSans 256 90 0 0 AVSS
port 5 nsew
flabel metal3 28626 -8204 28826 -8004 0 FreeSans 256 90 0 0 AVDD
port 0 nsew
<< end >>
