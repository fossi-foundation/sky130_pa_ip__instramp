magic
tech sky130A
magscale 1 2
timestamp 1729620069
<< pwell >>
rect -3043 -2182 3043 2182
<< psubdiff >>
rect -3007 2112 -2911 2146
rect 2911 2112 3007 2146
rect -3007 2050 -2973 2112
rect 2973 2050 3007 2112
rect -3007 -2112 -2973 -2050
rect 2973 -2112 3007 -2050
rect -3007 -2146 -2911 -2112
rect 2911 -2146 3007 -2112
<< psubdiffcont >>
rect -2911 2112 2911 2146
rect -3007 -2050 -2973 2050
rect 2973 -2050 3007 2050
rect -2911 -2146 2911 -2112
<< xpolycontact >>
rect -2877 1584 -2739 2016
rect -2877 -2016 -2739 -1584
rect -2643 1584 -2505 2016
rect -2643 -2016 -2505 -1584
rect -2409 1584 -2271 2016
rect -2409 -2016 -2271 -1584
rect -2175 1584 -2037 2016
rect -2175 -2016 -2037 -1584
rect -1941 1584 -1803 2016
rect -1941 -2016 -1803 -1584
rect -1707 1584 -1569 2016
rect -1707 -2016 -1569 -1584
rect -1473 1584 -1335 2016
rect -1473 -2016 -1335 -1584
rect -1239 1584 -1101 2016
rect -1239 -2016 -1101 -1584
rect -1005 1584 -867 2016
rect -1005 -2016 -867 -1584
rect -771 1584 -633 2016
rect -771 -2016 -633 -1584
rect -537 1584 -399 2016
rect -537 -2016 -399 -1584
rect -303 1584 -165 2016
rect -303 -2016 -165 -1584
rect -69 1584 69 2016
rect -69 -2016 69 -1584
rect 165 1584 303 2016
rect 165 -2016 303 -1584
rect 399 1584 537 2016
rect 399 -2016 537 -1584
rect 633 1584 771 2016
rect 633 -2016 771 -1584
rect 867 1584 1005 2016
rect 867 -2016 1005 -1584
rect 1101 1584 1239 2016
rect 1101 -2016 1239 -1584
rect 1335 1584 1473 2016
rect 1335 -2016 1473 -1584
rect 1569 1584 1707 2016
rect 1569 -2016 1707 -1584
rect 1803 1584 1941 2016
rect 1803 -2016 1941 -1584
rect 2037 1584 2175 2016
rect 2037 -2016 2175 -1584
rect 2271 1584 2409 2016
rect 2271 -2016 2409 -1584
rect 2505 1584 2643 2016
rect 2505 -2016 2643 -1584
rect 2739 1584 2877 2016
rect 2739 -2016 2877 -1584
<< ppolyres >>
rect -2877 -1584 -2739 1584
rect -2643 -1584 -2505 1584
rect -2409 -1584 -2271 1584
rect -2175 -1584 -2037 1584
rect -1941 -1584 -1803 1584
rect -1707 -1584 -1569 1584
rect -1473 -1584 -1335 1584
rect -1239 -1584 -1101 1584
rect -1005 -1584 -867 1584
rect -771 -1584 -633 1584
rect -537 -1584 -399 1584
rect -303 -1584 -165 1584
rect -69 -1584 69 1584
rect 165 -1584 303 1584
rect 399 -1584 537 1584
rect 633 -1584 771 1584
rect 867 -1584 1005 1584
rect 1101 -1584 1239 1584
rect 1335 -1584 1473 1584
rect 1569 -1584 1707 1584
rect 1803 -1584 1941 1584
rect 2037 -1584 2175 1584
rect 2271 -1584 2409 1584
rect 2505 -1584 2643 1584
rect 2739 -1584 2877 1584
<< locali >>
rect -3007 2112 -2911 2146
rect 2911 2112 3007 2146
rect -3007 2050 -2973 2112
rect 2973 2050 3007 2112
rect -3007 -2112 -2973 -2050
rect 2973 -2112 3007 -2050
rect -3007 -2146 -2911 -2112
rect 2911 -2146 3007 -2112
<< viali >>
rect -2861 1601 -2755 1998
rect -2627 1601 -2521 1998
rect -2393 1601 -2287 1998
rect -2159 1601 -2053 1998
rect -1925 1601 -1819 1998
rect -1691 1601 -1585 1998
rect -1457 1601 -1351 1998
rect -1223 1601 -1117 1998
rect -989 1601 -883 1998
rect -755 1601 -649 1998
rect -521 1601 -415 1998
rect -287 1601 -181 1998
rect -53 1601 53 1998
rect 181 1601 287 1998
rect 415 1601 521 1998
rect 649 1601 755 1998
rect 883 1601 989 1998
rect 1117 1601 1223 1998
rect 1351 1601 1457 1998
rect 1585 1601 1691 1998
rect 1819 1601 1925 1998
rect 2053 1601 2159 1998
rect 2287 1601 2393 1998
rect 2521 1601 2627 1998
rect 2755 1601 2861 1998
rect -2861 -1998 -2755 -1601
rect -2627 -1998 -2521 -1601
rect -2393 -1998 -2287 -1601
rect -2159 -1998 -2053 -1601
rect -1925 -1998 -1819 -1601
rect -1691 -1998 -1585 -1601
rect -1457 -1998 -1351 -1601
rect -1223 -1998 -1117 -1601
rect -989 -1998 -883 -1601
rect -755 -1998 -649 -1601
rect -521 -1998 -415 -1601
rect -287 -1998 -181 -1601
rect -53 -1998 53 -1601
rect 181 -1998 287 -1601
rect 415 -1998 521 -1601
rect 649 -1998 755 -1601
rect 883 -1998 989 -1601
rect 1117 -1998 1223 -1601
rect 1351 -1998 1457 -1601
rect 1585 -1998 1691 -1601
rect 1819 -1998 1925 -1601
rect 2053 -1998 2159 -1601
rect 2287 -1998 2393 -1601
rect 2521 -1998 2627 -1601
rect 2755 -1998 2861 -1601
<< metal1 >>
rect -2867 1998 -2749 2010
rect -2867 1601 -2861 1998
rect -2755 1601 -2749 1998
rect -2867 1589 -2749 1601
rect -2633 1998 -2515 2010
rect -2633 1601 -2627 1998
rect -2521 1601 -2515 1998
rect -2633 1589 -2515 1601
rect -2399 1998 -2281 2010
rect -2399 1601 -2393 1998
rect -2287 1601 -2281 1998
rect -2399 1589 -2281 1601
rect -2165 1998 -2047 2010
rect -2165 1601 -2159 1998
rect -2053 1601 -2047 1998
rect -2165 1589 -2047 1601
rect -1931 1998 -1813 2010
rect -1931 1601 -1925 1998
rect -1819 1601 -1813 1998
rect -1931 1589 -1813 1601
rect -1697 1998 -1579 2010
rect -1697 1601 -1691 1998
rect -1585 1601 -1579 1998
rect -1697 1589 -1579 1601
rect -1463 1998 -1345 2010
rect -1463 1601 -1457 1998
rect -1351 1601 -1345 1998
rect -1463 1589 -1345 1601
rect -1229 1998 -1111 2010
rect -1229 1601 -1223 1998
rect -1117 1601 -1111 1998
rect -1229 1589 -1111 1601
rect -995 1998 -877 2010
rect -995 1601 -989 1998
rect -883 1601 -877 1998
rect -995 1589 -877 1601
rect -761 1998 -643 2010
rect -761 1601 -755 1998
rect -649 1601 -643 1998
rect -761 1589 -643 1601
rect -527 1998 -409 2010
rect -527 1601 -521 1998
rect -415 1601 -409 1998
rect -527 1589 -409 1601
rect -293 1998 -175 2010
rect -293 1601 -287 1998
rect -181 1601 -175 1998
rect -293 1589 -175 1601
rect -59 1998 59 2010
rect -59 1601 -53 1998
rect 53 1601 59 1998
rect -59 1589 59 1601
rect 175 1998 293 2010
rect 175 1601 181 1998
rect 287 1601 293 1998
rect 175 1589 293 1601
rect 409 1998 527 2010
rect 409 1601 415 1998
rect 521 1601 527 1998
rect 409 1589 527 1601
rect 643 1998 761 2010
rect 643 1601 649 1998
rect 755 1601 761 1998
rect 643 1589 761 1601
rect 877 1998 995 2010
rect 877 1601 883 1998
rect 989 1601 995 1998
rect 877 1589 995 1601
rect 1111 1998 1229 2010
rect 1111 1601 1117 1998
rect 1223 1601 1229 1998
rect 1111 1589 1229 1601
rect 1345 1998 1463 2010
rect 1345 1601 1351 1998
rect 1457 1601 1463 1998
rect 1345 1589 1463 1601
rect 1579 1998 1697 2010
rect 1579 1601 1585 1998
rect 1691 1601 1697 1998
rect 1579 1589 1697 1601
rect 1813 1998 1931 2010
rect 1813 1601 1819 1998
rect 1925 1601 1931 1998
rect 1813 1589 1931 1601
rect 2047 1998 2165 2010
rect 2047 1601 2053 1998
rect 2159 1601 2165 1998
rect 2047 1589 2165 1601
rect 2281 1998 2399 2010
rect 2281 1601 2287 1998
rect 2393 1601 2399 1998
rect 2281 1589 2399 1601
rect 2515 1998 2633 2010
rect 2515 1601 2521 1998
rect 2627 1601 2633 1998
rect 2515 1589 2633 1601
rect 2749 1998 2867 2010
rect 2749 1601 2755 1998
rect 2861 1601 2867 1998
rect 2749 1589 2867 1601
rect -2867 -1601 -2749 -1589
rect -2867 -1998 -2861 -1601
rect -2755 -1998 -2749 -1601
rect -2867 -2010 -2749 -1998
rect -2633 -1601 -2515 -1589
rect -2633 -1998 -2627 -1601
rect -2521 -1998 -2515 -1601
rect -2633 -2010 -2515 -1998
rect -2399 -1601 -2281 -1589
rect -2399 -1998 -2393 -1601
rect -2287 -1998 -2281 -1601
rect -2399 -2010 -2281 -1998
rect -2165 -1601 -2047 -1589
rect -2165 -1998 -2159 -1601
rect -2053 -1998 -2047 -1601
rect -2165 -2010 -2047 -1998
rect -1931 -1601 -1813 -1589
rect -1931 -1998 -1925 -1601
rect -1819 -1998 -1813 -1601
rect -1931 -2010 -1813 -1998
rect -1697 -1601 -1579 -1589
rect -1697 -1998 -1691 -1601
rect -1585 -1998 -1579 -1601
rect -1697 -2010 -1579 -1998
rect -1463 -1601 -1345 -1589
rect -1463 -1998 -1457 -1601
rect -1351 -1998 -1345 -1601
rect -1463 -2010 -1345 -1998
rect -1229 -1601 -1111 -1589
rect -1229 -1998 -1223 -1601
rect -1117 -1998 -1111 -1601
rect -1229 -2010 -1111 -1998
rect -995 -1601 -877 -1589
rect -995 -1998 -989 -1601
rect -883 -1998 -877 -1601
rect -995 -2010 -877 -1998
rect -761 -1601 -643 -1589
rect -761 -1998 -755 -1601
rect -649 -1998 -643 -1601
rect -761 -2010 -643 -1998
rect -527 -1601 -409 -1589
rect -527 -1998 -521 -1601
rect -415 -1998 -409 -1601
rect -527 -2010 -409 -1998
rect -293 -1601 -175 -1589
rect -293 -1998 -287 -1601
rect -181 -1998 -175 -1601
rect -293 -2010 -175 -1998
rect -59 -1601 59 -1589
rect -59 -1998 -53 -1601
rect 53 -1998 59 -1601
rect -59 -2010 59 -1998
rect 175 -1601 293 -1589
rect 175 -1998 181 -1601
rect 287 -1998 293 -1601
rect 175 -2010 293 -1998
rect 409 -1601 527 -1589
rect 409 -1998 415 -1601
rect 521 -1998 527 -1601
rect 409 -2010 527 -1998
rect 643 -1601 761 -1589
rect 643 -1998 649 -1601
rect 755 -1998 761 -1601
rect 643 -2010 761 -1998
rect 877 -1601 995 -1589
rect 877 -1998 883 -1601
rect 989 -1998 995 -1601
rect 877 -2010 995 -1998
rect 1111 -1601 1229 -1589
rect 1111 -1998 1117 -1601
rect 1223 -1998 1229 -1601
rect 1111 -2010 1229 -1998
rect 1345 -1601 1463 -1589
rect 1345 -1998 1351 -1601
rect 1457 -1998 1463 -1601
rect 1345 -2010 1463 -1998
rect 1579 -1601 1697 -1589
rect 1579 -1998 1585 -1601
rect 1691 -1998 1697 -1601
rect 1579 -2010 1697 -1998
rect 1813 -1601 1931 -1589
rect 1813 -1998 1819 -1601
rect 1925 -1998 1931 -1601
rect 1813 -2010 1931 -1998
rect 2047 -1601 2165 -1589
rect 2047 -1998 2053 -1601
rect 2159 -1998 2165 -1601
rect 2047 -2010 2165 -1998
rect 2281 -1601 2399 -1589
rect 2281 -1998 2287 -1601
rect 2393 -1998 2399 -1601
rect 2281 -2010 2399 -1998
rect 2515 -1601 2633 -1589
rect 2515 -1998 2521 -1601
rect 2627 -1998 2633 -1601
rect 2515 -2010 2633 -1998
rect 2749 -1601 2867 -1589
rect 2749 -1998 2755 -1601
rect 2861 -1998 2867 -1601
rect 2749 -2010 2867 -1998
<< properties >>
string FIXED_BBOX -2990 -2129 2990 2129
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 16.0 m 1 nx 25 wmin 0.690 lmin 0.50 class resistor rho 319.8 val 7.98k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
