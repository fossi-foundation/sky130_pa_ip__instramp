magic
tech sky130A
timestamp 1730739923
<< pwell >>
rect -790 -597 790 597
<< mvnnmos >>
rect -676 368 -476 468
rect -388 368 -188 468
rect -100 368 100 468
rect 188 368 388 468
rect 476 368 676 468
rect -676 159 -476 259
rect -388 159 -188 259
rect -100 159 100 259
rect 188 159 388 259
rect 476 159 676 259
rect -676 -50 -476 50
rect -388 -50 -188 50
rect -100 -50 100 50
rect 188 -50 388 50
rect 476 -50 676 50
rect -676 -259 -476 -159
rect -388 -259 -188 -159
rect -100 -259 100 -159
rect 188 -259 388 -159
rect 476 -259 676 -159
rect -676 -468 -476 -368
rect -388 -468 -188 -368
rect -100 -468 100 -368
rect 188 -468 388 -368
rect 476 -468 676 -368
<< mvndiff >>
rect -705 462 -676 468
rect -705 374 -699 462
rect -682 374 -676 462
rect -705 368 -676 374
rect -476 462 -447 468
rect -476 374 -470 462
rect -453 374 -447 462
rect -476 368 -447 374
rect -417 462 -388 468
rect -417 374 -411 462
rect -394 374 -388 462
rect -417 368 -388 374
rect -188 462 -159 468
rect -188 374 -182 462
rect -165 374 -159 462
rect -188 368 -159 374
rect -129 462 -100 468
rect -129 374 -123 462
rect -106 374 -100 462
rect -129 368 -100 374
rect 100 462 129 468
rect 100 374 106 462
rect 123 374 129 462
rect 100 368 129 374
rect 159 462 188 468
rect 159 374 165 462
rect 182 374 188 462
rect 159 368 188 374
rect 388 462 417 468
rect 388 374 394 462
rect 411 374 417 462
rect 388 368 417 374
rect 447 462 476 468
rect 447 374 453 462
rect 470 374 476 462
rect 447 368 476 374
rect 676 462 705 468
rect 676 374 682 462
rect 699 374 705 462
rect 676 368 705 374
rect -705 253 -676 259
rect -705 165 -699 253
rect -682 165 -676 253
rect -705 159 -676 165
rect -476 253 -447 259
rect -476 165 -470 253
rect -453 165 -447 253
rect -476 159 -447 165
rect -417 253 -388 259
rect -417 165 -411 253
rect -394 165 -388 253
rect -417 159 -388 165
rect -188 253 -159 259
rect -188 165 -182 253
rect -165 165 -159 253
rect -188 159 -159 165
rect -129 253 -100 259
rect -129 165 -123 253
rect -106 165 -100 253
rect -129 159 -100 165
rect 100 253 129 259
rect 100 165 106 253
rect 123 165 129 253
rect 100 159 129 165
rect 159 253 188 259
rect 159 165 165 253
rect 182 165 188 253
rect 159 159 188 165
rect 388 253 417 259
rect 388 165 394 253
rect 411 165 417 253
rect 388 159 417 165
rect 447 253 476 259
rect 447 165 453 253
rect 470 165 476 253
rect 447 159 476 165
rect 676 253 705 259
rect 676 165 682 253
rect 699 165 705 253
rect 676 159 705 165
rect -705 44 -676 50
rect -705 -44 -699 44
rect -682 -44 -676 44
rect -705 -50 -676 -44
rect -476 44 -447 50
rect -476 -44 -470 44
rect -453 -44 -447 44
rect -476 -50 -447 -44
rect -417 44 -388 50
rect -417 -44 -411 44
rect -394 -44 -388 44
rect -417 -50 -388 -44
rect -188 44 -159 50
rect -188 -44 -182 44
rect -165 -44 -159 44
rect -188 -50 -159 -44
rect -129 44 -100 50
rect -129 -44 -123 44
rect -106 -44 -100 44
rect -129 -50 -100 -44
rect 100 44 129 50
rect 100 -44 106 44
rect 123 -44 129 44
rect 100 -50 129 -44
rect 159 44 188 50
rect 159 -44 165 44
rect 182 -44 188 44
rect 159 -50 188 -44
rect 388 44 417 50
rect 388 -44 394 44
rect 411 -44 417 44
rect 388 -50 417 -44
rect 447 44 476 50
rect 447 -44 453 44
rect 470 -44 476 44
rect 447 -50 476 -44
rect 676 44 705 50
rect 676 -44 682 44
rect 699 -44 705 44
rect 676 -50 705 -44
rect -705 -165 -676 -159
rect -705 -253 -699 -165
rect -682 -253 -676 -165
rect -705 -259 -676 -253
rect -476 -165 -447 -159
rect -476 -253 -470 -165
rect -453 -253 -447 -165
rect -476 -259 -447 -253
rect -417 -165 -388 -159
rect -417 -253 -411 -165
rect -394 -253 -388 -165
rect -417 -259 -388 -253
rect -188 -165 -159 -159
rect -188 -253 -182 -165
rect -165 -253 -159 -165
rect -188 -259 -159 -253
rect -129 -165 -100 -159
rect -129 -253 -123 -165
rect -106 -253 -100 -165
rect -129 -259 -100 -253
rect 100 -165 129 -159
rect 100 -253 106 -165
rect 123 -253 129 -165
rect 100 -259 129 -253
rect 159 -165 188 -159
rect 159 -253 165 -165
rect 182 -253 188 -165
rect 159 -259 188 -253
rect 388 -165 417 -159
rect 388 -253 394 -165
rect 411 -253 417 -165
rect 388 -259 417 -253
rect 447 -165 476 -159
rect 447 -253 453 -165
rect 470 -253 476 -165
rect 447 -259 476 -253
rect 676 -165 705 -159
rect 676 -253 682 -165
rect 699 -253 705 -165
rect 676 -259 705 -253
rect -705 -374 -676 -368
rect -705 -462 -699 -374
rect -682 -462 -676 -374
rect -705 -468 -676 -462
rect -476 -374 -447 -368
rect -476 -462 -470 -374
rect -453 -462 -447 -374
rect -476 -468 -447 -462
rect -417 -374 -388 -368
rect -417 -462 -411 -374
rect -394 -462 -388 -374
rect -417 -468 -388 -462
rect -188 -374 -159 -368
rect -188 -462 -182 -374
rect -165 -462 -159 -374
rect -188 -468 -159 -462
rect -129 -374 -100 -368
rect -129 -462 -123 -374
rect -106 -462 -100 -374
rect -129 -468 -100 -462
rect 100 -374 129 -368
rect 100 -462 106 -374
rect 123 -462 129 -374
rect 100 -468 129 -462
rect 159 -374 188 -368
rect 159 -462 165 -374
rect 182 -462 188 -374
rect 159 -468 188 -462
rect 388 -374 417 -368
rect 388 -462 394 -374
rect 411 -462 417 -374
rect 388 -468 417 -462
rect 447 -374 476 -368
rect 447 -462 453 -374
rect 470 -462 476 -374
rect 447 -468 476 -462
rect 676 -374 705 -368
rect 676 -462 682 -374
rect 699 -462 705 -374
rect 676 -468 705 -462
<< mvndiffc >>
rect -699 374 -682 462
rect -470 374 -453 462
rect -411 374 -394 462
rect -182 374 -165 462
rect -123 374 -106 462
rect 106 374 123 462
rect 165 374 182 462
rect 394 374 411 462
rect 453 374 470 462
rect 682 374 699 462
rect -699 165 -682 253
rect -470 165 -453 253
rect -411 165 -394 253
rect -182 165 -165 253
rect -123 165 -106 253
rect 106 165 123 253
rect 165 165 182 253
rect 394 165 411 253
rect 453 165 470 253
rect 682 165 699 253
rect -699 -44 -682 44
rect -470 -44 -453 44
rect -411 -44 -394 44
rect -182 -44 -165 44
rect -123 -44 -106 44
rect 106 -44 123 44
rect 165 -44 182 44
rect 394 -44 411 44
rect 453 -44 470 44
rect 682 -44 699 44
rect -699 -253 -682 -165
rect -470 -253 -453 -165
rect -411 -253 -394 -165
rect -182 -253 -165 -165
rect -123 -253 -106 -165
rect 106 -253 123 -165
rect 165 -253 182 -165
rect 394 -253 411 -165
rect 453 -253 470 -165
rect 682 -253 699 -165
rect -699 -462 -682 -374
rect -470 -462 -453 -374
rect -411 -462 -394 -374
rect -182 -462 -165 -374
rect -123 -462 -106 -374
rect 106 -462 123 -374
rect 165 -462 182 -374
rect 394 -462 411 -374
rect 453 -462 470 -374
rect 682 -462 699 -374
<< mvpsubdiff >>
rect -772 573 772 579
rect -772 556 -718 573
rect 718 556 772 573
rect -772 550 772 556
rect -772 525 -743 550
rect -772 -525 -766 525
rect -749 -525 -743 525
rect 743 525 772 550
rect -772 -550 -743 -525
rect 743 -525 749 525
rect 766 -525 772 525
rect 743 -550 772 -525
rect -772 -556 772 -550
rect -772 -573 -718 -556
rect 718 -573 772 -556
rect -772 -579 772 -573
<< mvpsubdiffcont >>
rect -718 556 718 573
rect -766 -525 -749 525
rect 749 -525 766 525
rect -718 -573 718 -556
<< poly >>
rect -676 504 -476 512
rect -676 487 -668 504
rect -484 487 -476 504
rect -676 468 -476 487
rect -388 504 -188 512
rect -388 487 -380 504
rect -196 487 -188 504
rect -388 468 -188 487
rect -100 504 100 512
rect -100 487 -92 504
rect 92 487 100 504
rect -100 468 100 487
rect 188 504 388 512
rect 188 487 196 504
rect 380 487 388 504
rect 188 468 388 487
rect 476 504 676 512
rect 476 487 484 504
rect 668 487 676 504
rect 476 468 676 487
rect -676 349 -476 368
rect -676 332 -668 349
rect -484 332 -476 349
rect -676 324 -476 332
rect -388 349 -188 368
rect -388 332 -380 349
rect -196 332 -188 349
rect -388 324 -188 332
rect -100 349 100 368
rect -100 332 -92 349
rect 92 332 100 349
rect -100 324 100 332
rect 188 349 388 368
rect 188 332 196 349
rect 380 332 388 349
rect 188 324 388 332
rect 476 349 676 368
rect 476 332 484 349
rect 668 332 676 349
rect 476 324 676 332
rect -676 295 -476 303
rect -676 278 -668 295
rect -484 278 -476 295
rect -676 259 -476 278
rect -388 295 -188 303
rect -388 278 -380 295
rect -196 278 -188 295
rect -388 259 -188 278
rect -100 295 100 303
rect -100 278 -92 295
rect 92 278 100 295
rect -100 259 100 278
rect 188 295 388 303
rect 188 278 196 295
rect 380 278 388 295
rect 188 259 388 278
rect 476 295 676 303
rect 476 278 484 295
rect 668 278 676 295
rect 476 259 676 278
rect -676 140 -476 159
rect -676 123 -668 140
rect -484 123 -476 140
rect -676 115 -476 123
rect -388 140 -188 159
rect -388 123 -380 140
rect -196 123 -188 140
rect -388 115 -188 123
rect -100 140 100 159
rect -100 123 -92 140
rect 92 123 100 140
rect -100 115 100 123
rect 188 140 388 159
rect 188 123 196 140
rect 380 123 388 140
rect 188 115 388 123
rect 476 140 676 159
rect 476 123 484 140
rect 668 123 676 140
rect 476 115 676 123
rect -676 86 -476 94
rect -676 69 -668 86
rect -484 69 -476 86
rect -676 50 -476 69
rect -388 86 -188 94
rect -388 69 -380 86
rect -196 69 -188 86
rect -388 50 -188 69
rect -100 86 100 94
rect -100 69 -92 86
rect 92 69 100 86
rect -100 50 100 69
rect 188 86 388 94
rect 188 69 196 86
rect 380 69 388 86
rect 188 50 388 69
rect 476 86 676 94
rect 476 69 484 86
rect 668 69 676 86
rect 476 50 676 69
rect -676 -69 -476 -50
rect -676 -86 -668 -69
rect -484 -86 -476 -69
rect -676 -94 -476 -86
rect -388 -69 -188 -50
rect -388 -86 -380 -69
rect -196 -86 -188 -69
rect -388 -94 -188 -86
rect -100 -69 100 -50
rect -100 -86 -92 -69
rect 92 -86 100 -69
rect -100 -94 100 -86
rect 188 -69 388 -50
rect 188 -86 196 -69
rect 380 -86 388 -69
rect 188 -94 388 -86
rect 476 -69 676 -50
rect 476 -86 484 -69
rect 668 -86 676 -69
rect 476 -94 676 -86
rect -676 -123 -476 -115
rect -676 -140 -668 -123
rect -484 -140 -476 -123
rect -676 -159 -476 -140
rect -388 -123 -188 -115
rect -388 -140 -380 -123
rect -196 -140 -188 -123
rect -388 -159 -188 -140
rect -100 -123 100 -115
rect -100 -140 -92 -123
rect 92 -140 100 -123
rect -100 -159 100 -140
rect 188 -123 388 -115
rect 188 -140 196 -123
rect 380 -140 388 -123
rect 188 -159 388 -140
rect 476 -123 676 -115
rect 476 -140 484 -123
rect 668 -140 676 -123
rect 476 -159 676 -140
rect -676 -278 -476 -259
rect -676 -295 -668 -278
rect -484 -295 -476 -278
rect -676 -303 -476 -295
rect -388 -278 -188 -259
rect -388 -295 -380 -278
rect -196 -295 -188 -278
rect -388 -303 -188 -295
rect -100 -278 100 -259
rect -100 -295 -92 -278
rect 92 -295 100 -278
rect -100 -303 100 -295
rect 188 -278 388 -259
rect 188 -295 196 -278
rect 380 -295 388 -278
rect 188 -303 388 -295
rect 476 -278 676 -259
rect 476 -295 484 -278
rect 668 -295 676 -278
rect 476 -303 676 -295
rect -676 -332 -476 -324
rect -676 -349 -668 -332
rect -484 -349 -476 -332
rect -676 -368 -476 -349
rect -388 -332 -188 -324
rect -388 -349 -380 -332
rect -196 -349 -188 -332
rect -388 -368 -188 -349
rect -100 -332 100 -324
rect -100 -349 -92 -332
rect 92 -349 100 -332
rect -100 -368 100 -349
rect 188 -332 388 -324
rect 188 -349 196 -332
rect 380 -349 388 -332
rect 188 -368 388 -349
rect 476 -332 676 -324
rect 476 -349 484 -332
rect 668 -349 676 -332
rect 476 -368 676 -349
rect -676 -487 -476 -468
rect -676 -504 -668 -487
rect -484 -504 -476 -487
rect -676 -512 -476 -504
rect -388 -487 -188 -468
rect -388 -504 -380 -487
rect -196 -504 -188 -487
rect -388 -512 -188 -504
rect -100 -487 100 -468
rect -100 -504 -92 -487
rect 92 -504 100 -487
rect -100 -512 100 -504
rect 188 -487 388 -468
rect 188 -504 196 -487
rect 380 -504 388 -487
rect 188 -512 388 -504
rect 476 -487 676 -468
rect 476 -504 484 -487
rect 668 -504 676 -487
rect 476 -512 676 -504
<< polycont >>
rect -668 487 -484 504
rect -380 487 -196 504
rect -92 487 92 504
rect 196 487 380 504
rect 484 487 668 504
rect -668 332 -484 349
rect -380 332 -196 349
rect -92 332 92 349
rect 196 332 380 349
rect 484 332 668 349
rect -668 278 -484 295
rect -380 278 -196 295
rect -92 278 92 295
rect 196 278 380 295
rect 484 278 668 295
rect -668 123 -484 140
rect -380 123 -196 140
rect -92 123 92 140
rect 196 123 380 140
rect 484 123 668 140
rect -668 69 -484 86
rect -380 69 -196 86
rect -92 69 92 86
rect 196 69 380 86
rect 484 69 668 86
rect -668 -86 -484 -69
rect -380 -86 -196 -69
rect -92 -86 92 -69
rect 196 -86 380 -69
rect 484 -86 668 -69
rect -668 -140 -484 -123
rect -380 -140 -196 -123
rect -92 -140 92 -123
rect 196 -140 380 -123
rect 484 -140 668 -123
rect -668 -295 -484 -278
rect -380 -295 -196 -278
rect -92 -295 92 -278
rect 196 -295 380 -278
rect 484 -295 668 -278
rect -668 -349 -484 -332
rect -380 -349 -196 -332
rect -92 -349 92 -332
rect 196 -349 380 -332
rect 484 -349 668 -332
rect -668 -504 -484 -487
rect -380 -504 -196 -487
rect -92 -504 92 -487
rect 196 -504 380 -487
rect 484 -504 668 -487
<< locali >>
rect -766 556 -718 573
rect 718 556 766 573
rect -766 525 -749 556
rect 749 525 766 556
rect -676 487 -668 504
rect -484 487 -476 504
rect -388 487 -380 504
rect -196 487 -188 504
rect -100 487 -92 504
rect 92 487 100 504
rect 188 487 196 504
rect 380 487 388 504
rect 476 487 484 504
rect 668 487 676 504
rect -699 462 -682 470
rect -699 366 -682 374
rect -470 462 -453 470
rect -470 366 -453 374
rect -411 462 -394 470
rect -411 366 -394 374
rect -182 462 -165 470
rect -182 366 -165 374
rect -123 462 -106 470
rect -123 366 -106 374
rect 106 462 123 470
rect 106 366 123 374
rect 165 462 182 470
rect 165 366 182 374
rect 394 462 411 470
rect 394 366 411 374
rect 453 462 470 470
rect 453 366 470 374
rect 682 462 699 470
rect 682 366 699 374
rect -676 332 -668 349
rect -484 332 -476 349
rect -388 332 -380 349
rect -196 332 -188 349
rect -100 332 -92 349
rect 92 332 100 349
rect 188 332 196 349
rect 380 332 388 349
rect 476 332 484 349
rect 668 332 676 349
rect -676 278 -668 295
rect -484 278 -476 295
rect -388 278 -380 295
rect -196 278 -188 295
rect -100 278 -92 295
rect 92 278 100 295
rect 188 278 196 295
rect 380 278 388 295
rect 476 278 484 295
rect 668 278 676 295
rect -699 253 -682 261
rect -699 157 -682 165
rect -470 253 -453 261
rect -470 157 -453 165
rect -411 253 -394 261
rect -411 157 -394 165
rect -182 253 -165 261
rect -182 157 -165 165
rect -123 253 -106 261
rect -123 157 -106 165
rect 106 253 123 261
rect 106 157 123 165
rect 165 253 182 261
rect 165 157 182 165
rect 394 253 411 261
rect 394 157 411 165
rect 453 253 470 261
rect 453 157 470 165
rect 682 253 699 261
rect 682 157 699 165
rect -676 123 -668 140
rect -484 123 -476 140
rect -388 123 -380 140
rect -196 123 -188 140
rect -100 123 -92 140
rect 92 123 100 140
rect 188 123 196 140
rect 380 123 388 140
rect 476 123 484 140
rect 668 123 676 140
rect -676 69 -668 86
rect -484 69 -476 86
rect -388 69 -380 86
rect -196 69 -188 86
rect -100 69 -92 86
rect 92 69 100 86
rect 188 69 196 86
rect 380 69 388 86
rect 476 69 484 86
rect 668 69 676 86
rect -699 44 -682 52
rect -699 -52 -682 -44
rect -470 44 -453 52
rect -470 -52 -453 -44
rect -411 44 -394 52
rect -411 -52 -394 -44
rect -182 44 -165 52
rect -182 -52 -165 -44
rect -123 44 -106 52
rect -123 -52 -106 -44
rect 106 44 123 52
rect 106 -52 123 -44
rect 165 44 182 52
rect 165 -52 182 -44
rect 394 44 411 52
rect 394 -52 411 -44
rect 453 44 470 52
rect 453 -52 470 -44
rect 682 44 699 52
rect 682 -52 699 -44
rect -676 -86 -668 -69
rect -484 -86 -476 -69
rect -388 -86 -380 -69
rect -196 -86 -188 -69
rect -100 -86 -92 -69
rect 92 -86 100 -69
rect 188 -86 196 -69
rect 380 -86 388 -69
rect 476 -86 484 -69
rect 668 -86 676 -69
rect -676 -140 -668 -123
rect -484 -140 -476 -123
rect -388 -140 -380 -123
rect -196 -140 -188 -123
rect -100 -140 -92 -123
rect 92 -140 100 -123
rect 188 -140 196 -123
rect 380 -140 388 -123
rect 476 -140 484 -123
rect 668 -140 676 -123
rect -699 -165 -682 -157
rect -699 -261 -682 -253
rect -470 -165 -453 -157
rect -470 -261 -453 -253
rect -411 -165 -394 -157
rect -411 -261 -394 -253
rect -182 -165 -165 -157
rect -182 -261 -165 -253
rect -123 -165 -106 -157
rect -123 -261 -106 -253
rect 106 -165 123 -157
rect 106 -261 123 -253
rect 165 -165 182 -157
rect 165 -261 182 -253
rect 394 -165 411 -157
rect 394 -261 411 -253
rect 453 -165 470 -157
rect 453 -261 470 -253
rect 682 -165 699 -157
rect 682 -261 699 -253
rect -676 -295 -668 -278
rect -484 -295 -476 -278
rect -388 -295 -380 -278
rect -196 -295 -188 -278
rect -100 -295 -92 -278
rect 92 -295 100 -278
rect 188 -295 196 -278
rect 380 -295 388 -278
rect 476 -295 484 -278
rect 668 -295 676 -278
rect -676 -349 -668 -332
rect -484 -349 -476 -332
rect -388 -349 -380 -332
rect -196 -349 -188 -332
rect -100 -349 -92 -332
rect 92 -349 100 -332
rect 188 -349 196 -332
rect 380 -349 388 -332
rect 476 -349 484 -332
rect 668 -349 676 -332
rect -699 -374 -682 -366
rect -699 -470 -682 -462
rect -470 -374 -453 -366
rect -470 -470 -453 -462
rect -411 -374 -394 -366
rect -411 -470 -394 -462
rect -182 -374 -165 -366
rect -182 -470 -165 -462
rect -123 -374 -106 -366
rect -123 -470 -106 -462
rect 106 -374 123 -366
rect 106 -470 123 -462
rect 165 -374 182 -366
rect 165 -470 182 -462
rect 394 -374 411 -366
rect 394 -470 411 -462
rect 453 -374 470 -366
rect 453 -470 470 -462
rect 682 -374 699 -366
rect 682 -470 699 -462
rect -676 -504 -668 -487
rect -484 -504 -476 -487
rect -388 -504 -380 -487
rect -196 -504 -188 -487
rect -100 -504 -92 -487
rect 92 -504 100 -487
rect 188 -504 196 -487
rect 380 -504 388 -487
rect 476 -504 484 -487
rect 668 -504 676 -487
rect -766 -556 -749 -525
rect 749 -556 766 -525
rect -766 -573 -718 -556
rect 718 -573 766 -556
<< viali >>
rect -668 487 -484 504
rect -380 487 -196 504
rect -92 487 92 504
rect 196 487 380 504
rect 484 487 668 504
rect -699 374 -682 462
rect -470 374 -453 462
rect -411 374 -394 462
rect -182 374 -165 462
rect -123 374 -106 462
rect 106 374 123 462
rect 165 374 182 462
rect 394 374 411 462
rect 453 374 470 462
rect 682 374 699 462
rect -668 332 -484 349
rect -380 332 -196 349
rect -92 332 92 349
rect 196 332 380 349
rect 484 332 668 349
rect -668 278 -484 295
rect -380 278 -196 295
rect -92 278 92 295
rect 196 278 380 295
rect 484 278 668 295
rect -699 165 -682 253
rect -470 165 -453 253
rect -411 165 -394 253
rect -182 165 -165 253
rect -123 165 -106 253
rect 106 165 123 253
rect 165 165 182 253
rect 394 165 411 253
rect 453 165 470 253
rect 682 165 699 253
rect -668 123 -484 140
rect -380 123 -196 140
rect -92 123 92 140
rect 196 123 380 140
rect 484 123 668 140
rect -668 69 -484 86
rect -380 69 -196 86
rect -92 69 92 86
rect 196 69 380 86
rect 484 69 668 86
rect -699 -44 -682 44
rect -470 -44 -453 44
rect -411 -44 -394 44
rect -182 -44 -165 44
rect -123 -44 -106 44
rect 106 -44 123 44
rect 165 -44 182 44
rect 394 -44 411 44
rect 453 -44 470 44
rect 682 -44 699 44
rect -668 -86 -484 -69
rect -380 -86 -196 -69
rect -92 -86 92 -69
rect 196 -86 380 -69
rect 484 -86 668 -69
rect -668 -140 -484 -123
rect -380 -140 -196 -123
rect -92 -140 92 -123
rect 196 -140 380 -123
rect 484 -140 668 -123
rect -699 -253 -682 -165
rect -470 -253 -453 -165
rect -411 -253 -394 -165
rect -182 -253 -165 -165
rect -123 -253 -106 -165
rect 106 -253 123 -165
rect 165 -253 182 -165
rect 394 -253 411 -165
rect 453 -253 470 -165
rect 682 -253 699 -165
rect -668 -295 -484 -278
rect -380 -295 -196 -278
rect -92 -295 92 -278
rect 196 -295 380 -278
rect 484 -295 668 -278
rect -668 -349 -484 -332
rect -380 -349 -196 -332
rect -92 -349 92 -332
rect 196 -349 380 -332
rect 484 -349 668 -332
rect -699 -462 -682 -374
rect -470 -462 -453 -374
rect -411 -462 -394 -374
rect -182 -462 -165 -374
rect -123 -462 -106 -374
rect 106 -462 123 -374
rect 165 -462 182 -374
rect 394 -462 411 -374
rect 453 -462 470 -374
rect 682 -462 699 -374
rect -668 -504 -484 -487
rect -380 -504 -196 -487
rect -92 -504 92 -487
rect 196 -504 380 -487
rect 484 -504 668 -487
<< metal1 >>
rect -674 504 -478 507
rect -674 487 -668 504
rect -484 487 -478 504
rect -674 484 -478 487
rect -386 504 -190 507
rect -386 487 -380 504
rect -196 487 -190 504
rect -386 484 -190 487
rect -98 504 98 507
rect -98 487 -92 504
rect 92 487 98 504
rect -98 484 98 487
rect 190 504 386 507
rect 190 487 196 504
rect 380 487 386 504
rect 190 484 386 487
rect 478 504 674 507
rect 478 487 484 504
rect 668 487 674 504
rect 478 484 674 487
rect -702 462 -679 468
rect -702 374 -699 462
rect -682 374 -679 462
rect -702 368 -679 374
rect -473 462 -450 468
rect -473 374 -470 462
rect -453 374 -450 462
rect -473 368 -450 374
rect -414 462 -391 468
rect -414 374 -411 462
rect -394 374 -391 462
rect -414 368 -391 374
rect -185 462 -162 468
rect -185 374 -182 462
rect -165 374 -162 462
rect -185 368 -162 374
rect -126 462 -103 468
rect -126 374 -123 462
rect -106 374 -103 462
rect -126 368 -103 374
rect 103 462 126 468
rect 103 374 106 462
rect 123 374 126 462
rect 103 368 126 374
rect 162 462 185 468
rect 162 374 165 462
rect 182 374 185 462
rect 162 368 185 374
rect 391 462 414 468
rect 391 374 394 462
rect 411 374 414 462
rect 391 368 414 374
rect 450 462 473 468
rect 450 374 453 462
rect 470 374 473 462
rect 450 368 473 374
rect 679 462 702 468
rect 679 374 682 462
rect 699 374 702 462
rect 679 368 702 374
rect -674 349 -478 352
rect -674 332 -668 349
rect -484 332 -478 349
rect -674 329 -478 332
rect -386 349 -190 352
rect -386 332 -380 349
rect -196 332 -190 349
rect -386 329 -190 332
rect -98 349 98 352
rect -98 332 -92 349
rect 92 332 98 349
rect -98 329 98 332
rect 190 349 386 352
rect 190 332 196 349
rect 380 332 386 349
rect 190 329 386 332
rect 478 349 674 352
rect 478 332 484 349
rect 668 332 674 349
rect 478 329 674 332
rect -674 295 -478 298
rect -674 278 -668 295
rect -484 278 -478 295
rect -674 275 -478 278
rect -386 295 -190 298
rect -386 278 -380 295
rect -196 278 -190 295
rect -386 275 -190 278
rect -98 295 98 298
rect -98 278 -92 295
rect 92 278 98 295
rect -98 275 98 278
rect 190 295 386 298
rect 190 278 196 295
rect 380 278 386 295
rect 190 275 386 278
rect 478 295 674 298
rect 478 278 484 295
rect 668 278 674 295
rect 478 275 674 278
rect -702 253 -679 259
rect -702 165 -699 253
rect -682 165 -679 253
rect -702 159 -679 165
rect -473 253 -450 259
rect -473 165 -470 253
rect -453 165 -450 253
rect -473 159 -450 165
rect -414 253 -391 259
rect -414 165 -411 253
rect -394 165 -391 253
rect -414 159 -391 165
rect -185 253 -162 259
rect -185 165 -182 253
rect -165 165 -162 253
rect -185 159 -162 165
rect -126 253 -103 259
rect -126 165 -123 253
rect -106 165 -103 253
rect -126 159 -103 165
rect 103 253 126 259
rect 103 165 106 253
rect 123 165 126 253
rect 103 159 126 165
rect 162 253 185 259
rect 162 165 165 253
rect 182 165 185 253
rect 162 159 185 165
rect 391 253 414 259
rect 391 165 394 253
rect 411 165 414 253
rect 391 159 414 165
rect 450 253 473 259
rect 450 165 453 253
rect 470 165 473 253
rect 450 159 473 165
rect 679 253 702 259
rect 679 165 682 253
rect 699 165 702 253
rect 679 159 702 165
rect -674 140 -478 143
rect -674 123 -668 140
rect -484 123 -478 140
rect -674 120 -478 123
rect -386 140 -190 143
rect -386 123 -380 140
rect -196 123 -190 140
rect -386 120 -190 123
rect -98 140 98 143
rect -98 123 -92 140
rect 92 123 98 140
rect -98 120 98 123
rect 190 140 386 143
rect 190 123 196 140
rect 380 123 386 140
rect 190 120 386 123
rect 478 140 674 143
rect 478 123 484 140
rect 668 123 674 140
rect 478 120 674 123
rect -674 86 -478 89
rect -674 69 -668 86
rect -484 69 -478 86
rect -674 66 -478 69
rect -386 86 -190 89
rect -386 69 -380 86
rect -196 69 -190 86
rect -386 66 -190 69
rect -98 86 98 89
rect -98 69 -92 86
rect 92 69 98 86
rect -98 66 98 69
rect 190 86 386 89
rect 190 69 196 86
rect 380 69 386 86
rect 190 66 386 69
rect 478 86 674 89
rect 478 69 484 86
rect 668 69 674 86
rect 478 66 674 69
rect -702 44 -679 50
rect -702 -44 -699 44
rect -682 -44 -679 44
rect -702 -50 -679 -44
rect -473 44 -450 50
rect -473 -44 -470 44
rect -453 -44 -450 44
rect -473 -50 -450 -44
rect -414 44 -391 50
rect -414 -44 -411 44
rect -394 -44 -391 44
rect -414 -50 -391 -44
rect -185 44 -162 50
rect -185 -44 -182 44
rect -165 -44 -162 44
rect -185 -50 -162 -44
rect -126 44 -103 50
rect -126 -44 -123 44
rect -106 -44 -103 44
rect -126 -50 -103 -44
rect 103 44 126 50
rect 103 -44 106 44
rect 123 -44 126 44
rect 103 -50 126 -44
rect 162 44 185 50
rect 162 -44 165 44
rect 182 -44 185 44
rect 162 -50 185 -44
rect 391 44 414 50
rect 391 -44 394 44
rect 411 -44 414 44
rect 391 -50 414 -44
rect 450 44 473 50
rect 450 -44 453 44
rect 470 -44 473 44
rect 450 -50 473 -44
rect 679 44 702 50
rect 679 -44 682 44
rect 699 -44 702 44
rect 679 -50 702 -44
rect -674 -69 -478 -66
rect -674 -86 -668 -69
rect -484 -86 -478 -69
rect -674 -89 -478 -86
rect -386 -69 -190 -66
rect -386 -86 -380 -69
rect -196 -86 -190 -69
rect -386 -89 -190 -86
rect -98 -69 98 -66
rect -98 -86 -92 -69
rect 92 -86 98 -69
rect -98 -89 98 -86
rect 190 -69 386 -66
rect 190 -86 196 -69
rect 380 -86 386 -69
rect 190 -89 386 -86
rect 478 -69 674 -66
rect 478 -86 484 -69
rect 668 -86 674 -69
rect 478 -89 674 -86
rect -674 -123 -478 -120
rect -674 -140 -668 -123
rect -484 -140 -478 -123
rect -674 -143 -478 -140
rect -386 -123 -190 -120
rect -386 -140 -380 -123
rect -196 -140 -190 -123
rect -386 -143 -190 -140
rect -98 -123 98 -120
rect -98 -140 -92 -123
rect 92 -140 98 -123
rect -98 -143 98 -140
rect 190 -123 386 -120
rect 190 -140 196 -123
rect 380 -140 386 -123
rect 190 -143 386 -140
rect 478 -123 674 -120
rect 478 -140 484 -123
rect 668 -140 674 -123
rect 478 -143 674 -140
rect -702 -165 -679 -159
rect -702 -253 -699 -165
rect -682 -253 -679 -165
rect -702 -259 -679 -253
rect -473 -165 -450 -159
rect -473 -253 -470 -165
rect -453 -253 -450 -165
rect -473 -259 -450 -253
rect -414 -165 -391 -159
rect -414 -253 -411 -165
rect -394 -253 -391 -165
rect -414 -259 -391 -253
rect -185 -165 -162 -159
rect -185 -253 -182 -165
rect -165 -253 -162 -165
rect -185 -259 -162 -253
rect -126 -165 -103 -159
rect -126 -253 -123 -165
rect -106 -253 -103 -165
rect -126 -259 -103 -253
rect 103 -165 126 -159
rect 103 -253 106 -165
rect 123 -253 126 -165
rect 103 -259 126 -253
rect 162 -165 185 -159
rect 162 -253 165 -165
rect 182 -253 185 -165
rect 162 -259 185 -253
rect 391 -165 414 -159
rect 391 -253 394 -165
rect 411 -253 414 -165
rect 391 -259 414 -253
rect 450 -165 473 -159
rect 450 -253 453 -165
rect 470 -253 473 -165
rect 450 -259 473 -253
rect 679 -165 702 -159
rect 679 -253 682 -165
rect 699 -253 702 -165
rect 679 -259 702 -253
rect -674 -278 -478 -275
rect -674 -295 -668 -278
rect -484 -295 -478 -278
rect -674 -298 -478 -295
rect -386 -278 -190 -275
rect -386 -295 -380 -278
rect -196 -295 -190 -278
rect -386 -298 -190 -295
rect -98 -278 98 -275
rect -98 -295 -92 -278
rect 92 -295 98 -278
rect -98 -298 98 -295
rect 190 -278 386 -275
rect 190 -295 196 -278
rect 380 -295 386 -278
rect 190 -298 386 -295
rect 478 -278 674 -275
rect 478 -295 484 -278
rect 668 -295 674 -278
rect 478 -298 674 -295
rect -674 -332 -478 -329
rect -674 -349 -668 -332
rect -484 -349 -478 -332
rect -674 -352 -478 -349
rect -386 -332 -190 -329
rect -386 -349 -380 -332
rect -196 -349 -190 -332
rect -386 -352 -190 -349
rect -98 -332 98 -329
rect -98 -349 -92 -332
rect 92 -349 98 -332
rect -98 -352 98 -349
rect 190 -332 386 -329
rect 190 -349 196 -332
rect 380 -349 386 -332
rect 190 -352 386 -349
rect 478 -332 674 -329
rect 478 -349 484 -332
rect 668 -349 674 -332
rect 478 -352 674 -349
rect -702 -374 -679 -368
rect -702 -462 -699 -374
rect -682 -462 -679 -374
rect -702 -468 -679 -462
rect -473 -374 -450 -368
rect -473 -462 -470 -374
rect -453 -462 -450 -374
rect -473 -468 -450 -462
rect -414 -374 -391 -368
rect -414 -462 -411 -374
rect -394 -462 -391 -374
rect -414 -468 -391 -462
rect -185 -374 -162 -368
rect -185 -462 -182 -374
rect -165 -462 -162 -374
rect -185 -468 -162 -462
rect -126 -374 -103 -368
rect -126 -462 -123 -374
rect -106 -462 -103 -374
rect -126 -468 -103 -462
rect 103 -374 126 -368
rect 103 -462 106 -374
rect 123 -462 126 -374
rect 103 -468 126 -462
rect 162 -374 185 -368
rect 162 -462 165 -374
rect 182 -462 185 -374
rect 162 -468 185 -462
rect 391 -374 414 -368
rect 391 -462 394 -374
rect 411 -462 414 -374
rect 391 -468 414 -462
rect 450 -374 473 -368
rect 450 -462 453 -374
rect 470 -462 473 -374
rect 450 -468 473 -462
rect 679 -374 702 -368
rect 679 -462 682 -374
rect 699 -462 702 -374
rect 679 -468 702 -462
rect -674 -487 -478 -484
rect -674 -504 -668 -487
rect -484 -504 -478 -487
rect -674 -507 -478 -504
rect -386 -487 -190 -484
rect -386 -504 -380 -487
rect -196 -504 -190 -487
rect -386 -507 -190 -504
rect -98 -487 98 -484
rect -98 -504 -92 -487
rect 92 -504 98 -487
rect -98 -507 98 -504
rect 190 -487 386 -484
rect 190 -504 196 -487
rect 380 -504 386 -487
rect 190 -507 386 -504
rect 478 -487 674 -484
rect 478 -504 484 -487
rect 668 -504 674 -487
rect 478 -507 674 -504
<< properties >>
string FIXED_BBOX -757 -564 757 564
string gencell sky130_fd_pr__nfet_05v0_nvt
string library sky130
string parameters w 1.0 l 2.0 m 5 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.90 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
