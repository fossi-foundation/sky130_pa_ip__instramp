magic
tech sky130A
magscale 1 2
timestamp 1730950751
<< error_s >>
rect 284 25778 24926 26064
rect 284 21668 570 25778
rect 24640 22998 24926 25778
rect 24638 22712 24926 22998
rect 24638 22052 24924 22712
rect 14720 21966 24924 22052
rect 14720 21766 24926 21966
rect 284 12994 488 21668
rect 14720 15142 15006 21766
rect 284 11948 570 12994
rect 14746 12500 15006 15142
rect 284 3274 486 11948
rect 14720 11930 15006 12500
rect 14720 11644 15320 11930
rect 15034 6818 15320 11644
rect 14736 6532 15320 6818
rect 14736 5422 15022 6532
rect 284 2200 570 3274
rect 14744 2780 15022 5422
rect 284 -6474 484 2200
rect 14736 -4326 15022 2780
rect 284 -11086 570 -6474
rect 14742 -6970 15022 -4326
rect 14736 -7036 15022 -6970
rect 14736 -7322 29514 -7036
rect 29228 -9354 29514 -7322
rect 29224 -9360 29514 -9354
rect 29218 -9366 29224 -9360
rect 29218 -10498 29224 -10492
rect 29228 -10498 29514 -9360
rect 29224 -10504 29514 -10498
rect 29228 -11086 29514 -10504
rect 284 -11372 29514 -11086
<< dnwell >>
rect 364 22792 24846 25984
rect 364 21886 24844 22792
rect 364 21846 24846 21886
rect 364 11850 14926 21846
rect 364 6612 15240 11850
rect 364 -7116 14942 6612
rect 364 -11292 29434 -7116
<< locali >>
rect 9813 21480 11041 21499
rect 9813 18386 9826 21480
rect 9874 21429 11041 21480
rect 9874 18424 9883 21429
rect 10971 20744 11041 21429
rect 10971 18424 10980 20744
rect 9874 18418 10980 18424
rect 9874 18386 9936 18418
rect 9813 18360 9936 18386
rect 10926 18378 10980 18418
rect 11032 18424 11041 20744
rect 11314 21425 12525 21495
rect 11314 20758 11384 21425
rect 11032 18378 11042 18424
rect 11314 18423 11324 20758
rect 10926 18360 11042 18378
rect 9813 18354 11042 18360
rect 11313 18392 11324 18423
rect 11376 18423 11384 20758
rect 12455 20600 12525 21425
rect 12455 18423 12470 20600
rect 11376 18422 12470 18423
rect 11376 18392 11428 18422
rect 11313 18364 11428 18392
rect 12418 18378 12470 18422
rect 12520 18378 12525 20600
rect 12418 18364 12525 18378
rect 11313 18353 12525 18364
rect 12782 21442 14009 21491
rect 12782 21421 13954 21442
rect 12782 21342 12852 21421
rect 12782 18378 12786 21342
rect 12842 18417 12852 21342
rect 13939 18417 13954 21421
rect 12842 18412 13954 18417
rect 12842 18378 12904 18412
rect 12782 18354 12904 18378
rect 13894 18390 13954 18412
rect 14006 18390 14009 21442
rect 13894 18354 14009 18390
rect 12782 18350 14009 18354
rect 12785 18347 14009 18350
rect 9696 11800 15209 11817
rect 9696 11796 9802 11800
rect 9696 6706 9708 11796
rect 9746 11764 9802 11796
rect 15110 11796 15209 11800
rect 15110 11764 15154 11796
rect 9746 11751 15154 11764
rect 9746 6746 9762 11751
rect 15143 6746 15154 11751
rect 9746 6730 15154 6746
rect 9746 6706 10038 6730
rect 9696 6694 10038 6706
rect 14892 6700 15154 6730
rect 15198 6700 15209 11796
rect 14892 6694 15209 6700
rect 9696 6681 15209 6694
rect 9696 6680 15208 6681
rect 466 -7194 29290 -7178
rect 466 -7242 594 -7194
rect 14694 -7234 14944 -7194
rect 29200 -7234 29290 -7194
rect 14694 -7242 29290 -7234
rect 466 -7254 29290 -7242
rect 466 -7340 542 -7254
rect 29214 -7278 29290 -7254
rect 466 -11166 494 -7340
rect 466 -11218 542 -11166
rect 29214 -11182 29238 -7278
rect 29274 -11182 29290 -7278
rect 29214 -11218 29290 -11182
rect 466 -11228 29290 -11218
rect 466 -11276 594 -11228
rect 29198 -11276 29290 -11228
rect 466 -11294 29290 -11276
<< viali >>
rect 9826 18386 9874 21480
rect 9936 18360 10926 18418
rect 10980 18378 11032 20744
rect 11324 18392 11376 20758
rect 11428 18364 12418 18422
rect 12470 18378 12520 20600
rect 12786 18378 12842 21342
rect 12904 18354 13894 18412
rect 13954 18390 14006 21442
rect 9708 6706 9746 11796
rect 9802 11764 15110 11800
rect 10038 6694 14892 6730
rect 15154 6700 15198 11796
rect 594 -7242 14694 -7194
rect 14944 -7234 29200 -7194
rect 494 -11166 548 -7340
rect 29238 -11182 29274 -7278
rect 594 -11276 29198 -11228
<< metal1 >>
rect 24648 28030 24848 28230
rect 24626 27603 24826 27746
rect 917 27546 24826 27603
rect 368 26054 384 26198
rect 598 26054 746 26198
rect 11168 22280 11372 22300
rect 840 22116 914 22206
rect 636 22102 1072 22116
rect 636 22010 652 22102
rect 1056 22010 1072 22102
rect 1225 22096 1299 22196
rect 3280 22096 3354 22196
rect 1225 22022 3354 22096
rect 3625 22096 3699 22196
rect 5680 22096 5754 22196
rect 3625 22022 5754 22096
rect 6025 22096 6099 22196
rect 8080 22096 8154 22196
rect 6025 22022 8154 22096
rect 8425 22096 8499 22196
rect 10480 22096 10554 22196
rect 8425 22022 10554 22096
rect 636 21996 1072 22010
rect 2816 21760 3016 21960
rect 10825 21940 10899 22196
rect 11168 22124 11190 22280
rect 11350 22124 11372 22280
rect 11168 22104 11372 22124
rect 12140 22288 12276 22300
rect 12140 22116 12152 22288
rect 12260 22116 12276 22288
rect 12140 22104 12276 22116
rect 9694 21916 9892 21940
rect 9694 21664 9716 21916
rect 9872 21664 9892 21916
rect 9694 21640 9892 21664
rect 9814 21504 9892 21640
rect 9812 21480 9892 21504
rect 9812 18430 9826 21480
rect 9338 18386 9826 18430
rect 9874 18434 9892 21480
rect 9974 21863 10899 21940
rect 9974 20898 10050 21863
rect 11182 21792 11258 22104
rect 10476 21716 11258 21792
rect 12155 21848 12233 22104
rect 12768 22100 12968 22218
rect 12768 21930 12786 22100
rect 12952 21930 12968 22100
rect 13225 22096 13299 22196
rect 15280 22096 15354 22196
rect 13225 22022 15354 22096
rect 15625 22096 15699 22196
rect 17680 22096 17754 22196
rect 15625 22022 17754 22096
rect 18025 22096 18099 22196
rect 20080 22096 20154 22196
rect 18025 22022 20154 22096
rect 20425 22096 20499 22223
rect 22480 22096 22554 22204
rect 20425 22022 22554 22096
rect 22798 22114 22998 22196
rect 22798 22104 23100 22114
rect 22798 22012 22808 22104
rect 23086 22012 23100 22104
rect 22798 22004 23100 22012
rect 12768 21914 12968 21930
rect 12155 21769 13348 21848
rect 14452 21788 14472 21912
rect 14672 21788 15066 21912
rect 10146 20906 10382 21338
rect 10476 20902 10552 21716
rect 12768 21710 12972 21720
rect 12768 21604 12782 21710
rect 12962 21691 12972 21710
rect 12962 21621 13177 21691
rect 12962 21620 13176 21621
rect 12962 21604 12972 21620
rect 12768 21594 12972 21604
rect 10642 21552 11024 21562
rect 10642 21466 10654 21552
rect 11010 21466 11024 21552
rect 10642 21456 11024 21466
rect 10642 20906 10718 21456
rect 12290 21444 13010 21514
rect 11002 21392 11332 21408
rect 11002 21338 11018 21392
rect 10810 21278 11018 21338
rect 11314 21338 11332 21392
rect 11314 21278 11530 21338
rect 10810 20904 11530 21278
rect 11626 20906 11862 21338
rect 11958 20906 12196 21338
rect 12124 20812 12196 20906
rect 12290 20904 12360 21444
rect 12764 21342 12864 21382
rect 10970 20744 11050 20786
rect 9982 18508 10220 18940
rect 10314 18508 10552 18940
rect 10646 18508 10884 18940
rect 10970 18434 10980 20744
rect 9874 18418 10980 18434
rect 9874 18386 9936 18418
rect 9338 18360 9936 18386
rect 10926 18378 10980 18418
rect 11032 18430 11050 20744
rect 11306 20758 11386 20792
rect 11306 18430 11324 20758
rect 11032 18392 11324 18430
rect 11376 18432 11386 20758
rect 12124 20704 12684 20812
rect 12450 20600 12534 20634
rect 11458 18506 11696 18938
rect 11790 18506 12028 18938
rect 12122 18506 12360 18938
rect 12450 18432 12470 20600
rect 11376 18422 12470 18432
rect 11376 18392 11428 18422
rect 11032 18378 11428 18392
rect 10926 18364 11428 18378
rect 12418 18378 12470 18422
rect 12520 18432 12534 20600
rect 12520 18378 12536 18432
rect 12418 18364 12536 18378
rect 10926 18360 12536 18364
rect 9338 18340 12536 18360
rect 12628 18284 12684 20704
rect 12764 18378 12786 21342
rect 12842 18432 12864 21342
rect 12940 20906 13010 21444
rect 13106 20906 13176 21620
rect 13270 20906 13348 21769
rect 13770 21610 14728 21728
rect 14908 21610 14933 21728
rect 13438 20902 13676 21340
rect 13770 20906 13844 21610
rect 14278 21530 14620 21546
rect 13932 21442 14034 21498
rect 12940 18506 13178 18938
rect 13272 18506 13510 18938
rect 13604 18506 13842 18938
rect 13932 18432 13954 21442
rect 12842 18412 13954 18432
rect 12842 18378 12904 18412
rect 12764 18354 12904 18378
rect 13894 18390 13954 18412
rect 14006 18390 14034 21442
rect 14278 21440 14298 21530
rect 14604 21440 14620 21530
rect 14278 21430 14620 21440
rect 13894 18354 14034 18390
rect 12764 18338 14034 18354
rect 12628 18228 13720 18284
rect 13664 15206 13720 18228
rect 13934 17780 14034 18338
rect 13934 17604 14034 17614
rect 14506 15290 14600 21430
rect 14980 21075 15066 21788
rect 14819 20989 15066 21075
rect 14820 15738 14906 20989
rect 14820 15643 14946 15738
rect 14505 15216 14826 15290
rect 10452 15150 13720 15206
rect 2950 12199 3016 12639
rect 7040 12496 7240 12568
rect 7040 12402 7240 12410
rect 14752 12020 14826 15216
rect 14870 12310 14946 15643
rect 14870 12302 15368 12310
rect 14870 12204 14878 12302
rect 15354 12204 15368 12302
rect 14870 12194 15368 12204
rect 15528 12302 15888 12312
rect 15528 12200 15540 12302
rect 15876 12200 15888 12302
rect 15528 12192 15888 12200
rect 14752 11943 15332 12020
rect 9694 11800 15210 11818
rect 9694 11796 9802 11800
rect 9694 6706 9708 11796
rect 9746 11764 9802 11796
rect 15110 11796 15210 11800
rect 15110 11764 15154 11796
rect 9746 11750 15154 11764
rect 9746 6706 9762 11750
rect 9836 11224 10072 11656
rect 10168 11224 10404 11656
rect 10500 11224 10736 11656
rect 10832 11224 11068 11656
rect 11164 11224 11400 11656
rect 11496 11224 11732 11656
rect 11828 11224 12064 11656
rect 12160 11224 12396 11656
rect 12492 11224 12728 11656
rect 12824 11224 13060 11656
rect 13156 11224 13392 11656
rect 13488 11224 13724 11656
rect 13820 11224 14056 11656
rect 14152 11224 14388 11656
rect 14484 11224 14720 11656
rect 14816 11224 15052 11656
rect 9694 6680 9762 6706
rect 9830 6656 9912 7260
rect 10002 6824 10238 7256
rect 10334 6824 10570 7256
rect 10666 6824 10902 7256
rect 10998 6824 11234 7256
rect 11330 6824 11566 7256
rect 11662 6824 11898 7256
rect 11994 6824 12230 7256
rect 12326 6824 12562 7256
rect 12658 6824 12894 7256
rect 12990 6824 13226 7256
rect 13322 6824 13558 7256
rect 13654 6824 13890 7256
rect 13986 6824 14222 7256
rect 14318 6824 14554 7256
rect 14650 6824 14886 7256
rect 10012 6730 14912 6748
rect 10012 6694 10038 6730
rect 14892 6694 14912 6730
rect 10012 6680 14912 6694
rect 9820 6646 9948 6656
rect 9820 6310 9832 6646
rect 9938 6310 9948 6646
rect 14980 6439 15052 7256
rect 15142 6700 15154 11750
rect 15198 6700 15210 11796
rect 15142 6682 15210 6700
rect 15254 6439 15332 11943
rect 14561 6361 15332 6439
rect 9820 6298 9948 6310
rect 14562 5486 14618 6361
rect 15542 6091 15634 12192
rect 10382 5430 14618 5486
rect 14976 6021 15634 6091
rect 2948 2437 3014 3119
rect 7038 2762 7238 2848
rect 7038 2684 7238 2694
rect 14976 2598 15042 6021
rect 14880 2590 15192 2598
rect 14880 2522 14894 2590
rect 15184 2522 15192 2590
rect 14880 2514 15192 2522
rect 7036 -6976 7236 -6900
rect 2536 -7000 2802 -6990
rect 2536 -7178 2550 -7000
rect 466 -7194 2550 -7178
rect 2792 -7178 2802 -7000
rect 7036 -7042 7046 -6976
rect 7328 -7042 7338 -6976
rect 7600 -7070 7800 -6862
rect 14978 -6886 15042 2514
rect 11578 -6950 15042 -6886
rect 7926 -7042 7942 -6976
rect 8264 -6978 8280 -6976
rect 11578 -6978 11642 -6950
rect 8264 -7042 11642 -6978
rect 13850 -7006 14474 -6994
rect 13850 -7070 13868 -7006
rect 7600 -7110 13868 -7070
rect 14454 -7058 14474 -7006
rect 14454 -7110 14856 -7058
rect 7600 -7142 14856 -7110
rect 2792 -7194 14710 -7178
rect 466 -7242 594 -7194
rect 14694 -7242 14710 -7194
rect 466 -7244 2550 -7242
rect 2792 -7244 14710 -7242
rect 466 -7254 14710 -7244
rect 466 -7340 566 -7254
rect 466 -9354 494 -7340
rect 466 -10500 480 -9354
rect 466 -11166 494 -10500
rect 548 -11166 566 -7340
rect 662 -7346 732 -7334
rect 14772 -7338 14856 -7142
rect 14916 -7194 29290 -7178
rect 14916 -7234 14944 -7194
rect 29200 -7234 29290 -7194
rect 14916 -7254 29290 -7234
rect 29214 -7278 29290 -7254
rect 662 -7770 732 -7756
rect 828 -7770 1064 -7338
rect 1160 -7770 1396 -7338
rect 1492 -7770 1728 -7338
rect 1824 -7770 2060 -7338
rect 2156 -7770 2392 -7338
rect 2488 -7770 2724 -7338
rect 2820 -7770 3056 -7338
rect 3152 -7770 3388 -7338
rect 3484 -7770 3720 -7338
rect 3816 -7770 4052 -7338
rect 4148 -7770 4384 -7338
rect 4480 -7770 4716 -7338
rect 4812 -7770 5048 -7338
rect 5144 -7770 5380 -7338
rect 5476 -7770 5712 -7338
rect 5808 -7770 6044 -7338
rect 6140 -7770 6376 -7338
rect 6472 -7770 6708 -7338
rect 6804 -7770 7040 -7338
rect 7136 -7770 7372 -7338
rect 7468 -7770 7704 -7338
rect 7800 -7770 8036 -7338
rect 8132 -7770 8368 -7338
rect 8464 -7770 8700 -7338
rect 8796 -7770 9032 -7338
rect 9128 -7770 9364 -7338
rect 9460 -7770 9696 -7338
rect 9792 -7770 10028 -7338
rect 10124 -7770 10360 -7338
rect 10456 -7770 10692 -7338
rect 10788 -7770 11024 -7338
rect 11120 -7770 11356 -7338
rect 11452 -7770 11688 -7338
rect 11784 -7770 12020 -7338
rect 12116 -7770 12352 -7338
rect 12448 -7770 12684 -7338
rect 12780 -7770 13016 -7338
rect 13112 -7770 13348 -7338
rect 13444 -7770 13680 -7338
rect 13776 -7770 14012 -7338
rect 14108 -7770 14344 -7338
rect 14440 -7770 14676 -7338
rect 14772 -7770 15008 -7338
rect 15104 -7770 15340 -7338
rect 15436 -7770 15672 -7338
rect 15768 -7770 16004 -7338
rect 16100 -7770 16336 -7338
rect 16432 -7770 16668 -7338
rect 16764 -7770 17000 -7338
rect 17096 -7770 17332 -7338
rect 17428 -7770 17664 -7338
rect 17760 -7770 17996 -7338
rect 18092 -7770 18328 -7338
rect 18424 -7770 18660 -7338
rect 18756 -7770 18992 -7338
rect 19088 -7770 19324 -7338
rect 19420 -7770 19656 -7338
rect 19752 -7770 19988 -7338
rect 20084 -7770 20320 -7338
rect 20416 -7770 20652 -7338
rect 20748 -7770 20984 -7338
rect 21080 -7770 21316 -7338
rect 21412 -7770 21648 -7338
rect 21744 -7770 21980 -7338
rect 22076 -7770 22312 -7338
rect 22408 -7770 22644 -7338
rect 22740 -7770 22976 -7338
rect 23072 -7770 23308 -7338
rect 23404 -7770 23640 -7338
rect 23736 -7770 23972 -7338
rect 24068 -7770 24304 -7338
rect 24400 -7770 24636 -7338
rect 24732 -7770 24968 -7338
rect 25064 -7770 25300 -7338
rect 25396 -7770 25632 -7338
rect 25728 -7770 25964 -7338
rect 26060 -7770 26296 -7338
rect 26392 -7770 26628 -7338
rect 26724 -7770 26960 -7338
rect 27056 -7770 27292 -7338
rect 27388 -7770 27624 -7338
rect 27720 -7770 27956 -7338
rect 28052 -7770 28288 -7338
rect 28384 -7770 28620 -7338
rect 28716 -7770 28952 -7338
rect 29048 -7350 29118 -7312
rect 29048 -7770 29118 -7756
rect 29214 -9360 29238 -7278
rect 29274 -9360 29290 -7278
rect 29214 -10498 29224 -9360
rect 29278 -10498 29290 -9360
rect 662 -11110 898 -10678
rect 994 -11110 1230 -10678
rect 1326 -11110 1562 -10678
rect 1658 -11110 1894 -10678
rect 1990 -11110 2226 -10678
rect 2322 -11110 2558 -10678
rect 2654 -11110 2890 -10678
rect 2986 -11110 3222 -10678
rect 3318 -11110 3554 -10678
rect 3650 -11110 3886 -10678
rect 3982 -11110 4218 -10678
rect 4314 -11110 4550 -10678
rect 4646 -11110 4882 -10678
rect 4978 -11110 5214 -10678
rect 5310 -11110 5546 -10678
rect 5642 -11110 5878 -10678
rect 5974 -11110 6210 -10678
rect 6306 -11110 6542 -10678
rect 6638 -11110 6874 -10678
rect 6970 -11110 7206 -10678
rect 7302 -11110 7538 -10678
rect 7634 -11110 7870 -10678
rect 7966 -11110 8202 -10678
rect 8298 -11110 8534 -10678
rect 8630 -11110 8866 -10678
rect 8962 -11110 9198 -10678
rect 9294 -11110 9530 -10678
rect 9626 -11110 9862 -10678
rect 9958 -11110 10194 -10678
rect 10290 -11110 10526 -10678
rect 10622 -11110 10858 -10678
rect 10954 -11110 11190 -10678
rect 11286 -11110 11522 -10678
rect 11618 -11110 11854 -10678
rect 11950 -11110 12186 -10678
rect 12282 -11110 12518 -10678
rect 12614 -11110 12850 -10678
rect 12946 -11110 13182 -10678
rect 13278 -11110 13514 -10678
rect 13610 -11110 13846 -10678
rect 13942 -11110 14178 -10678
rect 14274 -11110 14510 -10678
rect 14606 -11110 14842 -10678
rect 14938 -11110 15174 -10678
rect 15270 -11110 15506 -10678
rect 15602 -11110 15838 -10678
rect 15934 -11110 16170 -10678
rect 16266 -11110 16502 -10678
rect 16598 -11110 16834 -10678
rect 16930 -11110 17166 -10678
rect 17262 -11110 17498 -10678
rect 17594 -11110 17830 -10678
rect 17926 -11110 18162 -10678
rect 18258 -11110 18494 -10678
rect 18590 -11110 18826 -10678
rect 18922 -11110 19158 -10678
rect 19254 -11110 19490 -10678
rect 19586 -11110 19822 -10678
rect 19918 -11110 20154 -10678
rect 20250 -11110 20486 -10678
rect 20582 -11110 20818 -10678
rect 20914 -11110 21150 -10678
rect 21246 -11110 21482 -10678
rect 21578 -11110 21814 -10678
rect 21910 -11110 22146 -10678
rect 22242 -11110 22478 -10678
rect 22574 -11110 22810 -10678
rect 22906 -11110 23142 -10678
rect 23238 -11110 23474 -10678
rect 23570 -11110 23806 -10678
rect 23902 -11110 24138 -10678
rect 24234 -11110 24470 -10678
rect 24566 -11110 24802 -10678
rect 24898 -11110 25134 -10678
rect 25230 -11110 25466 -10678
rect 25562 -11110 25798 -10678
rect 25894 -11110 26130 -10678
rect 26226 -11110 26462 -10678
rect 26558 -11110 26794 -10678
rect 26890 -11110 27126 -10678
rect 27222 -11110 27458 -10678
rect 27554 -11110 27790 -10678
rect 27886 -11110 28122 -10678
rect 28218 -11110 28454 -10678
rect 28550 -11110 28786 -10678
rect 28882 -11110 29118 -10678
rect 466 -11206 566 -11166
rect 29214 -11182 29238 -10498
rect 29274 -11182 29290 -10498
rect 29214 -11206 29290 -11182
rect 466 -11228 29290 -11206
rect 466 -11276 594 -11228
rect 29198 -11276 29290 -11228
rect 466 -11294 29290 -11276
<< via1 >>
rect 384 26054 598 26198
rect 652 22010 1056 22102
rect 11190 22124 11350 22280
rect 12152 22116 12260 22288
rect 9716 21664 9872 21916
rect 12786 21930 12952 22100
rect 22808 22012 23086 22104
rect 14472 21788 14672 21912
rect 12782 21604 12962 21710
rect 10654 21466 11010 21552
rect 11018 21278 11314 21392
rect 14728 21610 14908 21728
rect 14298 21440 14604 21530
rect 13934 17614 14034 17780
rect 7040 12410 7240 12496
rect 14878 12204 15354 12302
rect 15540 12200 15876 12302
rect 9832 6310 9938 6646
rect 7038 2694 7238 2762
rect 14894 2522 15184 2590
rect 2550 -7194 2792 -7000
rect 7046 -7042 7328 -6976
rect 7942 -7042 8264 -6976
rect 13868 -7110 14454 -7006
rect 2550 -7242 2792 -7194
rect 2550 -7244 2792 -7242
rect 480 -10500 494 -9354
rect 494 -10500 540 -9354
rect 662 -7756 732 -7346
rect 29048 -7756 29118 -7350
rect 29224 -10498 29238 -9360
rect 29238 -10498 29274 -9360
rect 29274 -10498 29278 -9360
<< metal2 >>
rect 1028 28058 1228 28258
rect 3428 28058 3628 28258
rect 5828 28058 6028 28258
rect 8228 28058 8428 28258
rect 10628 28058 10828 28258
rect 13028 28058 13228 28258
rect 15428 28058 15628 28258
rect 17828 28058 18028 28258
rect 20228 28058 20428 28258
rect 22628 28058 22828 28258
rect 384 26198 598 26216
rect 384 21234 598 26054
rect 2718 22546 2922 22568
rect 2718 22390 2740 22546
rect 2902 22390 2922 22546
rect 2718 22372 2922 22390
rect 5118 22546 5322 22568
rect 5118 22390 5140 22546
rect 5302 22390 5322 22546
rect 5118 22372 5322 22390
rect 7518 22546 7722 22568
rect 7518 22390 7540 22546
rect 7702 22390 7722 22546
rect 7518 22372 7722 22390
rect 9918 22546 10122 22568
rect 9918 22390 9940 22546
rect 10102 22390 10122 22546
rect 9918 22372 10122 22390
rect 12318 22546 12522 22568
rect 12318 22390 12340 22546
rect 12502 22390 12522 22546
rect 12318 22372 12522 22390
rect 14718 22546 14922 22568
rect 14718 22390 14740 22546
rect 14902 22390 14922 22546
rect 14718 22372 14922 22390
rect 17118 22546 17322 22568
rect 17118 22390 17140 22546
rect 17302 22390 17322 22546
rect 17118 22372 17322 22390
rect 19518 22546 19722 22568
rect 19518 22390 19540 22546
rect 19702 22390 19722 22546
rect 19518 22372 19722 22390
rect 21918 22546 22122 22568
rect 21918 22390 21940 22546
rect 22102 22390 22122 22546
rect 21918 22372 22122 22390
rect 24318 22546 24522 22568
rect 24318 22390 24340 22546
rect 24502 22390 24522 22546
rect 24318 22372 24522 22390
rect 2472 22280 2676 22300
rect 2472 22124 2494 22280
rect 2654 22124 2676 22280
rect 638 22102 1072 22116
rect 2472 22104 2676 22124
rect 4872 22280 5076 22300
rect 4872 22124 4894 22280
rect 5054 22124 5076 22280
rect 4872 22104 5076 22124
rect 7272 22280 7476 22300
rect 7272 22124 7294 22280
rect 7454 22124 7476 22280
rect 7272 22104 7476 22124
rect 9672 22280 9876 22300
rect 9672 22124 9694 22280
rect 9854 22124 9876 22280
rect 9672 22104 9876 22124
rect 11168 22280 11372 22300
rect 11168 22124 11190 22280
rect 11350 22124 11372 22280
rect 11168 22104 11372 22124
rect 12072 22288 12276 22300
rect 12072 22280 12152 22288
rect 12072 22124 12094 22280
rect 12072 22116 12152 22124
rect 12260 22116 12276 22288
rect 12072 22104 12276 22116
rect 14472 22280 14676 22300
rect 14472 22122 14494 22280
rect 14654 22178 14676 22280
rect 16872 22280 17076 22300
rect 14654 22122 14674 22178
rect 638 22010 652 22102
rect 1056 22010 1072 22102
rect 638 21996 1072 22010
rect 12770 22100 12968 22114
rect 9308 21916 12502 21940
rect 12770 21930 12786 22100
rect 12952 21930 12968 22100
rect 12770 21920 12968 21930
rect 9308 21664 9716 21916
rect 9872 21664 12502 21916
rect 9308 21638 12502 21664
rect 12768 21720 12968 21920
rect 14472 22104 14674 22122
rect 16872 22124 16894 22280
rect 17054 22124 17076 22280
rect 16872 22104 17076 22124
rect 19272 22280 19476 22300
rect 19272 22124 19294 22280
rect 19454 22124 19476 22280
rect 19272 22104 19476 22124
rect 21672 22280 21876 22300
rect 21672 22124 21694 22280
rect 21854 22124 21876 22280
rect 21672 22104 21876 22124
rect 24072 22280 24276 22300
rect 24072 22124 24094 22280
rect 24254 22124 24276 22280
rect 22798 22104 23100 22114
rect 24072 22104 24276 22124
rect 14472 21912 14672 22104
rect 22798 22072 22808 22104
rect 14472 21774 14672 21788
rect 14728 22012 22808 22072
rect 23086 22012 23100 22104
rect 14728 21996 23100 22012
rect 14728 21728 14908 21996
rect 12768 21710 12972 21720
rect 12768 21604 12782 21710
rect 12962 21604 12972 21710
rect 12768 21594 12972 21604
rect 14728 21598 14908 21610
rect 10642 21552 11024 21562
rect 10642 21466 10654 21552
rect 11010 21542 11024 21552
rect 14278 21542 14620 21546
rect 11010 21530 14620 21542
rect 11010 21466 14298 21530
rect 10642 21456 14298 21466
rect 14278 21440 14298 21456
rect 14604 21440 14620 21530
rect 14278 21430 14620 21440
rect 11002 21392 11332 21408
rect 11002 21278 11018 21392
rect 11314 21346 11332 21392
rect 14894 21346 15094 21466
rect 11314 21278 15094 21346
rect 11002 21266 15094 21278
rect 14978 21058 15094 21266
rect 9320 17614 13934 17780
rect 14034 17614 14049 17780
rect 7027 12410 7040 12496
rect 7240 12410 14684 12496
rect 364 12370 490 12380
rect 364 12270 376 12370
rect 480 12354 490 12370
rect 480 12346 14392 12354
rect 480 12274 14194 12346
rect 480 12270 490 12274
rect 364 12256 490 12270
rect 14178 12154 14194 12274
rect 14382 12154 14392 12346
rect 14590 12300 14684 12410
rect 14870 12304 15368 12310
rect 15528 12304 15888 12312
rect 14870 12302 15888 12304
rect 14870 12300 14878 12302
rect 14590 12212 14878 12300
rect 14870 12204 14878 12212
rect 15354 12204 15540 12302
rect 14870 12194 15368 12204
rect 15528 12200 15540 12204
rect 15876 12200 15888 12302
rect 15528 12192 15888 12200
rect 14178 12142 14392 12154
rect 14646 12130 14870 12138
rect 9306 11748 14474 12062
rect 14646 11884 14656 12130
rect 14858 11884 14870 12130
rect 14646 11876 14870 11884
rect 7018 2694 7038 2762
rect 7238 2694 14498 2762
rect 14430 2598 14498 2694
rect 14430 2590 15192 2598
rect 14430 2530 14894 2590
rect 14880 2522 14894 2530
rect 15184 2522 15192 2590
rect 14880 2514 15192 2522
rect 2536 -7000 2802 -6990
rect 2536 -7244 2550 -7000
rect 2792 -7244 2802 -7000
rect 7036 -7042 7046 -6976
rect 7328 -7042 7942 -6976
rect 8264 -7042 8280 -6976
rect 13850 -7006 14474 -6994
rect 13850 -7110 13868 -7006
rect 14454 -7110 14474 -7006
rect 13850 -7124 14474 -7110
rect 14644 -7128 14662 -7016
rect 14860 -7042 14870 -7016
rect 14860 -7128 15206 -7042
rect 2536 -7254 2802 -7244
rect 15094 -7278 15206 -7128
rect 384 -7342 736 -7334
rect 384 -7756 394 -7342
rect 468 -7346 736 -7342
rect 468 -7756 662 -7346
rect 732 -7756 736 -7346
rect 15094 -7350 29138 -7278
rect 15094 -7390 29048 -7350
rect 384 -7770 736 -7756
rect 29036 -7756 29048 -7390
rect 29118 -7756 29138 -7350
rect 29036 -7770 29138 -7756
<< via2 >>
rect 2740 22390 2902 22546
rect 5140 22390 5302 22546
rect 7540 22390 7702 22546
rect 9940 22390 10102 22546
rect 12340 22390 12502 22546
rect 14740 22390 14902 22546
rect 17140 22390 17302 22546
rect 19540 22390 19702 22546
rect 21940 22390 22102 22546
rect 24340 22390 24502 22546
rect 2494 22124 2654 22280
rect 4894 22124 5054 22280
rect 7294 22124 7454 22280
rect 9694 22124 9854 22280
rect 11190 22124 11350 22280
rect 12094 22124 12152 22280
rect 12152 22124 12254 22280
rect 14494 22122 14654 22280
rect 652 22010 1056 22102
rect 12786 21930 12952 22100
rect 16894 22124 17054 22280
rect 19294 22124 19454 22280
rect 21694 22124 21854 22280
rect 24094 22124 24254 22280
rect 376 12270 480 12370
rect 14194 12154 14382 12346
rect 14656 11884 14858 12130
rect 2550 -7244 2792 -7000
rect 13868 -7110 14454 -7006
rect 14662 -7128 14860 -7016
rect 394 -7756 468 -7342
<< metal3 >>
rect 2718 22546 2922 22568
rect 2718 22508 2740 22546
rect 670 22396 2740 22508
rect 2718 22390 2740 22396
rect 2902 22508 2922 22546
rect 5118 22546 5322 22568
rect 5118 22508 5140 22546
rect 2902 22396 5140 22508
rect 2902 22390 2922 22396
rect 2718 22372 2922 22390
rect 5118 22390 5140 22396
rect 5302 22508 5322 22546
rect 7518 22546 7722 22568
rect 7518 22508 7540 22546
rect 5302 22396 7540 22508
rect 5302 22390 5322 22396
rect 5118 22372 5322 22390
rect 7518 22390 7540 22396
rect 7702 22508 7722 22546
rect 9918 22546 10122 22568
rect 9918 22508 9940 22546
rect 7702 22396 9940 22508
rect 7702 22390 7722 22396
rect 7518 22372 7722 22390
rect 9918 22390 9940 22396
rect 10102 22508 10122 22546
rect 12318 22546 12522 22568
rect 12318 22508 12340 22546
rect 10102 22396 12340 22508
rect 10102 22390 10122 22396
rect 9918 22372 10122 22390
rect 12318 22390 12340 22396
rect 12502 22508 12522 22546
rect 14718 22546 14922 22568
rect 14718 22508 14740 22546
rect 12502 22396 14740 22508
rect 12502 22390 12522 22396
rect 12318 22372 12522 22390
rect 14718 22390 14740 22396
rect 14902 22508 14922 22546
rect 15002 22554 15572 22574
rect 15002 22508 15030 22554
rect 14902 22412 15030 22508
rect 15548 22508 15572 22554
rect 17118 22546 17322 22568
rect 17118 22508 17140 22546
rect 15548 22412 17140 22508
rect 14902 22396 17140 22412
rect 14902 22390 14922 22396
rect 14718 22372 14922 22390
rect 17118 22390 17140 22396
rect 17302 22508 17322 22546
rect 19518 22546 19722 22568
rect 19518 22508 19540 22546
rect 17302 22396 19540 22508
rect 17302 22390 17322 22396
rect 17118 22372 17322 22390
rect 19518 22390 19540 22396
rect 19702 22508 19722 22546
rect 21918 22546 22122 22568
rect 21918 22508 21940 22546
rect 19702 22396 21940 22508
rect 19702 22390 19722 22396
rect 19518 22372 19722 22390
rect 21918 22390 21940 22396
rect 22102 22508 22122 22546
rect 24318 22546 24522 22568
rect 24318 22508 24340 22546
rect 22102 22396 24340 22508
rect 22102 22390 22122 22396
rect 21918 22372 22122 22390
rect 24318 22390 24340 22396
rect 24502 22508 24522 22546
rect 24502 22396 24664 22508
rect 24502 22390 24522 22396
rect 24318 22372 24522 22390
rect 2472 22290 2676 22300
rect 4872 22290 5076 22300
rect 7272 22290 7476 22300
rect 9672 22290 9876 22300
rect 11168 22290 11372 22300
rect 12072 22290 12276 22300
rect 14472 22290 14676 22300
rect 16872 22290 17076 22300
rect 19272 22290 19476 22300
rect 21672 22290 21876 22300
rect 24072 22290 24276 22300
rect 672 22280 24774 22290
rect 672 22178 2494 22280
rect 2472 22124 2494 22178
rect 2654 22178 4894 22280
rect 2654 22124 2676 22178
rect 636 22102 1072 22116
rect 2472 22104 2676 22124
rect 4872 22124 4894 22178
rect 5054 22178 7294 22280
rect 5054 22124 5076 22178
rect 4872 22104 5076 22124
rect 7272 22124 7294 22178
rect 7454 22178 9694 22280
rect 7454 22124 7476 22178
rect 7272 22104 7476 22124
rect 9672 22124 9694 22178
rect 9854 22178 11190 22280
rect 9854 22124 9876 22178
rect 9672 22104 9876 22124
rect 11168 22124 11190 22178
rect 11350 22178 12094 22280
rect 11350 22124 11372 22178
rect 11168 22104 11372 22124
rect 12072 22124 12094 22178
rect 12254 22178 14494 22280
rect 12254 22124 12276 22178
rect 12072 22104 12276 22124
rect 14472 22122 14494 22178
rect 14654 22178 16894 22280
rect 14654 22122 14676 22178
rect 636 22010 652 22102
rect 1056 22010 1072 22102
rect 636 21996 1072 22010
rect 12770 22100 12968 22114
rect 14472 22104 14676 22122
rect 16872 22124 16894 22178
rect 17054 22178 19294 22280
rect 17054 22124 17076 22178
rect 16872 22104 17076 22124
rect 19272 22124 19294 22178
rect 19454 22178 21694 22280
rect 19454 22124 19476 22178
rect 19272 22104 19476 22124
rect 21672 22124 21694 22178
rect 21854 22178 24094 22280
rect 21854 22124 21876 22178
rect 21672 22104 21876 22124
rect 24072 22124 24094 22178
rect 24254 22178 24774 22280
rect 24254 22124 24276 22178
rect 24072 22104 24276 22124
rect 12770 21930 12786 22100
rect 12952 22038 12968 22100
rect 24574 22090 24774 22178
rect 12952 21948 14870 22038
rect 12952 21930 12968 21948
rect 12770 21914 12968 21930
rect 726 21686 926 21886
rect 14658 21092 14870 21948
rect 2578 20814 2778 21014
rect 364 12370 490 12380
rect 364 12270 376 12370
rect 480 12270 490 12370
rect 364 12256 490 12270
rect 386 -7342 474 12256
rect 574 12216 1074 12564
rect 2538 12222 2808 13782
rect 14658 12490 14870 14044
rect 14180 12346 14870 12490
rect 14180 12154 14194 12346
rect 14382 12278 14870 12346
rect 14382 12154 14392 12278
rect 14180 12142 14392 12154
rect 14646 12130 14870 12138
rect 14646 11884 14656 12130
rect 14858 11884 14870 12130
rect 14646 11876 14870 11884
rect 14656 11378 14868 11876
rect 572 2454 1072 2850
rect 2536 2472 2806 4058
rect 386 -7756 394 -7342
rect 468 -7756 474 -7342
rect 386 -7770 474 -7756
rect 572 -11250 1072 -6892
rect 2534 -7000 2804 -5680
rect 2534 -7244 2550 -7000
rect 2792 -7244 2804 -7000
rect 13850 -7006 14474 -6994
rect 13850 -7110 13868 -7006
rect 14454 -7110 14474 -7006
rect 13850 -7124 14474 -7110
rect 14654 -7016 14866 -5412
rect 2534 -11244 2804 -7244
rect 14654 -7128 14662 -7016
rect 14860 -7128 14866 -7016
rect 14654 -11384 14866 -7128
<< via3 >>
rect 15030 22412 15548 22554
rect 652 22010 1056 22102
rect 14660 11886 14856 12124
rect 13868 -7110 14454 -7006
<< metal4 >>
rect 15002 22554 15572 22574
rect 15002 22412 15030 22554
rect 15548 22412 15572 22554
rect 15002 22396 15572 22412
rect 636 22102 1072 22116
rect 636 22010 652 22102
rect 1056 22096 1072 22102
rect 1056 22014 14900 22096
rect 1056 22010 1072 22014
rect 636 21996 1072 22010
rect 14784 12504 14900 22014
rect 14646 12280 14900 12504
rect 14646 12124 14870 12280
rect 14646 11886 14660 12124
rect 14856 11886 14870 12124
rect 14646 11876 14870 11886
rect 15002 -6994 15122 22396
rect 13850 -7006 15122 -6994
rect 13850 -7110 13868 -7006
rect 14454 -7110 15122 -7006
rect 13850 -7124 15122 -7110
<< comment >>
rect 14868 -10456 14928 -7948
use sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP  sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP_0 paramcells
timestamp 1730948043
transform 1 0 13390 0 1 19922
box -616 -1582 616 1582
use sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP  sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP_1
timestamp 1730948043
transform 1 0 10430 0 1 19922
box -616 -1582 616 1582
use sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP  sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP_2
timestamp 1730948043
transform 1 0 11910 0 1 19922
box -616 -1582 616 1582
use sky130_fd_pr__res_xhigh_po_0p35_QDMB52  sky130_fd_pr__res_xhigh_po_0p35_QDMB52_0 paramcells
timestamp 1730948043
transform 1 0 14890 0 1 -9224
box -14394 -2052 14394 2052
use sky130_fd_pr__res_xhigh_po_0p35_S4N9LQ  sky130_fd_pr__res_xhigh_po_0p35_S4N9LQ_0 paramcells
timestamp 1730948043
transform 1 0 12444 0 1 9240
box -2774 -2582 2774 2582
use Universal_R_2R_Block2  x1
timestamp 1730948043
transform 0 1 22546 -1 0 29868
box 1610 -2778 7848 -198
use Universal_R_2R_Block2  x2
timestamp 1730948043
transform 0 1 15346 -1 0 29868
box 1610 -2778 7848 -198
use Universal_R_2R_Block2  x3
timestamp 1730948043
transform 0 1 8146 -1 0 29868
box 1610 -2778 7848 -198
use Universal_R_2R_Block2  x4
timestamp 1730948043
transform 0 1 3346 -1 0 29868
box 1610 -2778 7848 -198
use Universal_R_2R_Block2  x5
timestamp 1730948043
transform 0 1 17746 -1 0 29868
box 1610 -2778 7848 -198
use x1_x32_OA  x6
timestamp 1730948043
transform -1 0 15498 0 1 13652
box 548 -1232 15090 8401
use Output_OA  x7
timestamp 1730948043
transform -1 0 15494 0 1 -5816
box 548 -1234 15090 8401
use x1_x32_OA  x8
timestamp 1730948043
transform -1 0 15496 0 1 3932
box 548 -1232 15090 8401
use Universal_R_2R_Block2  x9
timestamp 1730948043
transform 0 1 12946 -1 0 29868
box 1610 -2778 7848 -198
use Universal_R_2R_Block2  x10
timestamp 1730948043
transform 0 1 10546 -1 0 29868
box 1610 -2778 7848 -198
use Universal_R_2R_Block2  x11
timestamp 1730948043
transform 0 1 5746 -1 0 29868
box 1610 -2778 7848 -198
use Universal_R_2R_Block2  x12
timestamp 1730948043
transform 0 1 20146 -1 0 29868
box 1610 -2778 7848 -198
use Universal_R_2R_Block2  x13
timestamp 1730948043
transform 0 1 24946 -1 0 29868
box 1610 -2778 7848 -198
<< labels >>
flabel metal1 2816 21760 3016 21960 0 FreeSans 256 0 0 0 VBIAS
port 17 nsew
flabel metal3 14660 -11380 14860 -11180 0 FreeSans 256 0 0 0 VOUT
port 8 nsew
flabel metal2 22628 28058 22828 28258 0 FreeSans 256 270 0 0 V9
port 3 nsew
flabel metal2 20228 28058 20428 28258 0 FreeSans 256 270 0 0 V8
port 2 nsew
flabel metal2 17828 28058 18028 28258 0 FreeSans 256 270 0 0 V7
port 4 nsew
flabel metal2 15428 28058 15628 28258 0 FreeSans 256 270 0 0 V6
port 0 nsew
flabel metal2 13028 28058 13228 28258 0 FreeSans 256 270 0 0 V5
port 1 nsew
flabel metal2 10628 28058 10828 28258 0 FreeSans 256 270 0 0 V4
port 9 nsew
flabel metal2 8228 28058 8428 28258 0 FreeSans 256 270 0 0 V3
port 10 nsew
flabel metal2 5828 28058 6028 28258 0 FreeSans 256 270 0 0 V2
port 11 nsew
flabel metal2 3428 28058 3628 28258 0 FreeSans 256 270 0 0 V1
port 12 nsew
flabel metal2 1028 28058 1228 28258 0 FreeSans 256 270 0 0 V0
port 13 nsew
flabel metal2 14894 21266 15094 21466 0 FreeSans 256 0 0 0 VO1
port 5 nsew
flabel metal3 24574 22090 24774 22290 0 FreeSans 256 0 0 0 VCM
port 14 nsew
flabel metal3 2578 20814 2778 21014 0 FreeSans 256 0 0 0 AVSS
port 16 nsew
flabel metal3 726 21686 926 21886 0 FreeSans 256 0 0 0 AVDD
port 7 nsew
flabel metal1 24626 27546 24826 27746 0 FreeSans 256 0 0 0 DVDD
port 6 nsew
flabel metal1 24648 28030 24848 28230 0 FreeSans 256 0 0 0 DVSS
port 15 nsew
<< end >>
