magic
tech sky130A
timestamp 1730992408
<< pwell >>
rect -1583 -1489 1583 1489
<< mvnmos >>
rect -1469 860 -1369 1360
rect -1340 860 -1240 1360
rect -1211 860 -1111 1360
rect -1082 860 -982 1360
rect -953 860 -853 1360
rect -824 860 -724 1360
rect -695 860 -595 1360
rect -566 860 -466 1360
rect -437 860 -337 1360
rect -308 860 -208 1360
rect -179 860 -79 1360
rect -50 860 50 1360
rect 79 860 179 1360
rect 208 860 308 1360
rect 337 860 437 1360
rect 466 860 566 1360
rect 595 860 695 1360
rect 724 860 824 1360
rect 853 860 953 1360
rect 982 860 1082 1360
rect 1111 860 1211 1360
rect 1240 860 1340 1360
rect 1369 860 1469 1360
rect -1469 305 -1369 805
rect -1340 305 -1240 805
rect -1211 305 -1111 805
rect -1082 305 -982 805
rect -953 305 -853 805
rect -824 305 -724 805
rect -695 305 -595 805
rect -566 305 -466 805
rect -437 305 -337 805
rect -308 305 -208 805
rect -179 305 -79 805
rect -50 305 50 805
rect 79 305 179 805
rect 208 305 308 805
rect 337 305 437 805
rect 466 305 566 805
rect 595 305 695 805
rect 724 305 824 805
rect 853 305 953 805
rect 982 305 1082 805
rect 1111 305 1211 805
rect 1240 305 1340 805
rect 1369 305 1469 805
rect -1469 -250 -1369 250
rect -1340 -250 -1240 250
rect -1211 -250 -1111 250
rect -1082 -250 -982 250
rect -953 -250 -853 250
rect -824 -250 -724 250
rect -695 -250 -595 250
rect -566 -250 -466 250
rect -437 -250 -337 250
rect -308 -250 -208 250
rect -179 -250 -79 250
rect -50 -250 50 250
rect 79 -250 179 250
rect 208 -250 308 250
rect 337 -250 437 250
rect 466 -250 566 250
rect 595 -250 695 250
rect 724 -250 824 250
rect 853 -250 953 250
rect 982 -250 1082 250
rect 1111 -250 1211 250
rect 1240 -250 1340 250
rect 1369 -250 1469 250
rect -1469 -805 -1369 -305
rect -1340 -805 -1240 -305
rect -1211 -805 -1111 -305
rect -1082 -805 -982 -305
rect -953 -805 -853 -305
rect -824 -805 -724 -305
rect -695 -805 -595 -305
rect -566 -805 -466 -305
rect -437 -805 -337 -305
rect -308 -805 -208 -305
rect -179 -805 -79 -305
rect -50 -805 50 -305
rect 79 -805 179 -305
rect 208 -805 308 -305
rect 337 -805 437 -305
rect 466 -805 566 -305
rect 595 -805 695 -305
rect 724 -805 824 -305
rect 853 -805 953 -305
rect 982 -805 1082 -305
rect 1111 -805 1211 -305
rect 1240 -805 1340 -305
rect 1369 -805 1469 -305
rect -1469 -1360 -1369 -860
rect -1340 -1360 -1240 -860
rect -1211 -1360 -1111 -860
rect -1082 -1360 -982 -860
rect -953 -1360 -853 -860
rect -824 -1360 -724 -860
rect -695 -1360 -595 -860
rect -566 -1360 -466 -860
rect -437 -1360 -337 -860
rect -308 -1360 -208 -860
rect -179 -1360 -79 -860
rect -50 -1360 50 -860
rect 79 -1360 179 -860
rect 208 -1360 308 -860
rect 337 -1360 437 -860
rect 466 -1360 566 -860
rect 595 -1360 695 -860
rect 724 -1360 824 -860
rect 853 -1360 953 -860
rect 982 -1360 1082 -860
rect 1111 -1360 1211 -860
rect 1240 -1360 1340 -860
rect 1369 -1360 1469 -860
<< mvndiff >>
rect -1498 1354 -1469 1360
rect -1498 866 -1492 1354
rect -1475 866 -1469 1354
rect -1498 860 -1469 866
rect -1369 1354 -1340 1360
rect -1369 866 -1363 1354
rect -1346 866 -1340 1354
rect -1369 860 -1340 866
rect -1240 1354 -1211 1360
rect -1240 866 -1234 1354
rect -1217 866 -1211 1354
rect -1240 860 -1211 866
rect -1111 1354 -1082 1360
rect -1111 866 -1105 1354
rect -1088 866 -1082 1354
rect -1111 860 -1082 866
rect -982 1354 -953 1360
rect -982 866 -976 1354
rect -959 866 -953 1354
rect -982 860 -953 866
rect -853 1354 -824 1360
rect -853 866 -847 1354
rect -830 866 -824 1354
rect -853 860 -824 866
rect -724 1354 -695 1360
rect -724 866 -718 1354
rect -701 866 -695 1354
rect -724 860 -695 866
rect -595 1354 -566 1360
rect -595 866 -589 1354
rect -572 866 -566 1354
rect -595 860 -566 866
rect -466 1354 -437 1360
rect -466 866 -460 1354
rect -443 866 -437 1354
rect -466 860 -437 866
rect -337 1354 -308 1360
rect -337 866 -331 1354
rect -314 866 -308 1354
rect -337 860 -308 866
rect -208 1354 -179 1360
rect -208 866 -202 1354
rect -185 866 -179 1354
rect -208 860 -179 866
rect -79 1354 -50 1360
rect -79 866 -73 1354
rect -56 866 -50 1354
rect -79 860 -50 866
rect 50 1354 79 1360
rect 50 866 56 1354
rect 73 866 79 1354
rect 50 860 79 866
rect 179 1354 208 1360
rect 179 866 185 1354
rect 202 866 208 1354
rect 179 860 208 866
rect 308 1354 337 1360
rect 308 866 314 1354
rect 331 866 337 1354
rect 308 860 337 866
rect 437 1354 466 1360
rect 437 866 443 1354
rect 460 866 466 1354
rect 437 860 466 866
rect 566 1354 595 1360
rect 566 866 572 1354
rect 589 866 595 1354
rect 566 860 595 866
rect 695 1354 724 1360
rect 695 866 701 1354
rect 718 866 724 1354
rect 695 860 724 866
rect 824 1354 853 1360
rect 824 866 830 1354
rect 847 866 853 1354
rect 824 860 853 866
rect 953 1354 982 1360
rect 953 866 959 1354
rect 976 866 982 1354
rect 953 860 982 866
rect 1082 1354 1111 1360
rect 1082 866 1088 1354
rect 1105 866 1111 1354
rect 1082 860 1111 866
rect 1211 1354 1240 1360
rect 1211 866 1217 1354
rect 1234 866 1240 1354
rect 1211 860 1240 866
rect 1340 1354 1369 1360
rect 1340 866 1346 1354
rect 1363 866 1369 1354
rect 1340 860 1369 866
rect 1469 1354 1498 1360
rect 1469 866 1475 1354
rect 1492 866 1498 1354
rect 1469 860 1498 866
rect -1498 799 -1469 805
rect -1498 311 -1492 799
rect -1475 311 -1469 799
rect -1498 305 -1469 311
rect -1369 799 -1340 805
rect -1369 311 -1363 799
rect -1346 311 -1340 799
rect -1369 305 -1340 311
rect -1240 799 -1211 805
rect -1240 311 -1234 799
rect -1217 311 -1211 799
rect -1240 305 -1211 311
rect -1111 799 -1082 805
rect -1111 311 -1105 799
rect -1088 311 -1082 799
rect -1111 305 -1082 311
rect -982 799 -953 805
rect -982 311 -976 799
rect -959 311 -953 799
rect -982 305 -953 311
rect -853 799 -824 805
rect -853 311 -847 799
rect -830 311 -824 799
rect -853 305 -824 311
rect -724 799 -695 805
rect -724 311 -718 799
rect -701 311 -695 799
rect -724 305 -695 311
rect -595 799 -566 805
rect -595 311 -589 799
rect -572 311 -566 799
rect -595 305 -566 311
rect -466 799 -437 805
rect -466 311 -460 799
rect -443 311 -437 799
rect -466 305 -437 311
rect -337 799 -308 805
rect -337 311 -331 799
rect -314 311 -308 799
rect -337 305 -308 311
rect -208 799 -179 805
rect -208 311 -202 799
rect -185 311 -179 799
rect -208 305 -179 311
rect -79 799 -50 805
rect -79 311 -73 799
rect -56 311 -50 799
rect -79 305 -50 311
rect 50 799 79 805
rect 50 311 56 799
rect 73 311 79 799
rect 50 305 79 311
rect 179 799 208 805
rect 179 311 185 799
rect 202 311 208 799
rect 179 305 208 311
rect 308 799 337 805
rect 308 311 314 799
rect 331 311 337 799
rect 308 305 337 311
rect 437 799 466 805
rect 437 311 443 799
rect 460 311 466 799
rect 437 305 466 311
rect 566 799 595 805
rect 566 311 572 799
rect 589 311 595 799
rect 566 305 595 311
rect 695 799 724 805
rect 695 311 701 799
rect 718 311 724 799
rect 695 305 724 311
rect 824 799 853 805
rect 824 311 830 799
rect 847 311 853 799
rect 824 305 853 311
rect 953 799 982 805
rect 953 311 959 799
rect 976 311 982 799
rect 953 305 982 311
rect 1082 799 1111 805
rect 1082 311 1088 799
rect 1105 311 1111 799
rect 1082 305 1111 311
rect 1211 799 1240 805
rect 1211 311 1217 799
rect 1234 311 1240 799
rect 1211 305 1240 311
rect 1340 799 1369 805
rect 1340 311 1346 799
rect 1363 311 1369 799
rect 1340 305 1369 311
rect 1469 799 1498 805
rect 1469 311 1475 799
rect 1492 311 1498 799
rect 1469 305 1498 311
rect -1498 244 -1469 250
rect -1498 -244 -1492 244
rect -1475 -244 -1469 244
rect -1498 -250 -1469 -244
rect -1369 244 -1340 250
rect -1369 -244 -1363 244
rect -1346 -244 -1340 244
rect -1369 -250 -1340 -244
rect -1240 244 -1211 250
rect -1240 -244 -1234 244
rect -1217 -244 -1211 244
rect -1240 -250 -1211 -244
rect -1111 244 -1082 250
rect -1111 -244 -1105 244
rect -1088 -244 -1082 244
rect -1111 -250 -1082 -244
rect -982 244 -953 250
rect -982 -244 -976 244
rect -959 -244 -953 244
rect -982 -250 -953 -244
rect -853 244 -824 250
rect -853 -244 -847 244
rect -830 -244 -824 244
rect -853 -250 -824 -244
rect -724 244 -695 250
rect -724 -244 -718 244
rect -701 -244 -695 244
rect -724 -250 -695 -244
rect -595 244 -566 250
rect -595 -244 -589 244
rect -572 -244 -566 244
rect -595 -250 -566 -244
rect -466 244 -437 250
rect -466 -244 -460 244
rect -443 -244 -437 244
rect -466 -250 -437 -244
rect -337 244 -308 250
rect -337 -244 -331 244
rect -314 -244 -308 244
rect -337 -250 -308 -244
rect -208 244 -179 250
rect -208 -244 -202 244
rect -185 -244 -179 244
rect -208 -250 -179 -244
rect -79 244 -50 250
rect -79 -244 -73 244
rect -56 -244 -50 244
rect -79 -250 -50 -244
rect 50 244 79 250
rect 50 -244 56 244
rect 73 -244 79 244
rect 50 -250 79 -244
rect 179 244 208 250
rect 179 -244 185 244
rect 202 -244 208 244
rect 179 -250 208 -244
rect 308 244 337 250
rect 308 -244 314 244
rect 331 -244 337 244
rect 308 -250 337 -244
rect 437 244 466 250
rect 437 -244 443 244
rect 460 -244 466 244
rect 437 -250 466 -244
rect 566 244 595 250
rect 566 -244 572 244
rect 589 -244 595 244
rect 566 -250 595 -244
rect 695 244 724 250
rect 695 -244 701 244
rect 718 -244 724 244
rect 695 -250 724 -244
rect 824 244 853 250
rect 824 -244 830 244
rect 847 -244 853 244
rect 824 -250 853 -244
rect 953 244 982 250
rect 953 -244 959 244
rect 976 -244 982 244
rect 953 -250 982 -244
rect 1082 244 1111 250
rect 1082 -244 1088 244
rect 1105 -244 1111 244
rect 1082 -250 1111 -244
rect 1211 244 1240 250
rect 1211 -244 1217 244
rect 1234 -244 1240 244
rect 1211 -250 1240 -244
rect 1340 244 1369 250
rect 1340 -244 1346 244
rect 1363 -244 1369 244
rect 1340 -250 1369 -244
rect 1469 244 1498 250
rect 1469 -244 1475 244
rect 1492 -244 1498 244
rect 1469 -250 1498 -244
rect -1498 -311 -1469 -305
rect -1498 -799 -1492 -311
rect -1475 -799 -1469 -311
rect -1498 -805 -1469 -799
rect -1369 -311 -1340 -305
rect -1369 -799 -1363 -311
rect -1346 -799 -1340 -311
rect -1369 -805 -1340 -799
rect -1240 -311 -1211 -305
rect -1240 -799 -1234 -311
rect -1217 -799 -1211 -311
rect -1240 -805 -1211 -799
rect -1111 -311 -1082 -305
rect -1111 -799 -1105 -311
rect -1088 -799 -1082 -311
rect -1111 -805 -1082 -799
rect -982 -311 -953 -305
rect -982 -799 -976 -311
rect -959 -799 -953 -311
rect -982 -805 -953 -799
rect -853 -311 -824 -305
rect -853 -799 -847 -311
rect -830 -799 -824 -311
rect -853 -805 -824 -799
rect -724 -311 -695 -305
rect -724 -799 -718 -311
rect -701 -799 -695 -311
rect -724 -805 -695 -799
rect -595 -311 -566 -305
rect -595 -799 -589 -311
rect -572 -799 -566 -311
rect -595 -805 -566 -799
rect -466 -311 -437 -305
rect -466 -799 -460 -311
rect -443 -799 -437 -311
rect -466 -805 -437 -799
rect -337 -311 -308 -305
rect -337 -799 -331 -311
rect -314 -799 -308 -311
rect -337 -805 -308 -799
rect -208 -311 -179 -305
rect -208 -799 -202 -311
rect -185 -799 -179 -311
rect -208 -805 -179 -799
rect -79 -311 -50 -305
rect -79 -799 -73 -311
rect -56 -799 -50 -311
rect -79 -805 -50 -799
rect 50 -311 79 -305
rect 50 -799 56 -311
rect 73 -799 79 -311
rect 50 -805 79 -799
rect 179 -311 208 -305
rect 179 -799 185 -311
rect 202 -799 208 -311
rect 179 -805 208 -799
rect 308 -311 337 -305
rect 308 -799 314 -311
rect 331 -799 337 -311
rect 308 -805 337 -799
rect 437 -311 466 -305
rect 437 -799 443 -311
rect 460 -799 466 -311
rect 437 -805 466 -799
rect 566 -311 595 -305
rect 566 -799 572 -311
rect 589 -799 595 -311
rect 566 -805 595 -799
rect 695 -311 724 -305
rect 695 -799 701 -311
rect 718 -799 724 -311
rect 695 -805 724 -799
rect 824 -311 853 -305
rect 824 -799 830 -311
rect 847 -799 853 -311
rect 824 -805 853 -799
rect 953 -311 982 -305
rect 953 -799 959 -311
rect 976 -799 982 -311
rect 953 -805 982 -799
rect 1082 -311 1111 -305
rect 1082 -799 1088 -311
rect 1105 -799 1111 -311
rect 1082 -805 1111 -799
rect 1211 -311 1240 -305
rect 1211 -799 1217 -311
rect 1234 -799 1240 -311
rect 1211 -805 1240 -799
rect 1340 -311 1369 -305
rect 1340 -799 1346 -311
rect 1363 -799 1369 -311
rect 1340 -805 1369 -799
rect 1469 -311 1498 -305
rect 1469 -799 1475 -311
rect 1492 -799 1498 -311
rect 1469 -805 1498 -799
rect -1498 -866 -1469 -860
rect -1498 -1354 -1492 -866
rect -1475 -1354 -1469 -866
rect -1498 -1360 -1469 -1354
rect -1369 -866 -1340 -860
rect -1369 -1354 -1363 -866
rect -1346 -1354 -1340 -866
rect -1369 -1360 -1340 -1354
rect -1240 -866 -1211 -860
rect -1240 -1354 -1234 -866
rect -1217 -1354 -1211 -866
rect -1240 -1360 -1211 -1354
rect -1111 -866 -1082 -860
rect -1111 -1354 -1105 -866
rect -1088 -1354 -1082 -866
rect -1111 -1360 -1082 -1354
rect -982 -866 -953 -860
rect -982 -1354 -976 -866
rect -959 -1354 -953 -866
rect -982 -1360 -953 -1354
rect -853 -866 -824 -860
rect -853 -1354 -847 -866
rect -830 -1354 -824 -866
rect -853 -1360 -824 -1354
rect -724 -866 -695 -860
rect -724 -1354 -718 -866
rect -701 -1354 -695 -866
rect -724 -1360 -695 -1354
rect -595 -866 -566 -860
rect -595 -1354 -589 -866
rect -572 -1354 -566 -866
rect -595 -1360 -566 -1354
rect -466 -866 -437 -860
rect -466 -1354 -460 -866
rect -443 -1354 -437 -866
rect -466 -1360 -437 -1354
rect -337 -866 -308 -860
rect -337 -1354 -331 -866
rect -314 -1354 -308 -866
rect -337 -1360 -308 -1354
rect -208 -866 -179 -860
rect -208 -1354 -202 -866
rect -185 -1354 -179 -866
rect -208 -1360 -179 -1354
rect -79 -866 -50 -860
rect -79 -1354 -73 -866
rect -56 -1354 -50 -866
rect -79 -1360 -50 -1354
rect 50 -866 79 -860
rect 50 -1354 56 -866
rect 73 -1354 79 -866
rect 50 -1360 79 -1354
rect 179 -866 208 -860
rect 179 -1354 185 -866
rect 202 -1354 208 -866
rect 179 -1360 208 -1354
rect 308 -866 337 -860
rect 308 -1354 314 -866
rect 331 -1354 337 -866
rect 308 -1360 337 -1354
rect 437 -866 466 -860
rect 437 -1354 443 -866
rect 460 -1354 466 -866
rect 437 -1360 466 -1354
rect 566 -866 595 -860
rect 566 -1354 572 -866
rect 589 -1354 595 -866
rect 566 -1360 595 -1354
rect 695 -866 724 -860
rect 695 -1354 701 -866
rect 718 -1354 724 -866
rect 695 -1360 724 -1354
rect 824 -866 853 -860
rect 824 -1354 830 -866
rect 847 -1354 853 -866
rect 824 -1360 853 -1354
rect 953 -866 982 -860
rect 953 -1354 959 -866
rect 976 -1354 982 -866
rect 953 -1360 982 -1354
rect 1082 -866 1111 -860
rect 1082 -1354 1088 -866
rect 1105 -1354 1111 -866
rect 1082 -1360 1111 -1354
rect 1211 -866 1240 -860
rect 1211 -1354 1217 -866
rect 1234 -1354 1240 -866
rect 1211 -1360 1240 -1354
rect 1340 -866 1369 -860
rect 1340 -1354 1346 -866
rect 1363 -1354 1369 -866
rect 1340 -1360 1369 -1354
rect 1469 -866 1498 -860
rect 1469 -1354 1475 -866
rect 1492 -1354 1498 -866
rect 1469 -1360 1498 -1354
<< mvndiffc >>
rect -1492 866 -1475 1354
rect -1363 866 -1346 1354
rect -1234 866 -1217 1354
rect -1105 866 -1088 1354
rect -976 866 -959 1354
rect -847 866 -830 1354
rect -718 866 -701 1354
rect -589 866 -572 1354
rect -460 866 -443 1354
rect -331 866 -314 1354
rect -202 866 -185 1354
rect -73 866 -56 1354
rect 56 866 73 1354
rect 185 866 202 1354
rect 314 866 331 1354
rect 443 866 460 1354
rect 572 866 589 1354
rect 701 866 718 1354
rect 830 866 847 1354
rect 959 866 976 1354
rect 1088 866 1105 1354
rect 1217 866 1234 1354
rect 1346 866 1363 1354
rect 1475 866 1492 1354
rect -1492 311 -1475 799
rect -1363 311 -1346 799
rect -1234 311 -1217 799
rect -1105 311 -1088 799
rect -976 311 -959 799
rect -847 311 -830 799
rect -718 311 -701 799
rect -589 311 -572 799
rect -460 311 -443 799
rect -331 311 -314 799
rect -202 311 -185 799
rect -73 311 -56 799
rect 56 311 73 799
rect 185 311 202 799
rect 314 311 331 799
rect 443 311 460 799
rect 572 311 589 799
rect 701 311 718 799
rect 830 311 847 799
rect 959 311 976 799
rect 1088 311 1105 799
rect 1217 311 1234 799
rect 1346 311 1363 799
rect 1475 311 1492 799
rect -1492 -244 -1475 244
rect -1363 -244 -1346 244
rect -1234 -244 -1217 244
rect -1105 -244 -1088 244
rect -976 -244 -959 244
rect -847 -244 -830 244
rect -718 -244 -701 244
rect -589 -244 -572 244
rect -460 -244 -443 244
rect -331 -244 -314 244
rect -202 -244 -185 244
rect -73 -244 -56 244
rect 56 -244 73 244
rect 185 -244 202 244
rect 314 -244 331 244
rect 443 -244 460 244
rect 572 -244 589 244
rect 701 -244 718 244
rect 830 -244 847 244
rect 959 -244 976 244
rect 1088 -244 1105 244
rect 1217 -244 1234 244
rect 1346 -244 1363 244
rect 1475 -244 1492 244
rect -1492 -799 -1475 -311
rect -1363 -799 -1346 -311
rect -1234 -799 -1217 -311
rect -1105 -799 -1088 -311
rect -976 -799 -959 -311
rect -847 -799 -830 -311
rect -718 -799 -701 -311
rect -589 -799 -572 -311
rect -460 -799 -443 -311
rect -331 -799 -314 -311
rect -202 -799 -185 -311
rect -73 -799 -56 -311
rect 56 -799 73 -311
rect 185 -799 202 -311
rect 314 -799 331 -311
rect 443 -799 460 -311
rect 572 -799 589 -311
rect 701 -799 718 -311
rect 830 -799 847 -311
rect 959 -799 976 -311
rect 1088 -799 1105 -311
rect 1217 -799 1234 -311
rect 1346 -799 1363 -311
rect 1475 -799 1492 -311
rect -1492 -1354 -1475 -866
rect -1363 -1354 -1346 -866
rect -1234 -1354 -1217 -866
rect -1105 -1354 -1088 -866
rect -976 -1354 -959 -866
rect -847 -1354 -830 -866
rect -718 -1354 -701 -866
rect -589 -1354 -572 -866
rect -460 -1354 -443 -866
rect -331 -1354 -314 -866
rect -202 -1354 -185 -866
rect -73 -1354 -56 -866
rect 56 -1354 73 -866
rect 185 -1354 202 -866
rect 314 -1354 331 -866
rect 443 -1354 460 -866
rect 572 -1354 589 -866
rect 701 -1354 718 -866
rect 830 -1354 847 -866
rect 959 -1354 976 -866
rect 1088 -1354 1105 -866
rect 1217 -1354 1234 -866
rect 1346 -1354 1363 -866
rect 1475 -1354 1492 -866
<< mvpsubdiff >>
rect -1565 1465 1565 1471
rect -1565 1448 -1511 1465
rect 1511 1448 1565 1465
rect -1565 1442 1565 1448
rect -1565 1417 -1536 1442
rect -1565 -1417 -1559 1417
rect -1542 -1417 -1536 1417
rect 1536 1417 1565 1442
rect -1565 -1442 -1536 -1417
rect 1536 -1417 1542 1417
rect 1559 -1417 1565 1417
rect 1536 -1442 1565 -1417
rect -1565 -1448 1565 -1442
rect -1565 -1465 -1511 -1448
rect 1511 -1465 1565 -1448
rect -1565 -1471 1565 -1465
<< mvpsubdiffcont >>
rect -1511 1448 1511 1465
rect -1559 -1417 -1542 1417
rect 1542 -1417 1559 1417
rect -1511 -1465 1511 -1448
<< poly >>
rect -1469 1396 -1369 1404
rect -1469 1379 -1461 1396
rect -1377 1379 -1369 1396
rect -1469 1360 -1369 1379
rect -1340 1396 -1240 1404
rect -1340 1379 -1332 1396
rect -1248 1379 -1240 1396
rect -1340 1360 -1240 1379
rect -1211 1396 -1111 1404
rect -1211 1379 -1203 1396
rect -1119 1379 -1111 1396
rect -1211 1360 -1111 1379
rect -1082 1396 -982 1404
rect -1082 1379 -1074 1396
rect -990 1379 -982 1396
rect -1082 1360 -982 1379
rect -953 1396 -853 1404
rect -953 1379 -945 1396
rect -861 1379 -853 1396
rect -953 1360 -853 1379
rect -824 1396 -724 1404
rect -824 1379 -816 1396
rect -732 1379 -724 1396
rect -824 1360 -724 1379
rect -695 1396 -595 1404
rect -695 1379 -687 1396
rect -603 1379 -595 1396
rect -695 1360 -595 1379
rect -566 1396 -466 1404
rect -566 1379 -558 1396
rect -474 1379 -466 1396
rect -566 1360 -466 1379
rect -437 1396 -337 1404
rect -437 1379 -429 1396
rect -345 1379 -337 1396
rect -437 1360 -337 1379
rect -308 1396 -208 1404
rect -308 1379 -300 1396
rect -216 1379 -208 1396
rect -308 1360 -208 1379
rect -179 1396 -79 1404
rect -179 1379 -171 1396
rect -87 1379 -79 1396
rect -179 1360 -79 1379
rect -50 1396 50 1404
rect -50 1379 -42 1396
rect 42 1379 50 1396
rect -50 1360 50 1379
rect 79 1396 179 1404
rect 79 1379 87 1396
rect 171 1379 179 1396
rect 79 1360 179 1379
rect 208 1396 308 1404
rect 208 1379 216 1396
rect 300 1379 308 1396
rect 208 1360 308 1379
rect 337 1396 437 1404
rect 337 1379 345 1396
rect 429 1379 437 1396
rect 337 1360 437 1379
rect 466 1396 566 1404
rect 466 1379 474 1396
rect 558 1379 566 1396
rect 466 1360 566 1379
rect 595 1396 695 1404
rect 595 1379 603 1396
rect 687 1379 695 1396
rect 595 1360 695 1379
rect 724 1396 824 1404
rect 724 1379 732 1396
rect 816 1379 824 1396
rect 724 1360 824 1379
rect 853 1396 953 1404
rect 853 1379 861 1396
rect 945 1379 953 1396
rect 853 1360 953 1379
rect 982 1396 1082 1404
rect 982 1379 990 1396
rect 1074 1379 1082 1396
rect 982 1360 1082 1379
rect 1111 1396 1211 1404
rect 1111 1379 1119 1396
rect 1203 1379 1211 1396
rect 1111 1360 1211 1379
rect 1240 1396 1340 1404
rect 1240 1379 1248 1396
rect 1332 1379 1340 1396
rect 1240 1360 1340 1379
rect 1369 1396 1469 1404
rect 1369 1379 1377 1396
rect 1461 1379 1469 1396
rect 1369 1360 1469 1379
rect -1469 841 -1369 860
rect -1469 824 -1461 841
rect -1377 824 -1369 841
rect -1469 805 -1369 824
rect -1340 841 -1240 860
rect -1340 824 -1332 841
rect -1248 824 -1240 841
rect -1340 805 -1240 824
rect -1211 841 -1111 860
rect -1211 824 -1203 841
rect -1119 824 -1111 841
rect -1211 805 -1111 824
rect -1082 841 -982 860
rect -1082 824 -1074 841
rect -990 824 -982 841
rect -1082 805 -982 824
rect -953 841 -853 860
rect -953 824 -945 841
rect -861 824 -853 841
rect -953 805 -853 824
rect -824 841 -724 860
rect -824 824 -816 841
rect -732 824 -724 841
rect -824 805 -724 824
rect -695 841 -595 860
rect -695 824 -687 841
rect -603 824 -595 841
rect -695 805 -595 824
rect -566 841 -466 860
rect -566 824 -558 841
rect -474 824 -466 841
rect -566 805 -466 824
rect -437 841 -337 860
rect -437 824 -429 841
rect -345 824 -337 841
rect -437 805 -337 824
rect -308 841 -208 860
rect -308 824 -300 841
rect -216 824 -208 841
rect -308 805 -208 824
rect -179 841 -79 860
rect -179 824 -171 841
rect -87 824 -79 841
rect -179 805 -79 824
rect -50 841 50 860
rect -50 824 -42 841
rect 42 824 50 841
rect -50 805 50 824
rect 79 841 179 860
rect 79 824 87 841
rect 171 824 179 841
rect 79 805 179 824
rect 208 841 308 860
rect 208 824 216 841
rect 300 824 308 841
rect 208 805 308 824
rect 337 841 437 860
rect 337 824 345 841
rect 429 824 437 841
rect 337 805 437 824
rect 466 841 566 860
rect 466 824 474 841
rect 558 824 566 841
rect 466 805 566 824
rect 595 841 695 860
rect 595 824 603 841
rect 687 824 695 841
rect 595 805 695 824
rect 724 841 824 860
rect 724 824 732 841
rect 816 824 824 841
rect 724 805 824 824
rect 853 841 953 860
rect 853 824 861 841
rect 945 824 953 841
rect 853 805 953 824
rect 982 841 1082 860
rect 982 824 990 841
rect 1074 824 1082 841
rect 982 805 1082 824
rect 1111 841 1211 860
rect 1111 824 1119 841
rect 1203 824 1211 841
rect 1111 805 1211 824
rect 1240 841 1340 860
rect 1240 824 1248 841
rect 1332 824 1340 841
rect 1240 805 1340 824
rect 1369 841 1469 860
rect 1369 824 1377 841
rect 1461 824 1469 841
rect 1369 805 1469 824
rect -1469 286 -1369 305
rect -1469 269 -1461 286
rect -1377 269 -1369 286
rect -1469 250 -1369 269
rect -1340 286 -1240 305
rect -1340 269 -1332 286
rect -1248 269 -1240 286
rect -1340 250 -1240 269
rect -1211 286 -1111 305
rect -1211 269 -1203 286
rect -1119 269 -1111 286
rect -1211 250 -1111 269
rect -1082 286 -982 305
rect -1082 269 -1074 286
rect -990 269 -982 286
rect -1082 250 -982 269
rect -953 286 -853 305
rect -953 269 -945 286
rect -861 269 -853 286
rect -953 250 -853 269
rect -824 286 -724 305
rect -824 269 -816 286
rect -732 269 -724 286
rect -824 250 -724 269
rect -695 286 -595 305
rect -695 269 -687 286
rect -603 269 -595 286
rect -695 250 -595 269
rect -566 286 -466 305
rect -566 269 -558 286
rect -474 269 -466 286
rect -566 250 -466 269
rect -437 286 -337 305
rect -437 269 -429 286
rect -345 269 -337 286
rect -437 250 -337 269
rect -308 286 -208 305
rect -308 269 -300 286
rect -216 269 -208 286
rect -308 250 -208 269
rect -179 286 -79 305
rect -179 269 -171 286
rect -87 269 -79 286
rect -179 250 -79 269
rect -50 286 50 305
rect -50 269 -42 286
rect 42 269 50 286
rect -50 250 50 269
rect 79 286 179 305
rect 79 269 87 286
rect 171 269 179 286
rect 79 250 179 269
rect 208 286 308 305
rect 208 269 216 286
rect 300 269 308 286
rect 208 250 308 269
rect 337 286 437 305
rect 337 269 345 286
rect 429 269 437 286
rect 337 250 437 269
rect 466 286 566 305
rect 466 269 474 286
rect 558 269 566 286
rect 466 250 566 269
rect 595 286 695 305
rect 595 269 603 286
rect 687 269 695 286
rect 595 250 695 269
rect 724 286 824 305
rect 724 269 732 286
rect 816 269 824 286
rect 724 250 824 269
rect 853 286 953 305
rect 853 269 861 286
rect 945 269 953 286
rect 853 250 953 269
rect 982 286 1082 305
rect 982 269 990 286
rect 1074 269 1082 286
rect 982 250 1082 269
rect 1111 286 1211 305
rect 1111 269 1119 286
rect 1203 269 1211 286
rect 1111 250 1211 269
rect 1240 286 1340 305
rect 1240 269 1248 286
rect 1332 269 1340 286
rect 1240 250 1340 269
rect 1369 286 1469 305
rect 1369 269 1377 286
rect 1461 269 1469 286
rect 1369 250 1469 269
rect -1469 -269 -1369 -250
rect -1469 -286 -1461 -269
rect -1377 -286 -1369 -269
rect -1469 -305 -1369 -286
rect -1340 -269 -1240 -250
rect -1340 -286 -1332 -269
rect -1248 -286 -1240 -269
rect -1340 -305 -1240 -286
rect -1211 -269 -1111 -250
rect -1211 -286 -1203 -269
rect -1119 -286 -1111 -269
rect -1211 -305 -1111 -286
rect -1082 -269 -982 -250
rect -1082 -286 -1074 -269
rect -990 -286 -982 -269
rect -1082 -305 -982 -286
rect -953 -269 -853 -250
rect -953 -286 -945 -269
rect -861 -286 -853 -269
rect -953 -305 -853 -286
rect -824 -269 -724 -250
rect -824 -286 -816 -269
rect -732 -286 -724 -269
rect -824 -305 -724 -286
rect -695 -269 -595 -250
rect -695 -286 -687 -269
rect -603 -286 -595 -269
rect -695 -305 -595 -286
rect -566 -269 -466 -250
rect -566 -286 -558 -269
rect -474 -286 -466 -269
rect -566 -305 -466 -286
rect -437 -269 -337 -250
rect -437 -286 -429 -269
rect -345 -286 -337 -269
rect -437 -305 -337 -286
rect -308 -269 -208 -250
rect -308 -286 -300 -269
rect -216 -286 -208 -269
rect -308 -305 -208 -286
rect -179 -269 -79 -250
rect -179 -286 -171 -269
rect -87 -286 -79 -269
rect -179 -305 -79 -286
rect -50 -269 50 -250
rect -50 -286 -42 -269
rect 42 -286 50 -269
rect -50 -305 50 -286
rect 79 -269 179 -250
rect 79 -286 87 -269
rect 171 -286 179 -269
rect 79 -305 179 -286
rect 208 -269 308 -250
rect 208 -286 216 -269
rect 300 -286 308 -269
rect 208 -305 308 -286
rect 337 -269 437 -250
rect 337 -286 345 -269
rect 429 -286 437 -269
rect 337 -305 437 -286
rect 466 -269 566 -250
rect 466 -286 474 -269
rect 558 -286 566 -269
rect 466 -305 566 -286
rect 595 -269 695 -250
rect 595 -286 603 -269
rect 687 -286 695 -269
rect 595 -305 695 -286
rect 724 -269 824 -250
rect 724 -286 732 -269
rect 816 -286 824 -269
rect 724 -305 824 -286
rect 853 -269 953 -250
rect 853 -286 861 -269
rect 945 -286 953 -269
rect 853 -305 953 -286
rect 982 -269 1082 -250
rect 982 -286 990 -269
rect 1074 -286 1082 -269
rect 982 -305 1082 -286
rect 1111 -269 1211 -250
rect 1111 -286 1119 -269
rect 1203 -286 1211 -269
rect 1111 -305 1211 -286
rect 1240 -269 1340 -250
rect 1240 -286 1248 -269
rect 1332 -286 1340 -269
rect 1240 -305 1340 -286
rect 1369 -269 1469 -250
rect 1369 -286 1377 -269
rect 1461 -286 1469 -269
rect 1369 -305 1469 -286
rect -1469 -824 -1369 -805
rect -1469 -841 -1461 -824
rect -1377 -841 -1369 -824
rect -1469 -860 -1369 -841
rect -1340 -824 -1240 -805
rect -1340 -841 -1332 -824
rect -1248 -841 -1240 -824
rect -1340 -860 -1240 -841
rect -1211 -824 -1111 -805
rect -1211 -841 -1203 -824
rect -1119 -841 -1111 -824
rect -1211 -860 -1111 -841
rect -1082 -824 -982 -805
rect -1082 -841 -1074 -824
rect -990 -841 -982 -824
rect -1082 -860 -982 -841
rect -953 -824 -853 -805
rect -953 -841 -945 -824
rect -861 -841 -853 -824
rect -953 -860 -853 -841
rect -824 -824 -724 -805
rect -824 -841 -816 -824
rect -732 -841 -724 -824
rect -824 -860 -724 -841
rect -695 -824 -595 -805
rect -695 -841 -687 -824
rect -603 -841 -595 -824
rect -695 -860 -595 -841
rect -566 -824 -466 -805
rect -566 -841 -558 -824
rect -474 -841 -466 -824
rect -566 -860 -466 -841
rect -437 -824 -337 -805
rect -437 -841 -429 -824
rect -345 -841 -337 -824
rect -437 -860 -337 -841
rect -308 -824 -208 -805
rect -308 -841 -300 -824
rect -216 -841 -208 -824
rect -308 -860 -208 -841
rect -179 -824 -79 -805
rect -179 -841 -171 -824
rect -87 -841 -79 -824
rect -179 -860 -79 -841
rect -50 -824 50 -805
rect -50 -841 -42 -824
rect 42 -841 50 -824
rect -50 -860 50 -841
rect 79 -824 179 -805
rect 79 -841 87 -824
rect 171 -841 179 -824
rect 79 -860 179 -841
rect 208 -824 308 -805
rect 208 -841 216 -824
rect 300 -841 308 -824
rect 208 -860 308 -841
rect 337 -824 437 -805
rect 337 -841 345 -824
rect 429 -841 437 -824
rect 337 -860 437 -841
rect 466 -824 566 -805
rect 466 -841 474 -824
rect 558 -841 566 -824
rect 466 -860 566 -841
rect 595 -824 695 -805
rect 595 -841 603 -824
rect 687 -841 695 -824
rect 595 -860 695 -841
rect 724 -824 824 -805
rect 724 -841 732 -824
rect 816 -841 824 -824
rect 724 -860 824 -841
rect 853 -824 953 -805
rect 853 -841 861 -824
rect 945 -841 953 -824
rect 853 -860 953 -841
rect 982 -824 1082 -805
rect 982 -841 990 -824
rect 1074 -841 1082 -824
rect 982 -860 1082 -841
rect 1111 -824 1211 -805
rect 1111 -841 1119 -824
rect 1203 -841 1211 -824
rect 1111 -860 1211 -841
rect 1240 -824 1340 -805
rect 1240 -841 1248 -824
rect 1332 -841 1340 -824
rect 1240 -860 1340 -841
rect 1369 -824 1469 -805
rect 1369 -841 1377 -824
rect 1461 -841 1469 -824
rect 1369 -860 1469 -841
rect -1469 -1379 -1369 -1360
rect -1469 -1396 -1461 -1379
rect -1377 -1396 -1369 -1379
rect -1469 -1404 -1369 -1396
rect -1340 -1379 -1240 -1360
rect -1340 -1396 -1332 -1379
rect -1248 -1396 -1240 -1379
rect -1340 -1404 -1240 -1396
rect -1211 -1379 -1111 -1360
rect -1211 -1396 -1203 -1379
rect -1119 -1396 -1111 -1379
rect -1211 -1404 -1111 -1396
rect -1082 -1379 -982 -1360
rect -1082 -1396 -1074 -1379
rect -990 -1396 -982 -1379
rect -1082 -1404 -982 -1396
rect -953 -1379 -853 -1360
rect -953 -1396 -945 -1379
rect -861 -1396 -853 -1379
rect -953 -1404 -853 -1396
rect -824 -1379 -724 -1360
rect -824 -1396 -816 -1379
rect -732 -1396 -724 -1379
rect -824 -1404 -724 -1396
rect -695 -1379 -595 -1360
rect -695 -1396 -687 -1379
rect -603 -1396 -595 -1379
rect -695 -1404 -595 -1396
rect -566 -1379 -466 -1360
rect -566 -1396 -558 -1379
rect -474 -1396 -466 -1379
rect -566 -1404 -466 -1396
rect -437 -1379 -337 -1360
rect -437 -1396 -429 -1379
rect -345 -1396 -337 -1379
rect -437 -1404 -337 -1396
rect -308 -1379 -208 -1360
rect -308 -1396 -300 -1379
rect -216 -1396 -208 -1379
rect -308 -1404 -208 -1396
rect -179 -1379 -79 -1360
rect -179 -1396 -171 -1379
rect -87 -1396 -79 -1379
rect -179 -1404 -79 -1396
rect -50 -1379 50 -1360
rect -50 -1396 -42 -1379
rect 42 -1396 50 -1379
rect -50 -1404 50 -1396
rect 79 -1379 179 -1360
rect 79 -1396 87 -1379
rect 171 -1396 179 -1379
rect 79 -1404 179 -1396
rect 208 -1379 308 -1360
rect 208 -1396 216 -1379
rect 300 -1396 308 -1379
rect 208 -1404 308 -1396
rect 337 -1379 437 -1360
rect 337 -1396 345 -1379
rect 429 -1396 437 -1379
rect 337 -1404 437 -1396
rect 466 -1379 566 -1360
rect 466 -1396 474 -1379
rect 558 -1396 566 -1379
rect 466 -1404 566 -1396
rect 595 -1379 695 -1360
rect 595 -1396 603 -1379
rect 687 -1396 695 -1379
rect 595 -1404 695 -1396
rect 724 -1379 824 -1360
rect 724 -1396 732 -1379
rect 816 -1396 824 -1379
rect 724 -1404 824 -1396
rect 853 -1379 953 -1360
rect 853 -1396 861 -1379
rect 945 -1396 953 -1379
rect 853 -1404 953 -1396
rect 982 -1379 1082 -1360
rect 982 -1396 990 -1379
rect 1074 -1396 1082 -1379
rect 982 -1404 1082 -1396
rect 1111 -1379 1211 -1360
rect 1111 -1396 1119 -1379
rect 1203 -1396 1211 -1379
rect 1111 -1404 1211 -1396
rect 1240 -1379 1340 -1360
rect 1240 -1396 1248 -1379
rect 1332 -1396 1340 -1379
rect 1240 -1404 1340 -1396
rect 1369 -1379 1469 -1360
rect 1369 -1396 1377 -1379
rect 1461 -1396 1469 -1379
rect 1369 -1404 1469 -1396
<< polycont >>
rect -1461 1379 -1377 1396
rect -1332 1379 -1248 1396
rect -1203 1379 -1119 1396
rect -1074 1379 -990 1396
rect -945 1379 -861 1396
rect -816 1379 -732 1396
rect -687 1379 -603 1396
rect -558 1379 -474 1396
rect -429 1379 -345 1396
rect -300 1379 -216 1396
rect -171 1379 -87 1396
rect -42 1379 42 1396
rect 87 1379 171 1396
rect 216 1379 300 1396
rect 345 1379 429 1396
rect 474 1379 558 1396
rect 603 1379 687 1396
rect 732 1379 816 1396
rect 861 1379 945 1396
rect 990 1379 1074 1396
rect 1119 1379 1203 1396
rect 1248 1379 1332 1396
rect 1377 1379 1461 1396
rect -1461 824 -1377 841
rect -1332 824 -1248 841
rect -1203 824 -1119 841
rect -1074 824 -990 841
rect -945 824 -861 841
rect -816 824 -732 841
rect -687 824 -603 841
rect -558 824 -474 841
rect -429 824 -345 841
rect -300 824 -216 841
rect -171 824 -87 841
rect -42 824 42 841
rect 87 824 171 841
rect 216 824 300 841
rect 345 824 429 841
rect 474 824 558 841
rect 603 824 687 841
rect 732 824 816 841
rect 861 824 945 841
rect 990 824 1074 841
rect 1119 824 1203 841
rect 1248 824 1332 841
rect 1377 824 1461 841
rect -1461 269 -1377 286
rect -1332 269 -1248 286
rect -1203 269 -1119 286
rect -1074 269 -990 286
rect -945 269 -861 286
rect -816 269 -732 286
rect -687 269 -603 286
rect -558 269 -474 286
rect -429 269 -345 286
rect -300 269 -216 286
rect -171 269 -87 286
rect -42 269 42 286
rect 87 269 171 286
rect 216 269 300 286
rect 345 269 429 286
rect 474 269 558 286
rect 603 269 687 286
rect 732 269 816 286
rect 861 269 945 286
rect 990 269 1074 286
rect 1119 269 1203 286
rect 1248 269 1332 286
rect 1377 269 1461 286
rect -1461 -286 -1377 -269
rect -1332 -286 -1248 -269
rect -1203 -286 -1119 -269
rect -1074 -286 -990 -269
rect -945 -286 -861 -269
rect -816 -286 -732 -269
rect -687 -286 -603 -269
rect -558 -286 -474 -269
rect -429 -286 -345 -269
rect -300 -286 -216 -269
rect -171 -286 -87 -269
rect -42 -286 42 -269
rect 87 -286 171 -269
rect 216 -286 300 -269
rect 345 -286 429 -269
rect 474 -286 558 -269
rect 603 -286 687 -269
rect 732 -286 816 -269
rect 861 -286 945 -269
rect 990 -286 1074 -269
rect 1119 -286 1203 -269
rect 1248 -286 1332 -269
rect 1377 -286 1461 -269
rect -1461 -841 -1377 -824
rect -1332 -841 -1248 -824
rect -1203 -841 -1119 -824
rect -1074 -841 -990 -824
rect -945 -841 -861 -824
rect -816 -841 -732 -824
rect -687 -841 -603 -824
rect -558 -841 -474 -824
rect -429 -841 -345 -824
rect -300 -841 -216 -824
rect -171 -841 -87 -824
rect -42 -841 42 -824
rect 87 -841 171 -824
rect 216 -841 300 -824
rect 345 -841 429 -824
rect 474 -841 558 -824
rect 603 -841 687 -824
rect 732 -841 816 -824
rect 861 -841 945 -824
rect 990 -841 1074 -824
rect 1119 -841 1203 -824
rect 1248 -841 1332 -824
rect 1377 -841 1461 -824
rect -1461 -1396 -1377 -1379
rect -1332 -1396 -1248 -1379
rect -1203 -1396 -1119 -1379
rect -1074 -1396 -990 -1379
rect -945 -1396 -861 -1379
rect -816 -1396 -732 -1379
rect -687 -1396 -603 -1379
rect -558 -1396 -474 -1379
rect -429 -1396 -345 -1379
rect -300 -1396 -216 -1379
rect -171 -1396 -87 -1379
rect -42 -1396 42 -1379
rect 87 -1396 171 -1379
rect 216 -1396 300 -1379
rect 345 -1396 429 -1379
rect 474 -1396 558 -1379
rect 603 -1396 687 -1379
rect 732 -1396 816 -1379
rect 861 -1396 945 -1379
rect 990 -1396 1074 -1379
rect 1119 -1396 1203 -1379
rect 1248 -1396 1332 -1379
rect 1377 -1396 1461 -1379
<< locali >>
rect -1559 1448 -1511 1465
rect 1511 1448 1559 1465
rect -1559 1417 -1542 1448
rect 1542 1417 1559 1448
rect -1469 1379 -1461 1396
rect -1377 1379 -1369 1396
rect -1340 1379 -1332 1396
rect -1248 1379 -1240 1396
rect -1211 1379 -1203 1396
rect -1119 1379 -1111 1396
rect -1082 1379 -1074 1396
rect -990 1379 -982 1396
rect -953 1379 -945 1396
rect -861 1379 -853 1396
rect -824 1379 -816 1396
rect -732 1379 -724 1396
rect -695 1379 -687 1396
rect -603 1379 -595 1396
rect -566 1379 -558 1396
rect -474 1379 -466 1396
rect -437 1379 -429 1396
rect -345 1379 -337 1396
rect -308 1379 -300 1396
rect -216 1379 -208 1396
rect -179 1379 -171 1396
rect -87 1379 -79 1396
rect -50 1379 -42 1396
rect 42 1379 50 1396
rect 79 1379 87 1396
rect 171 1379 179 1396
rect 208 1379 216 1396
rect 300 1379 308 1396
rect 337 1379 345 1396
rect 429 1379 437 1396
rect 466 1379 474 1396
rect 558 1379 566 1396
rect 595 1379 603 1396
rect 687 1379 695 1396
rect 724 1379 732 1396
rect 816 1379 824 1396
rect 853 1379 861 1396
rect 945 1379 953 1396
rect 982 1379 990 1396
rect 1074 1379 1082 1396
rect 1111 1379 1119 1396
rect 1203 1379 1211 1396
rect 1240 1379 1248 1396
rect 1332 1379 1340 1396
rect 1369 1379 1377 1396
rect 1461 1379 1469 1396
rect -1492 1354 -1475 1362
rect -1492 858 -1475 866
rect -1363 1354 -1346 1362
rect -1363 858 -1346 866
rect -1234 1354 -1217 1362
rect -1234 858 -1217 866
rect -1105 1354 -1088 1362
rect -1105 858 -1088 866
rect -976 1354 -959 1362
rect -976 858 -959 866
rect -847 1354 -830 1362
rect -847 858 -830 866
rect -718 1354 -701 1362
rect -718 858 -701 866
rect -589 1354 -572 1362
rect -589 858 -572 866
rect -460 1354 -443 1362
rect -460 858 -443 866
rect -331 1354 -314 1362
rect -331 858 -314 866
rect -202 1354 -185 1362
rect -202 858 -185 866
rect -73 1354 -56 1362
rect -73 858 -56 866
rect 56 1354 73 1362
rect 56 858 73 866
rect 185 1354 202 1362
rect 185 858 202 866
rect 314 1354 331 1362
rect 314 858 331 866
rect 443 1354 460 1362
rect 443 858 460 866
rect 572 1354 589 1362
rect 572 858 589 866
rect 701 1354 718 1362
rect 701 858 718 866
rect 830 1354 847 1362
rect 830 858 847 866
rect 959 1354 976 1362
rect 959 858 976 866
rect 1088 1354 1105 1362
rect 1088 858 1105 866
rect 1217 1354 1234 1362
rect 1217 858 1234 866
rect 1346 1354 1363 1362
rect 1346 858 1363 866
rect 1475 1354 1492 1362
rect 1475 858 1492 866
rect -1469 824 -1461 841
rect -1377 824 -1369 841
rect -1340 824 -1332 841
rect -1248 824 -1240 841
rect -1211 824 -1203 841
rect -1119 824 -1111 841
rect -1082 824 -1074 841
rect -990 824 -982 841
rect -953 824 -945 841
rect -861 824 -853 841
rect -824 824 -816 841
rect -732 824 -724 841
rect -695 824 -687 841
rect -603 824 -595 841
rect -566 824 -558 841
rect -474 824 -466 841
rect -437 824 -429 841
rect -345 824 -337 841
rect -308 824 -300 841
rect -216 824 -208 841
rect -179 824 -171 841
rect -87 824 -79 841
rect -50 824 -42 841
rect 42 824 50 841
rect 79 824 87 841
rect 171 824 179 841
rect 208 824 216 841
rect 300 824 308 841
rect 337 824 345 841
rect 429 824 437 841
rect 466 824 474 841
rect 558 824 566 841
rect 595 824 603 841
rect 687 824 695 841
rect 724 824 732 841
rect 816 824 824 841
rect 853 824 861 841
rect 945 824 953 841
rect 982 824 990 841
rect 1074 824 1082 841
rect 1111 824 1119 841
rect 1203 824 1211 841
rect 1240 824 1248 841
rect 1332 824 1340 841
rect 1369 824 1377 841
rect 1461 824 1469 841
rect -1492 799 -1475 807
rect -1492 303 -1475 311
rect -1363 799 -1346 807
rect -1363 303 -1346 311
rect -1234 799 -1217 807
rect -1234 303 -1217 311
rect -1105 799 -1088 807
rect -1105 303 -1088 311
rect -976 799 -959 807
rect -976 303 -959 311
rect -847 799 -830 807
rect -847 303 -830 311
rect -718 799 -701 807
rect -718 303 -701 311
rect -589 799 -572 807
rect -589 303 -572 311
rect -460 799 -443 807
rect -460 303 -443 311
rect -331 799 -314 807
rect -331 303 -314 311
rect -202 799 -185 807
rect -202 303 -185 311
rect -73 799 -56 807
rect -73 303 -56 311
rect 56 799 73 807
rect 56 303 73 311
rect 185 799 202 807
rect 185 303 202 311
rect 314 799 331 807
rect 314 303 331 311
rect 443 799 460 807
rect 443 303 460 311
rect 572 799 589 807
rect 572 303 589 311
rect 701 799 718 807
rect 701 303 718 311
rect 830 799 847 807
rect 830 303 847 311
rect 959 799 976 807
rect 959 303 976 311
rect 1088 799 1105 807
rect 1088 303 1105 311
rect 1217 799 1234 807
rect 1217 303 1234 311
rect 1346 799 1363 807
rect 1346 303 1363 311
rect 1475 799 1492 807
rect 1475 303 1492 311
rect -1469 269 -1461 286
rect -1377 269 -1369 286
rect -1340 269 -1332 286
rect -1248 269 -1240 286
rect -1211 269 -1203 286
rect -1119 269 -1111 286
rect -1082 269 -1074 286
rect -990 269 -982 286
rect -953 269 -945 286
rect -861 269 -853 286
rect -824 269 -816 286
rect -732 269 -724 286
rect -695 269 -687 286
rect -603 269 -595 286
rect -566 269 -558 286
rect -474 269 -466 286
rect -437 269 -429 286
rect -345 269 -337 286
rect -308 269 -300 286
rect -216 269 -208 286
rect -179 269 -171 286
rect -87 269 -79 286
rect -50 269 -42 286
rect 42 269 50 286
rect 79 269 87 286
rect 171 269 179 286
rect 208 269 216 286
rect 300 269 308 286
rect 337 269 345 286
rect 429 269 437 286
rect 466 269 474 286
rect 558 269 566 286
rect 595 269 603 286
rect 687 269 695 286
rect 724 269 732 286
rect 816 269 824 286
rect 853 269 861 286
rect 945 269 953 286
rect 982 269 990 286
rect 1074 269 1082 286
rect 1111 269 1119 286
rect 1203 269 1211 286
rect 1240 269 1248 286
rect 1332 269 1340 286
rect 1369 269 1377 286
rect 1461 269 1469 286
rect -1492 244 -1475 252
rect -1492 -252 -1475 -244
rect -1363 244 -1346 252
rect -1363 -252 -1346 -244
rect -1234 244 -1217 252
rect -1234 -252 -1217 -244
rect -1105 244 -1088 252
rect -1105 -252 -1088 -244
rect -976 244 -959 252
rect -976 -252 -959 -244
rect -847 244 -830 252
rect -847 -252 -830 -244
rect -718 244 -701 252
rect -718 -252 -701 -244
rect -589 244 -572 252
rect -589 -252 -572 -244
rect -460 244 -443 252
rect -460 -252 -443 -244
rect -331 244 -314 252
rect -331 -252 -314 -244
rect -202 244 -185 252
rect -202 -252 -185 -244
rect -73 244 -56 252
rect -73 -252 -56 -244
rect 56 244 73 252
rect 56 -252 73 -244
rect 185 244 202 252
rect 185 -252 202 -244
rect 314 244 331 252
rect 314 -252 331 -244
rect 443 244 460 252
rect 443 -252 460 -244
rect 572 244 589 252
rect 572 -252 589 -244
rect 701 244 718 252
rect 701 -252 718 -244
rect 830 244 847 252
rect 830 -252 847 -244
rect 959 244 976 252
rect 959 -252 976 -244
rect 1088 244 1105 252
rect 1088 -252 1105 -244
rect 1217 244 1234 252
rect 1217 -252 1234 -244
rect 1346 244 1363 252
rect 1346 -252 1363 -244
rect 1475 244 1492 252
rect 1475 -252 1492 -244
rect -1469 -286 -1461 -269
rect -1377 -286 -1369 -269
rect -1340 -286 -1332 -269
rect -1248 -286 -1240 -269
rect -1211 -286 -1203 -269
rect -1119 -286 -1111 -269
rect -1082 -286 -1074 -269
rect -990 -286 -982 -269
rect -953 -286 -945 -269
rect -861 -286 -853 -269
rect -824 -286 -816 -269
rect -732 -286 -724 -269
rect -695 -286 -687 -269
rect -603 -286 -595 -269
rect -566 -286 -558 -269
rect -474 -286 -466 -269
rect -437 -286 -429 -269
rect -345 -286 -337 -269
rect -308 -286 -300 -269
rect -216 -286 -208 -269
rect -179 -286 -171 -269
rect -87 -286 -79 -269
rect -50 -286 -42 -269
rect 42 -286 50 -269
rect 79 -286 87 -269
rect 171 -286 179 -269
rect 208 -286 216 -269
rect 300 -286 308 -269
rect 337 -286 345 -269
rect 429 -286 437 -269
rect 466 -286 474 -269
rect 558 -286 566 -269
rect 595 -286 603 -269
rect 687 -286 695 -269
rect 724 -286 732 -269
rect 816 -286 824 -269
rect 853 -286 861 -269
rect 945 -286 953 -269
rect 982 -286 990 -269
rect 1074 -286 1082 -269
rect 1111 -286 1119 -269
rect 1203 -286 1211 -269
rect 1240 -286 1248 -269
rect 1332 -286 1340 -269
rect 1369 -286 1377 -269
rect 1461 -286 1469 -269
rect -1492 -311 -1475 -303
rect -1492 -807 -1475 -799
rect -1363 -311 -1346 -303
rect -1363 -807 -1346 -799
rect -1234 -311 -1217 -303
rect -1234 -807 -1217 -799
rect -1105 -311 -1088 -303
rect -1105 -807 -1088 -799
rect -976 -311 -959 -303
rect -976 -807 -959 -799
rect -847 -311 -830 -303
rect -847 -807 -830 -799
rect -718 -311 -701 -303
rect -718 -807 -701 -799
rect -589 -311 -572 -303
rect -589 -807 -572 -799
rect -460 -311 -443 -303
rect -460 -807 -443 -799
rect -331 -311 -314 -303
rect -331 -807 -314 -799
rect -202 -311 -185 -303
rect -202 -807 -185 -799
rect -73 -311 -56 -303
rect -73 -807 -56 -799
rect 56 -311 73 -303
rect 56 -807 73 -799
rect 185 -311 202 -303
rect 185 -807 202 -799
rect 314 -311 331 -303
rect 314 -807 331 -799
rect 443 -311 460 -303
rect 443 -807 460 -799
rect 572 -311 589 -303
rect 572 -807 589 -799
rect 701 -311 718 -303
rect 701 -807 718 -799
rect 830 -311 847 -303
rect 830 -807 847 -799
rect 959 -311 976 -303
rect 959 -807 976 -799
rect 1088 -311 1105 -303
rect 1088 -807 1105 -799
rect 1217 -311 1234 -303
rect 1217 -807 1234 -799
rect 1346 -311 1363 -303
rect 1346 -807 1363 -799
rect 1475 -311 1492 -303
rect 1475 -807 1492 -799
rect -1469 -841 -1461 -824
rect -1377 -841 -1369 -824
rect -1340 -841 -1332 -824
rect -1248 -841 -1240 -824
rect -1211 -841 -1203 -824
rect -1119 -841 -1111 -824
rect -1082 -841 -1074 -824
rect -990 -841 -982 -824
rect -953 -841 -945 -824
rect -861 -841 -853 -824
rect -824 -841 -816 -824
rect -732 -841 -724 -824
rect -695 -841 -687 -824
rect -603 -841 -595 -824
rect -566 -841 -558 -824
rect -474 -841 -466 -824
rect -437 -841 -429 -824
rect -345 -841 -337 -824
rect -308 -841 -300 -824
rect -216 -841 -208 -824
rect -179 -841 -171 -824
rect -87 -841 -79 -824
rect -50 -841 -42 -824
rect 42 -841 50 -824
rect 79 -841 87 -824
rect 171 -841 179 -824
rect 208 -841 216 -824
rect 300 -841 308 -824
rect 337 -841 345 -824
rect 429 -841 437 -824
rect 466 -841 474 -824
rect 558 -841 566 -824
rect 595 -841 603 -824
rect 687 -841 695 -824
rect 724 -841 732 -824
rect 816 -841 824 -824
rect 853 -841 861 -824
rect 945 -841 953 -824
rect 982 -841 990 -824
rect 1074 -841 1082 -824
rect 1111 -841 1119 -824
rect 1203 -841 1211 -824
rect 1240 -841 1248 -824
rect 1332 -841 1340 -824
rect 1369 -841 1377 -824
rect 1461 -841 1469 -824
rect -1492 -866 -1475 -858
rect -1492 -1362 -1475 -1354
rect -1363 -866 -1346 -858
rect -1363 -1362 -1346 -1354
rect -1234 -866 -1217 -858
rect -1234 -1362 -1217 -1354
rect -1105 -866 -1088 -858
rect -1105 -1362 -1088 -1354
rect -976 -866 -959 -858
rect -976 -1362 -959 -1354
rect -847 -866 -830 -858
rect -847 -1362 -830 -1354
rect -718 -866 -701 -858
rect -718 -1362 -701 -1354
rect -589 -866 -572 -858
rect -589 -1362 -572 -1354
rect -460 -866 -443 -858
rect -460 -1362 -443 -1354
rect -331 -866 -314 -858
rect -331 -1362 -314 -1354
rect -202 -866 -185 -858
rect -202 -1362 -185 -1354
rect -73 -866 -56 -858
rect -73 -1362 -56 -1354
rect 56 -866 73 -858
rect 56 -1362 73 -1354
rect 185 -866 202 -858
rect 185 -1362 202 -1354
rect 314 -866 331 -858
rect 314 -1362 331 -1354
rect 443 -866 460 -858
rect 443 -1362 460 -1354
rect 572 -866 589 -858
rect 572 -1362 589 -1354
rect 701 -866 718 -858
rect 701 -1362 718 -1354
rect 830 -866 847 -858
rect 830 -1362 847 -1354
rect 959 -866 976 -858
rect 959 -1362 976 -1354
rect 1088 -866 1105 -858
rect 1088 -1362 1105 -1354
rect 1217 -866 1234 -858
rect 1217 -1362 1234 -1354
rect 1346 -866 1363 -858
rect 1346 -1362 1363 -1354
rect 1475 -866 1492 -858
rect 1475 -1362 1492 -1354
rect -1469 -1396 -1461 -1379
rect -1377 -1396 -1369 -1379
rect -1340 -1396 -1332 -1379
rect -1248 -1396 -1240 -1379
rect -1211 -1396 -1203 -1379
rect -1119 -1396 -1111 -1379
rect -1082 -1396 -1074 -1379
rect -990 -1396 -982 -1379
rect -953 -1396 -945 -1379
rect -861 -1396 -853 -1379
rect -824 -1396 -816 -1379
rect -732 -1396 -724 -1379
rect -695 -1396 -687 -1379
rect -603 -1396 -595 -1379
rect -566 -1396 -558 -1379
rect -474 -1396 -466 -1379
rect -437 -1396 -429 -1379
rect -345 -1396 -337 -1379
rect -308 -1396 -300 -1379
rect -216 -1396 -208 -1379
rect -179 -1396 -171 -1379
rect -87 -1396 -79 -1379
rect -50 -1396 -42 -1379
rect 42 -1396 50 -1379
rect 79 -1396 87 -1379
rect 171 -1396 179 -1379
rect 208 -1396 216 -1379
rect 300 -1396 308 -1379
rect 337 -1396 345 -1379
rect 429 -1396 437 -1379
rect 466 -1396 474 -1379
rect 558 -1396 566 -1379
rect 595 -1396 603 -1379
rect 687 -1396 695 -1379
rect 724 -1396 732 -1379
rect 816 -1396 824 -1379
rect 853 -1396 861 -1379
rect 945 -1396 953 -1379
rect 982 -1396 990 -1379
rect 1074 -1396 1082 -1379
rect 1111 -1396 1119 -1379
rect 1203 -1396 1211 -1379
rect 1240 -1396 1248 -1379
rect 1332 -1396 1340 -1379
rect 1369 -1396 1377 -1379
rect 1461 -1396 1469 -1379
rect -1559 -1448 -1542 -1417
rect 1542 -1448 1559 -1417
rect -1559 -1465 -1511 -1448
rect 1511 -1465 1559 -1448
<< viali >>
rect -1461 1379 -1377 1396
rect -1332 1379 -1248 1396
rect -1203 1379 -1119 1396
rect -1074 1379 -990 1396
rect -945 1379 -861 1396
rect -816 1379 -732 1396
rect -687 1379 -603 1396
rect -558 1379 -474 1396
rect -429 1379 -345 1396
rect -300 1379 -216 1396
rect -171 1379 -87 1396
rect -42 1379 42 1396
rect 87 1379 171 1396
rect 216 1379 300 1396
rect 345 1379 429 1396
rect 474 1379 558 1396
rect 603 1379 687 1396
rect 732 1379 816 1396
rect 861 1379 945 1396
rect 990 1379 1074 1396
rect 1119 1379 1203 1396
rect 1248 1379 1332 1396
rect 1377 1379 1461 1396
rect -1492 866 -1475 1354
rect -1363 866 -1346 1354
rect -1234 866 -1217 1354
rect -1105 866 -1088 1354
rect -976 866 -959 1354
rect -847 866 -830 1354
rect -718 866 -701 1354
rect -589 866 -572 1354
rect -460 866 -443 1354
rect -331 866 -314 1354
rect -202 866 -185 1354
rect -73 866 -56 1354
rect 56 866 73 1354
rect 185 866 202 1354
rect 314 866 331 1354
rect 443 866 460 1354
rect 572 866 589 1354
rect 701 866 718 1354
rect 830 866 847 1354
rect 959 866 976 1354
rect 1088 866 1105 1354
rect 1217 866 1234 1354
rect 1346 866 1363 1354
rect 1475 866 1492 1354
rect -1461 824 -1377 841
rect -1332 824 -1248 841
rect -1203 824 -1119 841
rect -1074 824 -990 841
rect -945 824 -861 841
rect -816 824 -732 841
rect -687 824 -603 841
rect -558 824 -474 841
rect -429 824 -345 841
rect -300 824 -216 841
rect -171 824 -87 841
rect -42 824 42 841
rect 87 824 171 841
rect 216 824 300 841
rect 345 824 429 841
rect 474 824 558 841
rect 603 824 687 841
rect 732 824 816 841
rect 861 824 945 841
rect 990 824 1074 841
rect 1119 824 1203 841
rect 1248 824 1332 841
rect 1377 824 1461 841
rect -1492 311 -1475 799
rect -1363 311 -1346 799
rect -1234 311 -1217 799
rect -1105 311 -1088 799
rect -976 311 -959 799
rect -847 311 -830 799
rect -718 311 -701 799
rect -589 311 -572 799
rect -460 311 -443 799
rect -331 311 -314 799
rect -202 311 -185 799
rect -73 311 -56 799
rect 56 311 73 799
rect 185 311 202 799
rect 314 311 331 799
rect 443 311 460 799
rect 572 311 589 799
rect 701 311 718 799
rect 830 311 847 799
rect 959 311 976 799
rect 1088 311 1105 799
rect 1217 311 1234 799
rect 1346 311 1363 799
rect 1475 311 1492 799
rect -1461 269 -1377 286
rect -1332 269 -1248 286
rect -1203 269 -1119 286
rect -1074 269 -990 286
rect -945 269 -861 286
rect -816 269 -732 286
rect -687 269 -603 286
rect -558 269 -474 286
rect -429 269 -345 286
rect -300 269 -216 286
rect -171 269 -87 286
rect -42 269 42 286
rect 87 269 171 286
rect 216 269 300 286
rect 345 269 429 286
rect 474 269 558 286
rect 603 269 687 286
rect 732 269 816 286
rect 861 269 945 286
rect 990 269 1074 286
rect 1119 269 1203 286
rect 1248 269 1332 286
rect 1377 269 1461 286
rect -1492 -244 -1475 244
rect -1363 -244 -1346 244
rect -1234 -244 -1217 244
rect -1105 -244 -1088 244
rect -976 -244 -959 244
rect -847 -244 -830 244
rect -718 -244 -701 244
rect -589 -244 -572 244
rect -460 -244 -443 244
rect -331 -244 -314 244
rect -202 -244 -185 244
rect -73 -244 -56 244
rect 56 -244 73 244
rect 185 -244 202 244
rect 314 -244 331 244
rect 443 -244 460 244
rect 572 -244 589 244
rect 701 -244 718 244
rect 830 -244 847 244
rect 959 -244 976 244
rect 1088 -244 1105 244
rect 1217 -244 1234 244
rect 1346 -244 1363 244
rect 1475 -244 1492 244
rect -1461 -286 -1377 -269
rect -1332 -286 -1248 -269
rect -1203 -286 -1119 -269
rect -1074 -286 -990 -269
rect -945 -286 -861 -269
rect -816 -286 -732 -269
rect -687 -286 -603 -269
rect -558 -286 -474 -269
rect -429 -286 -345 -269
rect -300 -286 -216 -269
rect -171 -286 -87 -269
rect -42 -286 42 -269
rect 87 -286 171 -269
rect 216 -286 300 -269
rect 345 -286 429 -269
rect 474 -286 558 -269
rect 603 -286 687 -269
rect 732 -286 816 -269
rect 861 -286 945 -269
rect 990 -286 1074 -269
rect 1119 -286 1203 -269
rect 1248 -286 1332 -269
rect 1377 -286 1461 -269
rect -1492 -799 -1475 -311
rect -1363 -799 -1346 -311
rect -1234 -799 -1217 -311
rect -1105 -799 -1088 -311
rect -976 -799 -959 -311
rect -847 -799 -830 -311
rect -718 -799 -701 -311
rect -589 -799 -572 -311
rect -460 -799 -443 -311
rect -331 -799 -314 -311
rect -202 -799 -185 -311
rect -73 -799 -56 -311
rect 56 -799 73 -311
rect 185 -799 202 -311
rect 314 -799 331 -311
rect 443 -799 460 -311
rect 572 -799 589 -311
rect 701 -799 718 -311
rect 830 -799 847 -311
rect 959 -799 976 -311
rect 1088 -799 1105 -311
rect 1217 -799 1234 -311
rect 1346 -799 1363 -311
rect 1475 -799 1492 -311
rect -1461 -841 -1377 -824
rect -1332 -841 -1248 -824
rect -1203 -841 -1119 -824
rect -1074 -841 -990 -824
rect -945 -841 -861 -824
rect -816 -841 -732 -824
rect -687 -841 -603 -824
rect -558 -841 -474 -824
rect -429 -841 -345 -824
rect -300 -841 -216 -824
rect -171 -841 -87 -824
rect -42 -841 42 -824
rect 87 -841 171 -824
rect 216 -841 300 -824
rect 345 -841 429 -824
rect 474 -841 558 -824
rect 603 -841 687 -824
rect 732 -841 816 -824
rect 861 -841 945 -824
rect 990 -841 1074 -824
rect 1119 -841 1203 -824
rect 1248 -841 1332 -824
rect 1377 -841 1461 -824
rect -1492 -1354 -1475 -866
rect -1363 -1354 -1346 -866
rect -1234 -1354 -1217 -866
rect -1105 -1354 -1088 -866
rect -976 -1354 -959 -866
rect -847 -1354 -830 -866
rect -718 -1354 -701 -866
rect -589 -1354 -572 -866
rect -460 -1354 -443 -866
rect -331 -1354 -314 -866
rect -202 -1354 -185 -866
rect -73 -1354 -56 -866
rect 56 -1354 73 -866
rect 185 -1354 202 -866
rect 314 -1354 331 -866
rect 443 -1354 460 -866
rect 572 -1354 589 -866
rect 701 -1354 718 -866
rect 830 -1354 847 -866
rect 959 -1354 976 -866
rect 1088 -1354 1105 -866
rect 1217 -1354 1234 -866
rect 1346 -1354 1363 -866
rect 1475 -1354 1492 -866
rect -1461 -1396 -1377 -1379
rect -1332 -1396 -1248 -1379
rect -1203 -1396 -1119 -1379
rect -1074 -1396 -990 -1379
rect -945 -1396 -861 -1379
rect -816 -1396 -732 -1379
rect -687 -1396 -603 -1379
rect -558 -1396 -474 -1379
rect -429 -1396 -345 -1379
rect -300 -1396 -216 -1379
rect -171 -1396 -87 -1379
rect -42 -1396 42 -1379
rect 87 -1396 171 -1379
rect 216 -1396 300 -1379
rect 345 -1396 429 -1379
rect 474 -1396 558 -1379
rect 603 -1396 687 -1379
rect 732 -1396 816 -1379
rect 861 -1396 945 -1379
rect 990 -1396 1074 -1379
rect 1119 -1396 1203 -1379
rect 1248 -1396 1332 -1379
rect 1377 -1396 1461 -1379
<< metal1 >>
rect -1467 1396 -1371 1399
rect -1467 1379 -1461 1396
rect -1377 1379 -1371 1396
rect -1467 1376 -1371 1379
rect -1338 1396 -1242 1399
rect -1338 1379 -1332 1396
rect -1248 1379 -1242 1396
rect -1338 1376 -1242 1379
rect -1209 1396 -1113 1399
rect -1209 1379 -1203 1396
rect -1119 1379 -1113 1396
rect -1209 1376 -1113 1379
rect -1080 1396 -984 1399
rect -1080 1379 -1074 1396
rect -990 1379 -984 1396
rect -1080 1376 -984 1379
rect -951 1396 -855 1399
rect -951 1379 -945 1396
rect -861 1379 -855 1396
rect -951 1376 -855 1379
rect -822 1396 -726 1399
rect -822 1379 -816 1396
rect -732 1379 -726 1396
rect -822 1376 -726 1379
rect -693 1396 -597 1399
rect -693 1379 -687 1396
rect -603 1379 -597 1396
rect -693 1376 -597 1379
rect -564 1396 -468 1399
rect -564 1379 -558 1396
rect -474 1379 -468 1396
rect -564 1376 -468 1379
rect -435 1396 -339 1399
rect -435 1379 -429 1396
rect -345 1379 -339 1396
rect -435 1376 -339 1379
rect -306 1396 -210 1399
rect -306 1379 -300 1396
rect -216 1379 -210 1396
rect -306 1376 -210 1379
rect -177 1396 -81 1399
rect -177 1379 -171 1396
rect -87 1379 -81 1396
rect -177 1376 -81 1379
rect -48 1396 48 1399
rect -48 1379 -42 1396
rect 42 1379 48 1396
rect -48 1376 48 1379
rect 81 1396 177 1399
rect 81 1379 87 1396
rect 171 1379 177 1396
rect 81 1376 177 1379
rect 210 1396 306 1399
rect 210 1379 216 1396
rect 300 1379 306 1396
rect 210 1376 306 1379
rect 339 1396 435 1399
rect 339 1379 345 1396
rect 429 1379 435 1396
rect 339 1376 435 1379
rect 468 1396 564 1399
rect 468 1379 474 1396
rect 558 1379 564 1396
rect 468 1376 564 1379
rect 597 1396 693 1399
rect 597 1379 603 1396
rect 687 1379 693 1396
rect 597 1376 693 1379
rect 726 1396 822 1399
rect 726 1379 732 1396
rect 816 1379 822 1396
rect 726 1376 822 1379
rect 855 1396 951 1399
rect 855 1379 861 1396
rect 945 1379 951 1396
rect 855 1376 951 1379
rect 984 1396 1080 1399
rect 984 1379 990 1396
rect 1074 1379 1080 1396
rect 984 1376 1080 1379
rect 1113 1396 1209 1399
rect 1113 1379 1119 1396
rect 1203 1379 1209 1396
rect 1113 1376 1209 1379
rect 1242 1396 1338 1399
rect 1242 1379 1248 1396
rect 1332 1379 1338 1396
rect 1242 1376 1338 1379
rect 1371 1396 1467 1399
rect 1371 1379 1377 1396
rect 1461 1379 1467 1396
rect 1371 1376 1467 1379
rect -1495 1354 -1472 1360
rect -1495 866 -1492 1354
rect -1475 866 -1472 1354
rect -1495 860 -1472 866
rect -1366 1354 -1343 1360
rect -1366 866 -1363 1354
rect -1346 866 -1343 1354
rect -1366 860 -1343 866
rect -1237 1354 -1214 1360
rect -1237 866 -1234 1354
rect -1217 866 -1214 1354
rect -1237 860 -1214 866
rect -1108 1354 -1085 1360
rect -1108 866 -1105 1354
rect -1088 866 -1085 1354
rect -1108 860 -1085 866
rect -979 1354 -956 1360
rect -979 866 -976 1354
rect -959 866 -956 1354
rect -979 860 -956 866
rect -850 1354 -827 1360
rect -850 866 -847 1354
rect -830 866 -827 1354
rect -850 860 -827 866
rect -721 1354 -698 1360
rect -721 866 -718 1354
rect -701 866 -698 1354
rect -721 860 -698 866
rect -592 1354 -569 1360
rect -592 866 -589 1354
rect -572 866 -569 1354
rect -592 860 -569 866
rect -463 1354 -440 1360
rect -463 866 -460 1354
rect -443 866 -440 1354
rect -463 860 -440 866
rect -334 1354 -311 1360
rect -334 866 -331 1354
rect -314 866 -311 1354
rect -334 860 -311 866
rect -205 1354 -182 1360
rect -205 866 -202 1354
rect -185 866 -182 1354
rect -205 860 -182 866
rect -76 1354 -53 1360
rect -76 866 -73 1354
rect -56 866 -53 1354
rect -76 860 -53 866
rect 53 1354 76 1360
rect 53 866 56 1354
rect 73 866 76 1354
rect 53 860 76 866
rect 182 1354 205 1360
rect 182 866 185 1354
rect 202 866 205 1354
rect 182 860 205 866
rect 311 1354 334 1360
rect 311 866 314 1354
rect 331 866 334 1354
rect 311 860 334 866
rect 440 1354 463 1360
rect 440 866 443 1354
rect 460 866 463 1354
rect 440 860 463 866
rect 569 1354 592 1360
rect 569 866 572 1354
rect 589 866 592 1354
rect 569 860 592 866
rect 698 1354 721 1360
rect 698 866 701 1354
rect 718 866 721 1354
rect 698 860 721 866
rect 827 1354 850 1360
rect 827 866 830 1354
rect 847 866 850 1354
rect 827 860 850 866
rect 956 1354 979 1360
rect 956 866 959 1354
rect 976 866 979 1354
rect 956 860 979 866
rect 1085 1354 1108 1360
rect 1085 866 1088 1354
rect 1105 866 1108 1354
rect 1085 860 1108 866
rect 1214 1354 1237 1360
rect 1214 866 1217 1354
rect 1234 866 1237 1354
rect 1214 860 1237 866
rect 1343 1354 1366 1360
rect 1343 866 1346 1354
rect 1363 866 1366 1354
rect 1343 860 1366 866
rect 1472 1354 1495 1360
rect 1472 866 1475 1354
rect 1492 866 1495 1354
rect 1472 860 1495 866
rect -1467 841 -1371 844
rect -1467 824 -1461 841
rect -1377 824 -1371 841
rect -1467 821 -1371 824
rect -1338 841 -1242 844
rect -1338 824 -1332 841
rect -1248 824 -1242 841
rect -1338 821 -1242 824
rect -1209 841 -1113 844
rect -1209 824 -1203 841
rect -1119 824 -1113 841
rect -1209 821 -1113 824
rect -1080 841 -984 844
rect -1080 824 -1074 841
rect -990 824 -984 841
rect -1080 821 -984 824
rect -951 841 -855 844
rect -951 824 -945 841
rect -861 824 -855 841
rect -951 821 -855 824
rect -822 841 -726 844
rect -822 824 -816 841
rect -732 824 -726 841
rect -822 821 -726 824
rect -693 841 -597 844
rect -693 824 -687 841
rect -603 824 -597 841
rect -693 821 -597 824
rect -564 841 -468 844
rect -564 824 -558 841
rect -474 824 -468 841
rect -564 821 -468 824
rect -435 841 -339 844
rect -435 824 -429 841
rect -345 824 -339 841
rect -435 821 -339 824
rect -306 841 -210 844
rect -306 824 -300 841
rect -216 824 -210 841
rect -306 821 -210 824
rect -177 841 -81 844
rect -177 824 -171 841
rect -87 824 -81 841
rect -177 821 -81 824
rect -48 841 48 844
rect -48 824 -42 841
rect 42 824 48 841
rect -48 821 48 824
rect 81 841 177 844
rect 81 824 87 841
rect 171 824 177 841
rect 81 821 177 824
rect 210 841 306 844
rect 210 824 216 841
rect 300 824 306 841
rect 210 821 306 824
rect 339 841 435 844
rect 339 824 345 841
rect 429 824 435 841
rect 339 821 435 824
rect 468 841 564 844
rect 468 824 474 841
rect 558 824 564 841
rect 468 821 564 824
rect 597 841 693 844
rect 597 824 603 841
rect 687 824 693 841
rect 597 821 693 824
rect 726 841 822 844
rect 726 824 732 841
rect 816 824 822 841
rect 726 821 822 824
rect 855 841 951 844
rect 855 824 861 841
rect 945 824 951 841
rect 855 821 951 824
rect 984 841 1080 844
rect 984 824 990 841
rect 1074 824 1080 841
rect 984 821 1080 824
rect 1113 841 1209 844
rect 1113 824 1119 841
rect 1203 824 1209 841
rect 1113 821 1209 824
rect 1242 841 1338 844
rect 1242 824 1248 841
rect 1332 824 1338 841
rect 1242 821 1338 824
rect 1371 841 1467 844
rect 1371 824 1377 841
rect 1461 824 1467 841
rect 1371 821 1467 824
rect -1495 799 -1472 805
rect -1495 311 -1492 799
rect -1475 311 -1472 799
rect -1495 305 -1472 311
rect -1366 799 -1343 805
rect -1366 311 -1363 799
rect -1346 311 -1343 799
rect -1366 305 -1343 311
rect -1237 799 -1214 805
rect -1237 311 -1234 799
rect -1217 311 -1214 799
rect -1237 305 -1214 311
rect -1108 799 -1085 805
rect -1108 311 -1105 799
rect -1088 311 -1085 799
rect -1108 305 -1085 311
rect -979 799 -956 805
rect -979 311 -976 799
rect -959 311 -956 799
rect -979 305 -956 311
rect -850 799 -827 805
rect -850 311 -847 799
rect -830 311 -827 799
rect -850 305 -827 311
rect -721 799 -698 805
rect -721 311 -718 799
rect -701 311 -698 799
rect -721 305 -698 311
rect -592 799 -569 805
rect -592 311 -589 799
rect -572 311 -569 799
rect -592 305 -569 311
rect -463 799 -440 805
rect -463 311 -460 799
rect -443 311 -440 799
rect -463 305 -440 311
rect -334 799 -311 805
rect -334 311 -331 799
rect -314 311 -311 799
rect -334 305 -311 311
rect -205 799 -182 805
rect -205 311 -202 799
rect -185 311 -182 799
rect -205 305 -182 311
rect -76 799 -53 805
rect -76 311 -73 799
rect -56 311 -53 799
rect -76 305 -53 311
rect 53 799 76 805
rect 53 311 56 799
rect 73 311 76 799
rect 53 305 76 311
rect 182 799 205 805
rect 182 311 185 799
rect 202 311 205 799
rect 182 305 205 311
rect 311 799 334 805
rect 311 311 314 799
rect 331 311 334 799
rect 311 305 334 311
rect 440 799 463 805
rect 440 311 443 799
rect 460 311 463 799
rect 440 305 463 311
rect 569 799 592 805
rect 569 311 572 799
rect 589 311 592 799
rect 569 305 592 311
rect 698 799 721 805
rect 698 311 701 799
rect 718 311 721 799
rect 698 305 721 311
rect 827 799 850 805
rect 827 311 830 799
rect 847 311 850 799
rect 827 305 850 311
rect 956 799 979 805
rect 956 311 959 799
rect 976 311 979 799
rect 956 305 979 311
rect 1085 799 1108 805
rect 1085 311 1088 799
rect 1105 311 1108 799
rect 1085 305 1108 311
rect 1214 799 1237 805
rect 1214 311 1217 799
rect 1234 311 1237 799
rect 1214 305 1237 311
rect 1343 799 1366 805
rect 1343 311 1346 799
rect 1363 311 1366 799
rect 1343 305 1366 311
rect 1472 799 1495 805
rect 1472 311 1475 799
rect 1492 311 1495 799
rect 1472 305 1495 311
rect -1467 286 -1371 289
rect -1467 269 -1461 286
rect -1377 269 -1371 286
rect -1467 266 -1371 269
rect -1338 286 -1242 289
rect -1338 269 -1332 286
rect -1248 269 -1242 286
rect -1338 266 -1242 269
rect -1209 286 -1113 289
rect -1209 269 -1203 286
rect -1119 269 -1113 286
rect -1209 266 -1113 269
rect -1080 286 -984 289
rect -1080 269 -1074 286
rect -990 269 -984 286
rect -1080 266 -984 269
rect -951 286 -855 289
rect -951 269 -945 286
rect -861 269 -855 286
rect -951 266 -855 269
rect -822 286 -726 289
rect -822 269 -816 286
rect -732 269 -726 286
rect -822 266 -726 269
rect -693 286 -597 289
rect -693 269 -687 286
rect -603 269 -597 286
rect -693 266 -597 269
rect -564 286 -468 289
rect -564 269 -558 286
rect -474 269 -468 286
rect -564 266 -468 269
rect -435 286 -339 289
rect -435 269 -429 286
rect -345 269 -339 286
rect -435 266 -339 269
rect -306 286 -210 289
rect -306 269 -300 286
rect -216 269 -210 286
rect -306 266 -210 269
rect -177 286 -81 289
rect -177 269 -171 286
rect -87 269 -81 286
rect -177 266 -81 269
rect -48 286 48 289
rect -48 269 -42 286
rect 42 269 48 286
rect -48 266 48 269
rect 81 286 177 289
rect 81 269 87 286
rect 171 269 177 286
rect 81 266 177 269
rect 210 286 306 289
rect 210 269 216 286
rect 300 269 306 286
rect 210 266 306 269
rect 339 286 435 289
rect 339 269 345 286
rect 429 269 435 286
rect 339 266 435 269
rect 468 286 564 289
rect 468 269 474 286
rect 558 269 564 286
rect 468 266 564 269
rect 597 286 693 289
rect 597 269 603 286
rect 687 269 693 286
rect 597 266 693 269
rect 726 286 822 289
rect 726 269 732 286
rect 816 269 822 286
rect 726 266 822 269
rect 855 286 951 289
rect 855 269 861 286
rect 945 269 951 286
rect 855 266 951 269
rect 984 286 1080 289
rect 984 269 990 286
rect 1074 269 1080 286
rect 984 266 1080 269
rect 1113 286 1209 289
rect 1113 269 1119 286
rect 1203 269 1209 286
rect 1113 266 1209 269
rect 1242 286 1338 289
rect 1242 269 1248 286
rect 1332 269 1338 286
rect 1242 266 1338 269
rect 1371 286 1467 289
rect 1371 269 1377 286
rect 1461 269 1467 286
rect 1371 266 1467 269
rect -1495 244 -1472 250
rect -1495 -244 -1492 244
rect -1475 -244 -1472 244
rect -1495 -250 -1472 -244
rect -1366 244 -1343 250
rect -1366 -244 -1363 244
rect -1346 -244 -1343 244
rect -1366 -250 -1343 -244
rect -1237 244 -1214 250
rect -1237 -244 -1234 244
rect -1217 -244 -1214 244
rect -1237 -250 -1214 -244
rect -1108 244 -1085 250
rect -1108 -244 -1105 244
rect -1088 -244 -1085 244
rect -1108 -250 -1085 -244
rect -979 244 -956 250
rect -979 -244 -976 244
rect -959 -244 -956 244
rect -979 -250 -956 -244
rect -850 244 -827 250
rect -850 -244 -847 244
rect -830 -244 -827 244
rect -850 -250 -827 -244
rect -721 244 -698 250
rect -721 -244 -718 244
rect -701 -244 -698 244
rect -721 -250 -698 -244
rect -592 244 -569 250
rect -592 -244 -589 244
rect -572 -244 -569 244
rect -592 -250 -569 -244
rect -463 244 -440 250
rect -463 -244 -460 244
rect -443 -244 -440 244
rect -463 -250 -440 -244
rect -334 244 -311 250
rect -334 -244 -331 244
rect -314 -244 -311 244
rect -334 -250 -311 -244
rect -205 244 -182 250
rect -205 -244 -202 244
rect -185 -244 -182 244
rect -205 -250 -182 -244
rect -76 244 -53 250
rect -76 -244 -73 244
rect -56 -244 -53 244
rect -76 -250 -53 -244
rect 53 244 76 250
rect 53 -244 56 244
rect 73 -244 76 244
rect 53 -250 76 -244
rect 182 244 205 250
rect 182 -244 185 244
rect 202 -244 205 244
rect 182 -250 205 -244
rect 311 244 334 250
rect 311 -244 314 244
rect 331 -244 334 244
rect 311 -250 334 -244
rect 440 244 463 250
rect 440 -244 443 244
rect 460 -244 463 244
rect 440 -250 463 -244
rect 569 244 592 250
rect 569 -244 572 244
rect 589 -244 592 244
rect 569 -250 592 -244
rect 698 244 721 250
rect 698 -244 701 244
rect 718 -244 721 244
rect 698 -250 721 -244
rect 827 244 850 250
rect 827 -244 830 244
rect 847 -244 850 244
rect 827 -250 850 -244
rect 956 244 979 250
rect 956 -244 959 244
rect 976 -244 979 244
rect 956 -250 979 -244
rect 1085 244 1108 250
rect 1085 -244 1088 244
rect 1105 -244 1108 244
rect 1085 -250 1108 -244
rect 1214 244 1237 250
rect 1214 -244 1217 244
rect 1234 -244 1237 244
rect 1214 -250 1237 -244
rect 1343 244 1366 250
rect 1343 -244 1346 244
rect 1363 -244 1366 244
rect 1343 -250 1366 -244
rect 1472 244 1495 250
rect 1472 -244 1475 244
rect 1492 -244 1495 244
rect 1472 -250 1495 -244
rect -1467 -269 -1371 -266
rect -1467 -286 -1461 -269
rect -1377 -286 -1371 -269
rect -1467 -289 -1371 -286
rect -1338 -269 -1242 -266
rect -1338 -286 -1332 -269
rect -1248 -286 -1242 -269
rect -1338 -289 -1242 -286
rect -1209 -269 -1113 -266
rect -1209 -286 -1203 -269
rect -1119 -286 -1113 -269
rect -1209 -289 -1113 -286
rect -1080 -269 -984 -266
rect -1080 -286 -1074 -269
rect -990 -286 -984 -269
rect -1080 -289 -984 -286
rect -951 -269 -855 -266
rect -951 -286 -945 -269
rect -861 -286 -855 -269
rect -951 -289 -855 -286
rect -822 -269 -726 -266
rect -822 -286 -816 -269
rect -732 -286 -726 -269
rect -822 -289 -726 -286
rect -693 -269 -597 -266
rect -693 -286 -687 -269
rect -603 -286 -597 -269
rect -693 -289 -597 -286
rect -564 -269 -468 -266
rect -564 -286 -558 -269
rect -474 -286 -468 -269
rect -564 -289 -468 -286
rect -435 -269 -339 -266
rect -435 -286 -429 -269
rect -345 -286 -339 -269
rect -435 -289 -339 -286
rect -306 -269 -210 -266
rect -306 -286 -300 -269
rect -216 -286 -210 -269
rect -306 -289 -210 -286
rect -177 -269 -81 -266
rect -177 -286 -171 -269
rect -87 -286 -81 -269
rect -177 -289 -81 -286
rect -48 -269 48 -266
rect -48 -286 -42 -269
rect 42 -286 48 -269
rect -48 -289 48 -286
rect 81 -269 177 -266
rect 81 -286 87 -269
rect 171 -286 177 -269
rect 81 -289 177 -286
rect 210 -269 306 -266
rect 210 -286 216 -269
rect 300 -286 306 -269
rect 210 -289 306 -286
rect 339 -269 435 -266
rect 339 -286 345 -269
rect 429 -286 435 -269
rect 339 -289 435 -286
rect 468 -269 564 -266
rect 468 -286 474 -269
rect 558 -286 564 -269
rect 468 -289 564 -286
rect 597 -269 693 -266
rect 597 -286 603 -269
rect 687 -286 693 -269
rect 597 -289 693 -286
rect 726 -269 822 -266
rect 726 -286 732 -269
rect 816 -286 822 -269
rect 726 -289 822 -286
rect 855 -269 951 -266
rect 855 -286 861 -269
rect 945 -286 951 -269
rect 855 -289 951 -286
rect 984 -269 1080 -266
rect 984 -286 990 -269
rect 1074 -286 1080 -269
rect 984 -289 1080 -286
rect 1113 -269 1209 -266
rect 1113 -286 1119 -269
rect 1203 -286 1209 -269
rect 1113 -289 1209 -286
rect 1242 -269 1338 -266
rect 1242 -286 1248 -269
rect 1332 -286 1338 -269
rect 1242 -289 1338 -286
rect 1371 -269 1467 -266
rect 1371 -286 1377 -269
rect 1461 -286 1467 -269
rect 1371 -289 1467 -286
rect -1495 -311 -1472 -305
rect -1495 -799 -1492 -311
rect -1475 -799 -1472 -311
rect -1495 -805 -1472 -799
rect -1366 -311 -1343 -305
rect -1366 -799 -1363 -311
rect -1346 -799 -1343 -311
rect -1366 -805 -1343 -799
rect -1237 -311 -1214 -305
rect -1237 -799 -1234 -311
rect -1217 -799 -1214 -311
rect -1237 -805 -1214 -799
rect -1108 -311 -1085 -305
rect -1108 -799 -1105 -311
rect -1088 -799 -1085 -311
rect -1108 -805 -1085 -799
rect -979 -311 -956 -305
rect -979 -799 -976 -311
rect -959 -799 -956 -311
rect -979 -805 -956 -799
rect -850 -311 -827 -305
rect -850 -799 -847 -311
rect -830 -799 -827 -311
rect -850 -805 -827 -799
rect -721 -311 -698 -305
rect -721 -799 -718 -311
rect -701 -799 -698 -311
rect -721 -805 -698 -799
rect -592 -311 -569 -305
rect -592 -799 -589 -311
rect -572 -799 -569 -311
rect -592 -805 -569 -799
rect -463 -311 -440 -305
rect -463 -799 -460 -311
rect -443 -799 -440 -311
rect -463 -805 -440 -799
rect -334 -311 -311 -305
rect -334 -799 -331 -311
rect -314 -799 -311 -311
rect -334 -805 -311 -799
rect -205 -311 -182 -305
rect -205 -799 -202 -311
rect -185 -799 -182 -311
rect -205 -805 -182 -799
rect -76 -311 -53 -305
rect -76 -799 -73 -311
rect -56 -799 -53 -311
rect -76 -805 -53 -799
rect 53 -311 76 -305
rect 53 -799 56 -311
rect 73 -799 76 -311
rect 53 -805 76 -799
rect 182 -311 205 -305
rect 182 -799 185 -311
rect 202 -799 205 -311
rect 182 -805 205 -799
rect 311 -311 334 -305
rect 311 -799 314 -311
rect 331 -799 334 -311
rect 311 -805 334 -799
rect 440 -311 463 -305
rect 440 -799 443 -311
rect 460 -799 463 -311
rect 440 -805 463 -799
rect 569 -311 592 -305
rect 569 -799 572 -311
rect 589 -799 592 -311
rect 569 -805 592 -799
rect 698 -311 721 -305
rect 698 -799 701 -311
rect 718 -799 721 -311
rect 698 -805 721 -799
rect 827 -311 850 -305
rect 827 -799 830 -311
rect 847 -799 850 -311
rect 827 -805 850 -799
rect 956 -311 979 -305
rect 956 -799 959 -311
rect 976 -799 979 -311
rect 956 -805 979 -799
rect 1085 -311 1108 -305
rect 1085 -799 1088 -311
rect 1105 -799 1108 -311
rect 1085 -805 1108 -799
rect 1214 -311 1237 -305
rect 1214 -799 1217 -311
rect 1234 -799 1237 -311
rect 1214 -805 1237 -799
rect 1343 -311 1366 -305
rect 1343 -799 1346 -311
rect 1363 -799 1366 -311
rect 1343 -805 1366 -799
rect 1472 -311 1495 -305
rect 1472 -799 1475 -311
rect 1492 -799 1495 -311
rect 1472 -805 1495 -799
rect -1467 -824 -1371 -821
rect -1467 -841 -1461 -824
rect -1377 -841 -1371 -824
rect -1467 -844 -1371 -841
rect -1338 -824 -1242 -821
rect -1338 -841 -1332 -824
rect -1248 -841 -1242 -824
rect -1338 -844 -1242 -841
rect -1209 -824 -1113 -821
rect -1209 -841 -1203 -824
rect -1119 -841 -1113 -824
rect -1209 -844 -1113 -841
rect -1080 -824 -984 -821
rect -1080 -841 -1074 -824
rect -990 -841 -984 -824
rect -1080 -844 -984 -841
rect -951 -824 -855 -821
rect -951 -841 -945 -824
rect -861 -841 -855 -824
rect -951 -844 -855 -841
rect -822 -824 -726 -821
rect -822 -841 -816 -824
rect -732 -841 -726 -824
rect -822 -844 -726 -841
rect -693 -824 -597 -821
rect -693 -841 -687 -824
rect -603 -841 -597 -824
rect -693 -844 -597 -841
rect -564 -824 -468 -821
rect -564 -841 -558 -824
rect -474 -841 -468 -824
rect -564 -844 -468 -841
rect -435 -824 -339 -821
rect -435 -841 -429 -824
rect -345 -841 -339 -824
rect -435 -844 -339 -841
rect -306 -824 -210 -821
rect -306 -841 -300 -824
rect -216 -841 -210 -824
rect -306 -844 -210 -841
rect -177 -824 -81 -821
rect -177 -841 -171 -824
rect -87 -841 -81 -824
rect -177 -844 -81 -841
rect -48 -824 48 -821
rect -48 -841 -42 -824
rect 42 -841 48 -824
rect -48 -844 48 -841
rect 81 -824 177 -821
rect 81 -841 87 -824
rect 171 -841 177 -824
rect 81 -844 177 -841
rect 210 -824 306 -821
rect 210 -841 216 -824
rect 300 -841 306 -824
rect 210 -844 306 -841
rect 339 -824 435 -821
rect 339 -841 345 -824
rect 429 -841 435 -824
rect 339 -844 435 -841
rect 468 -824 564 -821
rect 468 -841 474 -824
rect 558 -841 564 -824
rect 468 -844 564 -841
rect 597 -824 693 -821
rect 597 -841 603 -824
rect 687 -841 693 -824
rect 597 -844 693 -841
rect 726 -824 822 -821
rect 726 -841 732 -824
rect 816 -841 822 -824
rect 726 -844 822 -841
rect 855 -824 951 -821
rect 855 -841 861 -824
rect 945 -841 951 -824
rect 855 -844 951 -841
rect 984 -824 1080 -821
rect 984 -841 990 -824
rect 1074 -841 1080 -824
rect 984 -844 1080 -841
rect 1113 -824 1209 -821
rect 1113 -841 1119 -824
rect 1203 -841 1209 -824
rect 1113 -844 1209 -841
rect 1242 -824 1338 -821
rect 1242 -841 1248 -824
rect 1332 -841 1338 -824
rect 1242 -844 1338 -841
rect 1371 -824 1467 -821
rect 1371 -841 1377 -824
rect 1461 -841 1467 -824
rect 1371 -844 1467 -841
rect -1495 -866 -1472 -860
rect -1495 -1354 -1492 -866
rect -1475 -1354 -1472 -866
rect -1495 -1360 -1472 -1354
rect -1366 -866 -1343 -860
rect -1366 -1354 -1363 -866
rect -1346 -1354 -1343 -866
rect -1366 -1360 -1343 -1354
rect -1237 -866 -1214 -860
rect -1237 -1354 -1234 -866
rect -1217 -1354 -1214 -866
rect -1237 -1360 -1214 -1354
rect -1108 -866 -1085 -860
rect -1108 -1354 -1105 -866
rect -1088 -1354 -1085 -866
rect -1108 -1360 -1085 -1354
rect -979 -866 -956 -860
rect -979 -1354 -976 -866
rect -959 -1354 -956 -866
rect -979 -1360 -956 -1354
rect -850 -866 -827 -860
rect -850 -1354 -847 -866
rect -830 -1354 -827 -866
rect -850 -1360 -827 -1354
rect -721 -866 -698 -860
rect -721 -1354 -718 -866
rect -701 -1354 -698 -866
rect -721 -1360 -698 -1354
rect -592 -866 -569 -860
rect -592 -1354 -589 -866
rect -572 -1354 -569 -866
rect -592 -1360 -569 -1354
rect -463 -866 -440 -860
rect -463 -1354 -460 -866
rect -443 -1354 -440 -866
rect -463 -1360 -440 -1354
rect -334 -866 -311 -860
rect -334 -1354 -331 -866
rect -314 -1354 -311 -866
rect -334 -1360 -311 -1354
rect -205 -866 -182 -860
rect -205 -1354 -202 -866
rect -185 -1354 -182 -866
rect -205 -1360 -182 -1354
rect -76 -866 -53 -860
rect -76 -1354 -73 -866
rect -56 -1354 -53 -866
rect -76 -1360 -53 -1354
rect 53 -866 76 -860
rect 53 -1354 56 -866
rect 73 -1354 76 -866
rect 53 -1360 76 -1354
rect 182 -866 205 -860
rect 182 -1354 185 -866
rect 202 -1354 205 -866
rect 182 -1360 205 -1354
rect 311 -866 334 -860
rect 311 -1354 314 -866
rect 331 -1354 334 -866
rect 311 -1360 334 -1354
rect 440 -866 463 -860
rect 440 -1354 443 -866
rect 460 -1354 463 -866
rect 440 -1360 463 -1354
rect 569 -866 592 -860
rect 569 -1354 572 -866
rect 589 -1354 592 -866
rect 569 -1360 592 -1354
rect 698 -866 721 -860
rect 698 -1354 701 -866
rect 718 -1354 721 -866
rect 698 -1360 721 -1354
rect 827 -866 850 -860
rect 827 -1354 830 -866
rect 847 -1354 850 -866
rect 827 -1360 850 -1354
rect 956 -866 979 -860
rect 956 -1354 959 -866
rect 976 -1354 979 -866
rect 956 -1360 979 -1354
rect 1085 -866 1108 -860
rect 1085 -1354 1088 -866
rect 1105 -1354 1108 -866
rect 1085 -1360 1108 -1354
rect 1214 -866 1237 -860
rect 1214 -1354 1217 -866
rect 1234 -1354 1237 -866
rect 1214 -1360 1237 -1354
rect 1343 -866 1366 -860
rect 1343 -1354 1346 -866
rect 1363 -1354 1366 -866
rect 1343 -1360 1366 -1354
rect 1472 -866 1495 -860
rect 1472 -1354 1475 -866
rect 1492 -1354 1495 -866
rect 1472 -1360 1495 -1354
rect -1467 -1379 -1371 -1376
rect -1467 -1396 -1461 -1379
rect -1377 -1396 -1371 -1379
rect -1467 -1399 -1371 -1396
rect -1338 -1379 -1242 -1376
rect -1338 -1396 -1332 -1379
rect -1248 -1396 -1242 -1379
rect -1338 -1399 -1242 -1396
rect -1209 -1379 -1113 -1376
rect -1209 -1396 -1203 -1379
rect -1119 -1396 -1113 -1379
rect -1209 -1399 -1113 -1396
rect -1080 -1379 -984 -1376
rect -1080 -1396 -1074 -1379
rect -990 -1396 -984 -1379
rect -1080 -1399 -984 -1396
rect -951 -1379 -855 -1376
rect -951 -1396 -945 -1379
rect -861 -1396 -855 -1379
rect -951 -1399 -855 -1396
rect -822 -1379 -726 -1376
rect -822 -1396 -816 -1379
rect -732 -1396 -726 -1379
rect -822 -1399 -726 -1396
rect -693 -1379 -597 -1376
rect -693 -1396 -687 -1379
rect -603 -1396 -597 -1379
rect -693 -1399 -597 -1396
rect -564 -1379 -468 -1376
rect -564 -1396 -558 -1379
rect -474 -1396 -468 -1379
rect -564 -1399 -468 -1396
rect -435 -1379 -339 -1376
rect -435 -1396 -429 -1379
rect -345 -1396 -339 -1379
rect -435 -1399 -339 -1396
rect -306 -1379 -210 -1376
rect -306 -1396 -300 -1379
rect -216 -1396 -210 -1379
rect -306 -1399 -210 -1396
rect -177 -1379 -81 -1376
rect -177 -1396 -171 -1379
rect -87 -1396 -81 -1379
rect -177 -1399 -81 -1396
rect -48 -1379 48 -1376
rect -48 -1396 -42 -1379
rect 42 -1396 48 -1379
rect -48 -1399 48 -1396
rect 81 -1379 177 -1376
rect 81 -1396 87 -1379
rect 171 -1396 177 -1379
rect 81 -1399 177 -1396
rect 210 -1379 306 -1376
rect 210 -1396 216 -1379
rect 300 -1396 306 -1379
rect 210 -1399 306 -1396
rect 339 -1379 435 -1376
rect 339 -1396 345 -1379
rect 429 -1396 435 -1379
rect 339 -1399 435 -1396
rect 468 -1379 564 -1376
rect 468 -1396 474 -1379
rect 558 -1396 564 -1379
rect 468 -1399 564 -1396
rect 597 -1379 693 -1376
rect 597 -1396 603 -1379
rect 687 -1396 693 -1379
rect 597 -1399 693 -1396
rect 726 -1379 822 -1376
rect 726 -1396 732 -1379
rect 816 -1396 822 -1379
rect 726 -1399 822 -1396
rect 855 -1379 951 -1376
rect 855 -1396 861 -1379
rect 945 -1396 951 -1379
rect 855 -1399 951 -1396
rect 984 -1379 1080 -1376
rect 984 -1396 990 -1379
rect 1074 -1396 1080 -1379
rect 984 -1399 1080 -1396
rect 1113 -1379 1209 -1376
rect 1113 -1396 1119 -1379
rect 1203 -1396 1209 -1379
rect 1113 -1399 1209 -1396
rect 1242 -1379 1338 -1376
rect 1242 -1396 1248 -1379
rect 1332 -1396 1338 -1379
rect 1242 -1399 1338 -1396
rect 1371 -1379 1467 -1376
rect 1371 -1396 1377 -1379
rect 1461 -1396 1467 -1379
rect 1371 -1399 1467 -1396
<< properties >>
string FIXED_BBOX -1550 -1456 1550 1456
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 1.0 m 5 nf 23 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
