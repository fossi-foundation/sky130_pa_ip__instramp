magic
tech sky130A
magscale 1 2
timestamp 1730992408
<< pwell >>
rect -4434 -2307 4434 2307
<< psubdiff >>
rect -4398 2237 -4302 2271
rect 4302 2237 4398 2271
rect -4398 2175 -4364 2237
rect 4364 2175 4398 2237
rect -4398 -2237 -4364 -2175
rect 4364 -2237 4398 -2175
rect -4398 -2271 -4302 -2237
rect 4302 -2271 4398 -2237
<< psubdiffcont >>
rect -4302 2237 4302 2271
rect -4398 -2175 -4364 2175
rect 4364 -2175 4398 2175
rect -4302 -2271 4302 -2237
<< xpolycontact >>
rect -4268 1709 -4198 2141
rect -4268 -2141 -4198 -1709
rect -4102 1709 -4032 2141
rect -4102 -2141 -4032 -1709
rect -3936 1709 -3866 2141
rect -3936 -2141 -3866 -1709
rect -3770 1709 -3700 2141
rect -3770 -2141 -3700 -1709
rect -3604 1709 -3534 2141
rect -3604 -2141 -3534 -1709
rect -3438 1709 -3368 2141
rect -3438 -2141 -3368 -1709
rect -3272 1709 -3202 2141
rect -3272 -2141 -3202 -1709
rect -3106 1709 -3036 2141
rect -3106 -2141 -3036 -1709
rect -2940 1709 -2870 2141
rect -2940 -2141 -2870 -1709
rect -2774 1709 -2704 2141
rect -2774 -2141 -2704 -1709
rect -2608 1709 -2538 2141
rect -2608 -2141 -2538 -1709
rect -2442 1709 -2372 2141
rect -2442 -2141 -2372 -1709
rect -2276 1709 -2206 2141
rect -2276 -2141 -2206 -1709
rect -2110 1709 -2040 2141
rect -2110 -2141 -2040 -1709
rect -1944 1709 -1874 2141
rect -1944 -2141 -1874 -1709
rect -1778 1709 -1708 2141
rect -1778 -2141 -1708 -1709
rect -1612 1709 -1542 2141
rect -1612 -2141 -1542 -1709
rect -1446 1709 -1376 2141
rect -1446 -2141 -1376 -1709
rect -1280 1709 -1210 2141
rect -1280 -2141 -1210 -1709
rect -1114 1709 -1044 2141
rect -1114 -2141 -1044 -1709
rect -948 1709 -878 2141
rect -948 -2141 -878 -1709
rect -782 1709 -712 2141
rect -782 -2141 -712 -1709
rect -616 1709 -546 2141
rect -616 -2141 -546 -1709
rect -450 1709 -380 2141
rect -450 -2141 -380 -1709
rect -284 1709 -214 2141
rect -284 -2141 -214 -1709
rect -118 1709 -48 2141
rect -118 -2141 -48 -1709
rect 48 1709 118 2141
rect 48 -2141 118 -1709
rect 214 1709 284 2141
rect 214 -2141 284 -1709
rect 380 1709 450 2141
rect 380 -2141 450 -1709
rect 546 1709 616 2141
rect 546 -2141 616 -1709
rect 712 1709 782 2141
rect 712 -2141 782 -1709
rect 878 1709 948 2141
rect 878 -2141 948 -1709
rect 1044 1709 1114 2141
rect 1044 -2141 1114 -1709
rect 1210 1709 1280 2141
rect 1210 -2141 1280 -1709
rect 1376 1709 1446 2141
rect 1376 -2141 1446 -1709
rect 1542 1709 1612 2141
rect 1542 -2141 1612 -1709
rect 1708 1709 1778 2141
rect 1708 -2141 1778 -1709
rect 1874 1709 1944 2141
rect 1874 -2141 1944 -1709
rect 2040 1709 2110 2141
rect 2040 -2141 2110 -1709
rect 2206 1709 2276 2141
rect 2206 -2141 2276 -1709
rect 2372 1709 2442 2141
rect 2372 -2141 2442 -1709
rect 2538 1709 2608 2141
rect 2538 -2141 2608 -1709
rect 2704 1709 2774 2141
rect 2704 -2141 2774 -1709
rect 2870 1709 2940 2141
rect 2870 -2141 2940 -1709
rect 3036 1709 3106 2141
rect 3036 -2141 3106 -1709
rect 3202 1709 3272 2141
rect 3202 -2141 3272 -1709
rect 3368 1709 3438 2141
rect 3368 -2141 3438 -1709
rect 3534 1709 3604 2141
rect 3534 -2141 3604 -1709
rect 3700 1709 3770 2141
rect 3700 -2141 3770 -1709
rect 3866 1709 3936 2141
rect 3866 -2141 3936 -1709
rect 4032 1709 4102 2141
rect 4032 -2141 4102 -1709
rect 4198 1709 4268 2141
rect 4198 -2141 4268 -1709
<< xpolyres >>
rect -4268 -1709 -4198 1709
rect -4102 -1709 -4032 1709
rect -3936 -1709 -3866 1709
rect -3770 -1709 -3700 1709
rect -3604 -1709 -3534 1709
rect -3438 -1709 -3368 1709
rect -3272 -1709 -3202 1709
rect -3106 -1709 -3036 1709
rect -2940 -1709 -2870 1709
rect -2774 -1709 -2704 1709
rect -2608 -1709 -2538 1709
rect -2442 -1709 -2372 1709
rect -2276 -1709 -2206 1709
rect -2110 -1709 -2040 1709
rect -1944 -1709 -1874 1709
rect -1778 -1709 -1708 1709
rect -1612 -1709 -1542 1709
rect -1446 -1709 -1376 1709
rect -1280 -1709 -1210 1709
rect -1114 -1709 -1044 1709
rect -948 -1709 -878 1709
rect -782 -1709 -712 1709
rect -616 -1709 -546 1709
rect -450 -1709 -380 1709
rect -284 -1709 -214 1709
rect -118 -1709 -48 1709
rect 48 -1709 118 1709
rect 214 -1709 284 1709
rect 380 -1709 450 1709
rect 546 -1709 616 1709
rect 712 -1709 782 1709
rect 878 -1709 948 1709
rect 1044 -1709 1114 1709
rect 1210 -1709 1280 1709
rect 1376 -1709 1446 1709
rect 1542 -1709 1612 1709
rect 1708 -1709 1778 1709
rect 1874 -1709 1944 1709
rect 2040 -1709 2110 1709
rect 2206 -1709 2276 1709
rect 2372 -1709 2442 1709
rect 2538 -1709 2608 1709
rect 2704 -1709 2774 1709
rect 2870 -1709 2940 1709
rect 3036 -1709 3106 1709
rect 3202 -1709 3272 1709
rect 3368 -1709 3438 1709
rect 3534 -1709 3604 1709
rect 3700 -1709 3770 1709
rect 3866 -1709 3936 1709
rect 4032 -1709 4102 1709
rect 4198 -1709 4268 1709
<< locali >>
rect -4398 2237 -4302 2271
rect 4302 2237 4398 2271
rect -4398 2175 -4364 2237
rect 4364 2175 4398 2237
rect -4398 -2237 -4364 -2175
rect 4364 -2237 4398 -2175
rect -4398 -2271 -4302 -2237
rect 4302 -2271 4398 -2237
<< viali >>
rect -4252 1726 -4214 2123
rect -4086 1726 -4048 2123
rect -3920 1726 -3882 2123
rect -3754 1726 -3716 2123
rect -3588 1726 -3550 2123
rect -3422 1726 -3384 2123
rect -3256 1726 -3218 2123
rect -3090 1726 -3052 2123
rect -2924 1726 -2886 2123
rect -2758 1726 -2720 2123
rect -2592 1726 -2554 2123
rect -2426 1726 -2388 2123
rect -2260 1726 -2222 2123
rect -2094 1726 -2056 2123
rect -1928 1726 -1890 2123
rect -1762 1726 -1724 2123
rect -1596 1726 -1558 2123
rect -1430 1726 -1392 2123
rect -1264 1726 -1226 2123
rect -1098 1726 -1060 2123
rect -932 1726 -894 2123
rect -766 1726 -728 2123
rect -600 1726 -562 2123
rect -434 1726 -396 2123
rect -268 1726 -230 2123
rect -102 1726 -64 2123
rect 64 1726 102 2123
rect 230 1726 268 2123
rect 396 1726 434 2123
rect 562 1726 600 2123
rect 728 1726 766 2123
rect 894 1726 932 2123
rect 1060 1726 1098 2123
rect 1226 1726 1264 2123
rect 1392 1726 1430 2123
rect 1558 1726 1596 2123
rect 1724 1726 1762 2123
rect 1890 1726 1928 2123
rect 2056 1726 2094 2123
rect 2222 1726 2260 2123
rect 2388 1726 2426 2123
rect 2554 1726 2592 2123
rect 2720 1726 2758 2123
rect 2886 1726 2924 2123
rect 3052 1726 3090 2123
rect 3218 1726 3256 2123
rect 3384 1726 3422 2123
rect 3550 1726 3588 2123
rect 3716 1726 3754 2123
rect 3882 1726 3920 2123
rect 4048 1726 4086 2123
rect 4214 1726 4252 2123
rect -4252 -2123 -4214 -1726
rect -4086 -2123 -4048 -1726
rect -3920 -2123 -3882 -1726
rect -3754 -2123 -3716 -1726
rect -3588 -2123 -3550 -1726
rect -3422 -2123 -3384 -1726
rect -3256 -2123 -3218 -1726
rect -3090 -2123 -3052 -1726
rect -2924 -2123 -2886 -1726
rect -2758 -2123 -2720 -1726
rect -2592 -2123 -2554 -1726
rect -2426 -2123 -2388 -1726
rect -2260 -2123 -2222 -1726
rect -2094 -2123 -2056 -1726
rect -1928 -2123 -1890 -1726
rect -1762 -2123 -1724 -1726
rect -1596 -2123 -1558 -1726
rect -1430 -2123 -1392 -1726
rect -1264 -2123 -1226 -1726
rect -1098 -2123 -1060 -1726
rect -932 -2123 -894 -1726
rect -766 -2123 -728 -1726
rect -600 -2123 -562 -1726
rect -434 -2123 -396 -1726
rect -268 -2123 -230 -1726
rect -102 -2123 -64 -1726
rect 64 -2123 102 -1726
rect 230 -2123 268 -1726
rect 396 -2123 434 -1726
rect 562 -2123 600 -1726
rect 728 -2123 766 -1726
rect 894 -2123 932 -1726
rect 1060 -2123 1098 -1726
rect 1226 -2123 1264 -1726
rect 1392 -2123 1430 -1726
rect 1558 -2123 1596 -1726
rect 1724 -2123 1762 -1726
rect 1890 -2123 1928 -1726
rect 2056 -2123 2094 -1726
rect 2222 -2123 2260 -1726
rect 2388 -2123 2426 -1726
rect 2554 -2123 2592 -1726
rect 2720 -2123 2758 -1726
rect 2886 -2123 2924 -1726
rect 3052 -2123 3090 -1726
rect 3218 -2123 3256 -1726
rect 3384 -2123 3422 -1726
rect 3550 -2123 3588 -1726
rect 3716 -2123 3754 -1726
rect 3882 -2123 3920 -1726
rect 4048 -2123 4086 -1726
rect 4214 -2123 4252 -1726
<< metal1 >>
rect -4258 2123 -4208 2135
rect -4258 1726 -4252 2123
rect -4214 1726 -4208 2123
rect -4258 1714 -4208 1726
rect -4092 2123 -4042 2135
rect -4092 1726 -4086 2123
rect -4048 1726 -4042 2123
rect -4092 1714 -4042 1726
rect -3926 2123 -3876 2135
rect -3926 1726 -3920 2123
rect -3882 1726 -3876 2123
rect -3926 1714 -3876 1726
rect -3760 2123 -3710 2135
rect -3760 1726 -3754 2123
rect -3716 1726 -3710 2123
rect -3760 1714 -3710 1726
rect -3594 2123 -3544 2135
rect -3594 1726 -3588 2123
rect -3550 1726 -3544 2123
rect -3594 1714 -3544 1726
rect -3428 2123 -3378 2135
rect -3428 1726 -3422 2123
rect -3384 1726 -3378 2123
rect -3428 1714 -3378 1726
rect -3262 2123 -3212 2135
rect -3262 1726 -3256 2123
rect -3218 1726 -3212 2123
rect -3262 1714 -3212 1726
rect -3096 2123 -3046 2135
rect -3096 1726 -3090 2123
rect -3052 1726 -3046 2123
rect -3096 1714 -3046 1726
rect -2930 2123 -2880 2135
rect -2930 1726 -2924 2123
rect -2886 1726 -2880 2123
rect -2930 1714 -2880 1726
rect -2764 2123 -2714 2135
rect -2764 1726 -2758 2123
rect -2720 1726 -2714 2123
rect -2764 1714 -2714 1726
rect -2598 2123 -2548 2135
rect -2598 1726 -2592 2123
rect -2554 1726 -2548 2123
rect -2598 1714 -2548 1726
rect -2432 2123 -2382 2135
rect -2432 1726 -2426 2123
rect -2388 1726 -2382 2123
rect -2432 1714 -2382 1726
rect -2266 2123 -2216 2135
rect -2266 1726 -2260 2123
rect -2222 1726 -2216 2123
rect -2266 1714 -2216 1726
rect -2100 2123 -2050 2135
rect -2100 1726 -2094 2123
rect -2056 1726 -2050 2123
rect -2100 1714 -2050 1726
rect -1934 2123 -1884 2135
rect -1934 1726 -1928 2123
rect -1890 1726 -1884 2123
rect -1934 1714 -1884 1726
rect -1768 2123 -1718 2135
rect -1768 1726 -1762 2123
rect -1724 1726 -1718 2123
rect -1768 1714 -1718 1726
rect -1602 2123 -1552 2135
rect -1602 1726 -1596 2123
rect -1558 1726 -1552 2123
rect -1602 1714 -1552 1726
rect -1436 2123 -1386 2135
rect -1436 1726 -1430 2123
rect -1392 1726 -1386 2123
rect -1436 1714 -1386 1726
rect -1270 2123 -1220 2135
rect -1270 1726 -1264 2123
rect -1226 1726 -1220 2123
rect -1270 1714 -1220 1726
rect -1104 2123 -1054 2135
rect -1104 1726 -1098 2123
rect -1060 1726 -1054 2123
rect -1104 1714 -1054 1726
rect -938 2123 -888 2135
rect -938 1726 -932 2123
rect -894 1726 -888 2123
rect -938 1714 -888 1726
rect -772 2123 -722 2135
rect -772 1726 -766 2123
rect -728 1726 -722 2123
rect -772 1714 -722 1726
rect -606 2123 -556 2135
rect -606 1726 -600 2123
rect -562 1726 -556 2123
rect -606 1714 -556 1726
rect -440 2123 -390 2135
rect -440 1726 -434 2123
rect -396 1726 -390 2123
rect -440 1714 -390 1726
rect -274 2123 -224 2135
rect -274 1726 -268 2123
rect -230 1726 -224 2123
rect -274 1714 -224 1726
rect -108 2123 -58 2135
rect -108 1726 -102 2123
rect -64 1726 -58 2123
rect -108 1714 -58 1726
rect 58 2123 108 2135
rect 58 1726 64 2123
rect 102 1726 108 2123
rect 58 1714 108 1726
rect 224 2123 274 2135
rect 224 1726 230 2123
rect 268 1726 274 2123
rect 224 1714 274 1726
rect 390 2123 440 2135
rect 390 1726 396 2123
rect 434 1726 440 2123
rect 390 1714 440 1726
rect 556 2123 606 2135
rect 556 1726 562 2123
rect 600 1726 606 2123
rect 556 1714 606 1726
rect 722 2123 772 2135
rect 722 1726 728 2123
rect 766 1726 772 2123
rect 722 1714 772 1726
rect 888 2123 938 2135
rect 888 1726 894 2123
rect 932 1726 938 2123
rect 888 1714 938 1726
rect 1054 2123 1104 2135
rect 1054 1726 1060 2123
rect 1098 1726 1104 2123
rect 1054 1714 1104 1726
rect 1220 2123 1270 2135
rect 1220 1726 1226 2123
rect 1264 1726 1270 2123
rect 1220 1714 1270 1726
rect 1386 2123 1436 2135
rect 1386 1726 1392 2123
rect 1430 1726 1436 2123
rect 1386 1714 1436 1726
rect 1552 2123 1602 2135
rect 1552 1726 1558 2123
rect 1596 1726 1602 2123
rect 1552 1714 1602 1726
rect 1718 2123 1768 2135
rect 1718 1726 1724 2123
rect 1762 1726 1768 2123
rect 1718 1714 1768 1726
rect 1884 2123 1934 2135
rect 1884 1726 1890 2123
rect 1928 1726 1934 2123
rect 1884 1714 1934 1726
rect 2050 2123 2100 2135
rect 2050 1726 2056 2123
rect 2094 1726 2100 2123
rect 2050 1714 2100 1726
rect 2216 2123 2266 2135
rect 2216 1726 2222 2123
rect 2260 1726 2266 2123
rect 2216 1714 2266 1726
rect 2382 2123 2432 2135
rect 2382 1726 2388 2123
rect 2426 1726 2432 2123
rect 2382 1714 2432 1726
rect 2548 2123 2598 2135
rect 2548 1726 2554 2123
rect 2592 1726 2598 2123
rect 2548 1714 2598 1726
rect 2714 2123 2764 2135
rect 2714 1726 2720 2123
rect 2758 1726 2764 2123
rect 2714 1714 2764 1726
rect 2880 2123 2930 2135
rect 2880 1726 2886 2123
rect 2924 1726 2930 2123
rect 2880 1714 2930 1726
rect 3046 2123 3096 2135
rect 3046 1726 3052 2123
rect 3090 1726 3096 2123
rect 3046 1714 3096 1726
rect 3212 2123 3262 2135
rect 3212 1726 3218 2123
rect 3256 1726 3262 2123
rect 3212 1714 3262 1726
rect 3378 2123 3428 2135
rect 3378 1726 3384 2123
rect 3422 1726 3428 2123
rect 3378 1714 3428 1726
rect 3544 2123 3594 2135
rect 3544 1726 3550 2123
rect 3588 1726 3594 2123
rect 3544 1714 3594 1726
rect 3710 2123 3760 2135
rect 3710 1726 3716 2123
rect 3754 1726 3760 2123
rect 3710 1714 3760 1726
rect 3876 2123 3926 2135
rect 3876 1726 3882 2123
rect 3920 1726 3926 2123
rect 3876 1714 3926 1726
rect 4042 2123 4092 2135
rect 4042 1726 4048 2123
rect 4086 1726 4092 2123
rect 4042 1714 4092 1726
rect 4208 2123 4258 2135
rect 4208 1726 4214 2123
rect 4252 1726 4258 2123
rect 4208 1714 4258 1726
rect -4258 -1726 -4208 -1714
rect -4258 -2123 -4252 -1726
rect -4214 -2123 -4208 -1726
rect -4258 -2135 -4208 -2123
rect -4092 -1726 -4042 -1714
rect -4092 -2123 -4086 -1726
rect -4048 -2123 -4042 -1726
rect -4092 -2135 -4042 -2123
rect -3926 -1726 -3876 -1714
rect -3926 -2123 -3920 -1726
rect -3882 -2123 -3876 -1726
rect -3926 -2135 -3876 -2123
rect -3760 -1726 -3710 -1714
rect -3760 -2123 -3754 -1726
rect -3716 -2123 -3710 -1726
rect -3760 -2135 -3710 -2123
rect -3594 -1726 -3544 -1714
rect -3594 -2123 -3588 -1726
rect -3550 -2123 -3544 -1726
rect -3594 -2135 -3544 -2123
rect -3428 -1726 -3378 -1714
rect -3428 -2123 -3422 -1726
rect -3384 -2123 -3378 -1726
rect -3428 -2135 -3378 -2123
rect -3262 -1726 -3212 -1714
rect -3262 -2123 -3256 -1726
rect -3218 -2123 -3212 -1726
rect -3262 -2135 -3212 -2123
rect -3096 -1726 -3046 -1714
rect -3096 -2123 -3090 -1726
rect -3052 -2123 -3046 -1726
rect -3096 -2135 -3046 -2123
rect -2930 -1726 -2880 -1714
rect -2930 -2123 -2924 -1726
rect -2886 -2123 -2880 -1726
rect -2930 -2135 -2880 -2123
rect -2764 -1726 -2714 -1714
rect -2764 -2123 -2758 -1726
rect -2720 -2123 -2714 -1726
rect -2764 -2135 -2714 -2123
rect -2598 -1726 -2548 -1714
rect -2598 -2123 -2592 -1726
rect -2554 -2123 -2548 -1726
rect -2598 -2135 -2548 -2123
rect -2432 -1726 -2382 -1714
rect -2432 -2123 -2426 -1726
rect -2388 -2123 -2382 -1726
rect -2432 -2135 -2382 -2123
rect -2266 -1726 -2216 -1714
rect -2266 -2123 -2260 -1726
rect -2222 -2123 -2216 -1726
rect -2266 -2135 -2216 -2123
rect -2100 -1726 -2050 -1714
rect -2100 -2123 -2094 -1726
rect -2056 -2123 -2050 -1726
rect -2100 -2135 -2050 -2123
rect -1934 -1726 -1884 -1714
rect -1934 -2123 -1928 -1726
rect -1890 -2123 -1884 -1726
rect -1934 -2135 -1884 -2123
rect -1768 -1726 -1718 -1714
rect -1768 -2123 -1762 -1726
rect -1724 -2123 -1718 -1726
rect -1768 -2135 -1718 -2123
rect -1602 -1726 -1552 -1714
rect -1602 -2123 -1596 -1726
rect -1558 -2123 -1552 -1726
rect -1602 -2135 -1552 -2123
rect -1436 -1726 -1386 -1714
rect -1436 -2123 -1430 -1726
rect -1392 -2123 -1386 -1726
rect -1436 -2135 -1386 -2123
rect -1270 -1726 -1220 -1714
rect -1270 -2123 -1264 -1726
rect -1226 -2123 -1220 -1726
rect -1270 -2135 -1220 -2123
rect -1104 -1726 -1054 -1714
rect -1104 -2123 -1098 -1726
rect -1060 -2123 -1054 -1726
rect -1104 -2135 -1054 -2123
rect -938 -1726 -888 -1714
rect -938 -2123 -932 -1726
rect -894 -2123 -888 -1726
rect -938 -2135 -888 -2123
rect -772 -1726 -722 -1714
rect -772 -2123 -766 -1726
rect -728 -2123 -722 -1726
rect -772 -2135 -722 -2123
rect -606 -1726 -556 -1714
rect -606 -2123 -600 -1726
rect -562 -2123 -556 -1726
rect -606 -2135 -556 -2123
rect -440 -1726 -390 -1714
rect -440 -2123 -434 -1726
rect -396 -2123 -390 -1726
rect -440 -2135 -390 -2123
rect -274 -1726 -224 -1714
rect -274 -2123 -268 -1726
rect -230 -2123 -224 -1726
rect -274 -2135 -224 -2123
rect -108 -1726 -58 -1714
rect -108 -2123 -102 -1726
rect -64 -2123 -58 -1726
rect -108 -2135 -58 -2123
rect 58 -1726 108 -1714
rect 58 -2123 64 -1726
rect 102 -2123 108 -1726
rect 58 -2135 108 -2123
rect 224 -1726 274 -1714
rect 224 -2123 230 -1726
rect 268 -2123 274 -1726
rect 224 -2135 274 -2123
rect 390 -1726 440 -1714
rect 390 -2123 396 -1726
rect 434 -2123 440 -1726
rect 390 -2135 440 -2123
rect 556 -1726 606 -1714
rect 556 -2123 562 -1726
rect 600 -2123 606 -1726
rect 556 -2135 606 -2123
rect 722 -1726 772 -1714
rect 722 -2123 728 -1726
rect 766 -2123 772 -1726
rect 722 -2135 772 -2123
rect 888 -1726 938 -1714
rect 888 -2123 894 -1726
rect 932 -2123 938 -1726
rect 888 -2135 938 -2123
rect 1054 -1726 1104 -1714
rect 1054 -2123 1060 -1726
rect 1098 -2123 1104 -1726
rect 1054 -2135 1104 -2123
rect 1220 -1726 1270 -1714
rect 1220 -2123 1226 -1726
rect 1264 -2123 1270 -1726
rect 1220 -2135 1270 -2123
rect 1386 -1726 1436 -1714
rect 1386 -2123 1392 -1726
rect 1430 -2123 1436 -1726
rect 1386 -2135 1436 -2123
rect 1552 -1726 1602 -1714
rect 1552 -2123 1558 -1726
rect 1596 -2123 1602 -1726
rect 1552 -2135 1602 -2123
rect 1718 -1726 1768 -1714
rect 1718 -2123 1724 -1726
rect 1762 -2123 1768 -1726
rect 1718 -2135 1768 -2123
rect 1884 -1726 1934 -1714
rect 1884 -2123 1890 -1726
rect 1928 -2123 1934 -1726
rect 1884 -2135 1934 -2123
rect 2050 -1726 2100 -1714
rect 2050 -2123 2056 -1726
rect 2094 -2123 2100 -1726
rect 2050 -2135 2100 -2123
rect 2216 -1726 2266 -1714
rect 2216 -2123 2222 -1726
rect 2260 -2123 2266 -1726
rect 2216 -2135 2266 -2123
rect 2382 -1726 2432 -1714
rect 2382 -2123 2388 -1726
rect 2426 -2123 2432 -1726
rect 2382 -2135 2432 -2123
rect 2548 -1726 2598 -1714
rect 2548 -2123 2554 -1726
rect 2592 -2123 2598 -1726
rect 2548 -2135 2598 -2123
rect 2714 -1726 2764 -1714
rect 2714 -2123 2720 -1726
rect 2758 -2123 2764 -1726
rect 2714 -2135 2764 -2123
rect 2880 -1726 2930 -1714
rect 2880 -2123 2886 -1726
rect 2924 -2123 2930 -1726
rect 2880 -2135 2930 -2123
rect 3046 -1726 3096 -1714
rect 3046 -2123 3052 -1726
rect 3090 -2123 3096 -1726
rect 3046 -2135 3096 -2123
rect 3212 -1726 3262 -1714
rect 3212 -2123 3218 -1726
rect 3256 -2123 3262 -1726
rect 3212 -2135 3262 -2123
rect 3378 -1726 3428 -1714
rect 3378 -2123 3384 -1726
rect 3422 -2123 3428 -1726
rect 3378 -2135 3428 -2123
rect 3544 -1726 3594 -1714
rect 3544 -2123 3550 -1726
rect 3588 -2123 3594 -1726
rect 3544 -2135 3594 -2123
rect 3710 -1726 3760 -1714
rect 3710 -2123 3716 -1726
rect 3754 -2123 3760 -1726
rect 3710 -2135 3760 -2123
rect 3876 -1726 3926 -1714
rect 3876 -2123 3882 -1726
rect 3920 -2123 3926 -1726
rect 3876 -2135 3926 -2123
rect 4042 -1726 4092 -1714
rect 4042 -2123 4048 -1726
rect 4086 -2123 4092 -1726
rect 4042 -2135 4092 -2123
rect 4208 -1726 4258 -1714
rect 4208 -2123 4214 -1726
rect 4252 -2123 4258 -1726
rect 4208 -2135 4258 -2123
<< properties >>
string FIXED_BBOX -4381 -2254 4381 2254
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 17.25 m 1 nx 52 wmin 0.350 lmin 0.50 class resistor rho 2000 val 99.646k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
