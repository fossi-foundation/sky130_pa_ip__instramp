magic
tech sky130A
magscale 1 2
timestamp 1729620069
<< pwell >>
rect -23635 -2182 23635 2182
<< psubdiff >>
rect -23599 2112 -23503 2146
rect 23503 2112 23599 2146
rect -23599 2050 -23565 2112
rect 23565 2050 23599 2112
rect -23599 -2112 -23565 -2050
rect 23565 -2112 23599 -2050
rect -23599 -2146 -23503 -2112
rect 23503 -2146 23599 -2112
<< psubdiffcont >>
rect -23503 2112 23503 2146
rect -23599 -2050 -23565 2050
rect 23565 -2050 23599 2050
rect -23503 -2146 23503 -2112
<< xpolycontact >>
rect -23469 1584 -23331 2016
rect -23469 -2016 -23331 -1584
rect -23235 1584 -23097 2016
rect -23235 -2016 -23097 -1584
rect -23001 1584 -22863 2016
rect -23001 -2016 -22863 -1584
rect -22767 1584 -22629 2016
rect -22767 -2016 -22629 -1584
rect -22533 1584 -22395 2016
rect -22533 -2016 -22395 -1584
rect -22299 1584 -22161 2016
rect -22299 -2016 -22161 -1584
rect -22065 1584 -21927 2016
rect -22065 -2016 -21927 -1584
rect -21831 1584 -21693 2016
rect -21831 -2016 -21693 -1584
rect -21597 1584 -21459 2016
rect -21597 -2016 -21459 -1584
rect -21363 1584 -21225 2016
rect -21363 -2016 -21225 -1584
rect -21129 1584 -20991 2016
rect -21129 -2016 -20991 -1584
rect -20895 1584 -20757 2016
rect -20895 -2016 -20757 -1584
rect -20661 1584 -20523 2016
rect -20661 -2016 -20523 -1584
rect -20427 1584 -20289 2016
rect -20427 -2016 -20289 -1584
rect -20193 1584 -20055 2016
rect -20193 -2016 -20055 -1584
rect -19959 1584 -19821 2016
rect -19959 -2016 -19821 -1584
rect -19725 1584 -19587 2016
rect -19725 -2016 -19587 -1584
rect -19491 1584 -19353 2016
rect -19491 -2016 -19353 -1584
rect -19257 1584 -19119 2016
rect -19257 -2016 -19119 -1584
rect -19023 1584 -18885 2016
rect -19023 -2016 -18885 -1584
rect -18789 1584 -18651 2016
rect -18789 -2016 -18651 -1584
rect -18555 1584 -18417 2016
rect -18555 -2016 -18417 -1584
rect -18321 1584 -18183 2016
rect -18321 -2016 -18183 -1584
rect -18087 1584 -17949 2016
rect -18087 -2016 -17949 -1584
rect -17853 1584 -17715 2016
rect -17853 -2016 -17715 -1584
rect -17619 1584 -17481 2016
rect -17619 -2016 -17481 -1584
rect -17385 1584 -17247 2016
rect -17385 -2016 -17247 -1584
rect -17151 1584 -17013 2016
rect -17151 -2016 -17013 -1584
rect -16917 1584 -16779 2016
rect -16917 -2016 -16779 -1584
rect -16683 1584 -16545 2016
rect -16683 -2016 -16545 -1584
rect -16449 1584 -16311 2016
rect -16449 -2016 -16311 -1584
rect -16215 1584 -16077 2016
rect -16215 -2016 -16077 -1584
rect -15981 1584 -15843 2016
rect -15981 -2016 -15843 -1584
rect -15747 1584 -15609 2016
rect -15747 -2016 -15609 -1584
rect -15513 1584 -15375 2016
rect -15513 -2016 -15375 -1584
rect -15279 1584 -15141 2016
rect -15279 -2016 -15141 -1584
rect -15045 1584 -14907 2016
rect -15045 -2016 -14907 -1584
rect -14811 1584 -14673 2016
rect -14811 -2016 -14673 -1584
rect -14577 1584 -14439 2016
rect -14577 -2016 -14439 -1584
rect -14343 1584 -14205 2016
rect -14343 -2016 -14205 -1584
rect -14109 1584 -13971 2016
rect -14109 -2016 -13971 -1584
rect -13875 1584 -13737 2016
rect -13875 -2016 -13737 -1584
rect -13641 1584 -13503 2016
rect -13641 -2016 -13503 -1584
rect -13407 1584 -13269 2016
rect -13407 -2016 -13269 -1584
rect -13173 1584 -13035 2016
rect -13173 -2016 -13035 -1584
rect -12939 1584 -12801 2016
rect -12939 -2016 -12801 -1584
rect -12705 1584 -12567 2016
rect -12705 -2016 -12567 -1584
rect -12471 1584 -12333 2016
rect -12471 -2016 -12333 -1584
rect -12237 1584 -12099 2016
rect -12237 -2016 -12099 -1584
rect -12003 1584 -11865 2016
rect -12003 -2016 -11865 -1584
rect -11769 1584 -11631 2016
rect -11769 -2016 -11631 -1584
rect -11535 1584 -11397 2016
rect -11535 -2016 -11397 -1584
rect -11301 1584 -11163 2016
rect -11301 -2016 -11163 -1584
rect -11067 1584 -10929 2016
rect -11067 -2016 -10929 -1584
rect -10833 1584 -10695 2016
rect -10833 -2016 -10695 -1584
rect -10599 1584 -10461 2016
rect -10599 -2016 -10461 -1584
rect -10365 1584 -10227 2016
rect -10365 -2016 -10227 -1584
rect -10131 1584 -9993 2016
rect -10131 -2016 -9993 -1584
rect -9897 1584 -9759 2016
rect -9897 -2016 -9759 -1584
rect -9663 1584 -9525 2016
rect -9663 -2016 -9525 -1584
rect -9429 1584 -9291 2016
rect -9429 -2016 -9291 -1584
rect -9195 1584 -9057 2016
rect -9195 -2016 -9057 -1584
rect -8961 1584 -8823 2016
rect -8961 -2016 -8823 -1584
rect -8727 1584 -8589 2016
rect -8727 -2016 -8589 -1584
rect -8493 1584 -8355 2016
rect -8493 -2016 -8355 -1584
rect -8259 1584 -8121 2016
rect -8259 -2016 -8121 -1584
rect -8025 1584 -7887 2016
rect -8025 -2016 -7887 -1584
rect -7791 1584 -7653 2016
rect -7791 -2016 -7653 -1584
rect -7557 1584 -7419 2016
rect -7557 -2016 -7419 -1584
rect -7323 1584 -7185 2016
rect -7323 -2016 -7185 -1584
rect -7089 1584 -6951 2016
rect -7089 -2016 -6951 -1584
rect -6855 1584 -6717 2016
rect -6855 -2016 -6717 -1584
rect -6621 1584 -6483 2016
rect -6621 -2016 -6483 -1584
rect -6387 1584 -6249 2016
rect -6387 -2016 -6249 -1584
rect -6153 1584 -6015 2016
rect -6153 -2016 -6015 -1584
rect -5919 1584 -5781 2016
rect -5919 -2016 -5781 -1584
rect -5685 1584 -5547 2016
rect -5685 -2016 -5547 -1584
rect -5451 1584 -5313 2016
rect -5451 -2016 -5313 -1584
rect -5217 1584 -5079 2016
rect -5217 -2016 -5079 -1584
rect -4983 1584 -4845 2016
rect -4983 -2016 -4845 -1584
rect -4749 1584 -4611 2016
rect -4749 -2016 -4611 -1584
rect -4515 1584 -4377 2016
rect -4515 -2016 -4377 -1584
rect -4281 1584 -4143 2016
rect -4281 -2016 -4143 -1584
rect -4047 1584 -3909 2016
rect -4047 -2016 -3909 -1584
rect -3813 1584 -3675 2016
rect -3813 -2016 -3675 -1584
rect -3579 1584 -3441 2016
rect -3579 -2016 -3441 -1584
rect -3345 1584 -3207 2016
rect -3345 -2016 -3207 -1584
rect -3111 1584 -2973 2016
rect -3111 -2016 -2973 -1584
rect -2877 1584 -2739 2016
rect -2877 -2016 -2739 -1584
rect -2643 1584 -2505 2016
rect -2643 -2016 -2505 -1584
rect -2409 1584 -2271 2016
rect -2409 -2016 -2271 -1584
rect -2175 1584 -2037 2016
rect -2175 -2016 -2037 -1584
rect -1941 1584 -1803 2016
rect -1941 -2016 -1803 -1584
rect -1707 1584 -1569 2016
rect -1707 -2016 -1569 -1584
rect -1473 1584 -1335 2016
rect -1473 -2016 -1335 -1584
rect -1239 1584 -1101 2016
rect -1239 -2016 -1101 -1584
rect -1005 1584 -867 2016
rect -1005 -2016 -867 -1584
rect -771 1584 -633 2016
rect -771 -2016 -633 -1584
rect -537 1584 -399 2016
rect -537 -2016 -399 -1584
rect -303 1584 -165 2016
rect -303 -2016 -165 -1584
rect -69 1584 69 2016
rect -69 -2016 69 -1584
rect 165 1584 303 2016
rect 165 -2016 303 -1584
rect 399 1584 537 2016
rect 399 -2016 537 -1584
rect 633 1584 771 2016
rect 633 -2016 771 -1584
rect 867 1584 1005 2016
rect 867 -2016 1005 -1584
rect 1101 1584 1239 2016
rect 1101 -2016 1239 -1584
rect 1335 1584 1473 2016
rect 1335 -2016 1473 -1584
rect 1569 1584 1707 2016
rect 1569 -2016 1707 -1584
rect 1803 1584 1941 2016
rect 1803 -2016 1941 -1584
rect 2037 1584 2175 2016
rect 2037 -2016 2175 -1584
rect 2271 1584 2409 2016
rect 2271 -2016 2409 -1584
rect 2505 1584 2643 2016
rect 2505 -2016 2643 -1584
rect 2739 1584 2877 2016
rect 2739 -2016 2877 -1584
rect 2973 1584 3111 2016
rect 2973 -2016 3111 -1584
rect 3207 1584 3345 2016
rect 3207 -2016 3345 -1584
rect 3441 1584 3579 2016
rect 3441 -2016 3579 -1584
rect 3675 1584 3813 2016
rect 3675 -2016 3813 -1584
rect 3909 1584 4047 2016
rect 3909 -2016 4047 -1584
rect 4143 1584 4281 2016
rect 4143 -2016 4281 -1584
rect 4377 1584 4515 2016
rect 4377 -2016 4515 -1584
rect 4611 1584 4749 2016
rect 4611 -2016 4749 -1584
rect 4845 1584 4983 2016
rect 4845 -2016 4983 -1584
rect 5079 1584 5217 2016
rect 5079 -2016 5217 -1584
rect 5313 1584 5451 2016
rect 5313 -2016 5451 -1584
rect 5547 1584 5685 2016
rect 5547 -2016 5685 -1584
rect 5781 1584 5919 2016
rect 5781 -2016 5919 -1584
rect 6015 1584 6153 2016
rect 6015 -2016 6153 -1584
rect 6249 1584 6387 2016
rect 6249 -2016 6387 -1584
rect 6483 1584 6621 2016
rect 6483 -2016 6621 -1584
rect 6717 1584 6855 2016
rect 6717 -2016 6855 -1584
rect 6951 1584 7089 2016
rect 6951 -2016 7089 -1584
rect 7185 1584 7323 2016
rect 7185 -2016 7323 -1584
rect 7419 1584 7557 2016
rect 7419 -2016 7557 -1584
rect 7653 1584 7791 2016
rect 7653 -2016 7791 -1584
rect 7887 1584 8025 2016
rect 7887 -2016 8025 -1584
rect 8121 1584 8259 2016
rect 8121 -2016 8259 -1584
rect 8355 1584 8493 2016
rect 8355 -2016 8493 -1584
rect 8589 1584 8727 2016
rect 8589 -2016 8727 -1584
rect 8823 1584 8961 2016
rect 8823 -2016 8961 -1584
rect 9057 1584 9195 2016
rect 9057 -2016 9195 -1584
rect 9291 1584 9429 2016
rect 9291 -2016 9429 -1584
rect 9525 1584 9663 2016
rect 9525 -2016 9663 -1584
rect 9759 1584 9897 2016
rect 9759 -2016 9897 -1584
rect 9993 1584 10131 2016
rect 9993 -2016 10131 -1584
rect 10227 1584 10365 2016
rect 10227 -2016 10365 -1584
rect 10461 1584 10599 2016
rect 10461 -2016 10599 -1584
rect 10695 1584 10833 2016
rect 10695 -2016 10833 -1584
rect 10929 1584 11067 2016
rect 10929 -2016 11067 -1584
rect 11163 1584 11301 2016
rect 11163 -2016 11301 -1584
rect 11397 1584 11535 2016
rect 11397 -2016 11535 -1584
rect 11631 1584 11769 2016
rect 11631 -2016 11769 -1584
rect 11865 1584 12003 2016
rect 11865 -2016 12003 -1584
rect 12099 1584 12237 2016
rect 12099 -2016 12237 -1584
rect 12333 1584 12471 2016
rect 12333 -2016 12471 -1584
rect 12567 1584 12705 2016
rect 12567 -2016 12705 -1584
rect 12801 1584 12939 2016
rect 12801 -2016 12939 -1584
rect 13035 1584 13173 2016
rect 13035 -2016 13173 -1584
rect 13269 1584 13407 2016
rect 13269 -2016 13407 -1584
rect 13503 1584 13641 2016
rect 13503 -2016 13641 -1584
rect 13737 1584 13875 2016
rect 13737 -2016 13875 -1584
rect 13971 1584 14109 2016
rect 13971 -2016 14109 -1584
rect 14205 1584 14343 2016
rect 14205 -2016 14343 -1584
rect 14439 1584 14577 2016
rect 14439 -2016 14577 -1584
rect 14673 1584 14811 2016
rect 14673 -2016 14811 -1584
rect 14907 1584 15045 2016
rect 14907 -2016 15045 -1584
rect 15141 1584 15279 2016
rect 15141 -2016 15279 -1584
rect 15375 1584 15513 2016
rect 15375 -2016 15513 -1584
rect 15609 1584 15747 2016
rect 15609 -2016 15747 -1584
rect 15843 1584 15981 2016
rect 15843 -2016 15981 -1584
rect 16077 1584 16215 2016
rect 16077 -2016 16215 -1584
rect 16311 1584 16449 2016
rect 16311 -2016 16449 -1584
rect 16545 1584 16683 2016
rect 16545 -2016 16683 -1584
rect 16779 1584 16917 2016
rect 16779 -2016 16917 -1584
rect 17013 1584 17151 2016
rect 17013 -2016 17151 -1584
rect 17247 1584 17385 2016
rect 17247 -2016 17385 -1584
rect 17481 1584 17619 2016
rect 17481 -2016 17619 -1584
rect 17715 1584 17853 2016
rect 17715 -2016 17853 -1584
rect 17949 1584 18087 2016
rect 17949 -2016 18087 -1584
rect 18183 1584 18321 2016
rect 18183 -2016 18321 -1584
rect 18417 1584 18555 2016
rect 18417 -2016 18555 -1584
rect 18651 1584 18789 2016
rect 18651 -2016 18789 -1584
rect 18885 1584 19023 2016
rect 18885 -2016 19023 -1584
rect 19119 1584 19257 2016
rect 19119 -2016 19257 -1584
rect 19353 1584 19491 2016
rect 19353 -2016 19491 -1584
rect 19587 1584 19725 2016
rect 19587 -2016 19725 -1584
rect 19821 1584 19959 2016
rect 19821 -2016 19959 -1584
rect 20055 1584 20193 2016
rect 20055 -2016 20193 -1584
rect 20289 1584 20427 2016
rect 20289 -2016 20427 -1584
rect 20523 1584 20661 2016
rect 20523 -2016 20661 -1584
rect 20757 1584 20895 2016
rect 20757 -2016 20895 -1584
rect 20991 1584 21129 2016
rect 20991 -2016 21129 -1584
rect 21225 1584 21363 2016
rect 21225 -2016 21363 -1584
rect 21459 1584 21597 2016
rect 21459 -2016 21597 -1584
rect 21693 1584 21831 2016
rect 21693 -2016 21831 -1584
rect 21927 1584 22065 2016
rect 21927 -2016 22065 -1584
rect 22161 1584 22299 2016
rect 22161 -2016 22299 -1584
rect 22395 1584 22533 2016
rect 22395 -2016 22533 -1584
rect 22629 1584 22767 2016
rect 22629 -2016 22767 -1584
rect 22863 1584 23001 2016
rect 22863 -2016 23001 -1584
rect 23097 1584 23235 2016
rect 23097 -2016 23235 -1584
rect 23331 1584 23469 2016
rect 23331 -2016 23469 -1584
<< ppolyres >>
rect -23469 -1584 -23331 1584
rect -23235 -1584 -23097 1584
rect -23001 -1584 -22863 1584
rect -22767 -1584 -22629 1584
rect -22533 -1584 -22395 1584
rect -22299 -1584 -22161 1584
rect -22065 -1584 -21927 1584
rect -21831 -1584 -21693 1584
rect -21597 -1584 -21459 1584
rect -21363 -1584 -21225 1584
rect -21129 -1584 -20991 1584
rect -20895 -1584 -20757 1584
rect -20661 -1584 -20523 1584
rect -20427 -1584 -20289 1584
rect -20193 -1584 -20055 1584
rect -19959 -1584 -19821 1584
rect -19725 -1584 -19587 1584
rect -19491 -1584 -19353 1584
rect -19257 -1584 -19119 1584
rect -19023 -1584 -18885 1584
rect -18789 -1584 -18651 1584
rect -18555 -1584 -18417 1584
rect -18321 -1584 -18183 1584
rect -18087 -1584 -17949 1584
rect -17853 -1584 -17715 1584
rect -17619 -1584 -17481 1584
rect -17385 -1584 -17247 1584
rect -17151 -1584 -17013 1584
rect -16917 -1584 -16779 1584
rect -16683 -1584 -16545 1584
rect -16449 -1584 -16311 1584
rect -16215 -1584 -16077 1584
rect -15981 -1584 -15843 1584
rect -15747 -1584 -15609 1584
rect -15513 -1584 -15375 1584
rect -15279 -1584 -15141 1584
rect -15045 -1584 -14907 1584
rect -14811 -1584 -14673 1584
rect -14577 -1584 -14439 1584
rect -14343 -1584 -14205 1584
rect -14109 -1584 -13971 1584
rect -13875 -1584 -13737 1584
rect -13641 -1584 -13503 1584
rect -13407 -1584 -13269 1584
rect -13173 -1584 -13035 1584
rect -12939 -1584 -12801 1584
rect -12705 -1584 -12567 1584
rect -12471 -1584 -12333 1584
rect -12237 -1584 -12099 1584
rect -12003 -1584 -11865 1584
rect -11769 -1584 -11631 1584
rect -11535 -1584 -11397 1584
rect -11301 -1584 -11163 1584
rect -11067 -1584 -10929 1584
rect -10833 -1584 -10695 1584
rect -10599 -1584 -10461 1584
rect -10365 -1584 -10227 1584
rect -10131 -1584 -9993 1584
rect -9897 -1584 -9759 1584
rect -9663 -1584 -9525 1584
rect -9429 -1584 -9291 1584
rect -9195 -1584 -9057 1584
rect -8961 -1584 -8823 1584
rect -8727 -1584 -8589 1584
rect -8493 -1584 -8355 1584
rect -8259 -1584 -8121 1584
rect -8025 -1584 -7887 1584
rect -7791 -1584 -7653 1584
rect -7557 -1584 -7419 1584
rect -7323 -1584 -7185 1584
rect -7089 -1584 -6951 1584
rect -6855 -1584 -6717 1584
rect -6621 -1584 -6483 1584
rect -6387 -1584 -6249 1584
rect -6153 -1584 -6015 1584
rect -5919 -1584 -5781 1584
rect -5685 -1584 -5547 1584
rect -5451 -1584 -5313 1584
rect -5217 -1584 -5079 1584
rect -4983 -1584 -4845 1584
rect -4749 -1584 -4611 1584
rect -4515 -1584 -4377 1584
rect -4281 -1584 -4143 1584
rect -4047 -1584 -3909 1584
rect -3813 -1584 -3675 1584
rect -3579 -1584 -3441 1584
rect -3345 -1584 -3207 1584
rect -3111 -1584 -2973 1584
rect -2877 -1584 -2739 1584
rect -2643 -1584 -2505 1584
rect -2409 -1584 -2271 1584
rect -2175 -1584 -2037 1584
rect -1941 -1584 -1803 1584
rect -1707 -1584 -1569 1584
rect -1473 -1584 -1335 1584
rect -1239 -1584 -1101 1584
rect -1005 -1584 -867 1584
rect -771 -1584 -633 1584
rect -537 -1584 -399 1584
rect -303 -1584 -165 1584
rect -69 -1584 69 1584
rect 165 -1584 303 1584
rect 399 -1584 537 1584
rect 633 -1584 771 1584
rect 867 -1584 1005 1584
rect 1101 -1584 1239 1584
rect 1335 -1584 1473 1584
rect 1569 -1584 1707 1584
rect 1803 -1584 1941 1584
rect 2037 -1584 2175 1584
rect 2271 -1584 2409 1584
rect 2505 -1584 2643 1584
rect 2739 -1584 2877 1584
rect 2973 -1584 3111 1584
rect 3207 -1584 3345 1584
rect 3441 -1584 3579 1584
rect 3675 -1584 3813 1584
rect 3909 -1584 4047 1584
rect 4143 -1584 4281 1584
rect 4377 -1584 4515 1584
rect 4611 -1584 4749 1584
rect 4845 -1584 4983 1584
rect 5079 -1584 5217 1584
rect 5313 -1584 5451 1584
rect 5547 -1584 5685 1584
rect 5781 -1584 5919 1584
rect 6015 -1584 6153 1584
rect 6249 -1584 6387 1584
rect 6483 -1584 6621 1584
rect 6717 -1584 6855 1584
rect 6951 -1584 7089 1584
rect 7185 -1584 7323 1584
rect 7419 -1584 7557 1584
rect 7653 -1584 7791 1584
rect 7887 -1584 8025 1584
rect 8121 -1584 8259 1584
rect 8355 -1584 8493 1584
rect 8589 -1584 8727 1584
rect 8823 -1584 8961 1584
rect 9057 -1584 9195 1584
rect 9291 -1584 9429 1584
rect 9525 -1584 9663 1584
rect 9759 -1584 9897 1584
rect 9993 -1584 10131 1584
rect 10227 -1584 10365 1584
rect 10461 -1584 10599 1584
rect 10695 -1584 10833 1584
rect 10929 -1584 11067 1584
rect 11163 -1584 11301 1584
rect 11397 -1584 11535 1584
rect 11631 -1584 11769 1584
rect 11865 -1584 12003 1584
rect 12099 -1584 12237 1584
rect 12333 -1584 12471 1584
rect 12567 -1584 12705 1584
rect 12801 -1584 12939 1584
rect 13035 -1584 13173 1584
rect 13269 -1584 13407 1584
rect 13503 -1584 13641 1584
rect 13737 -1584 13875 1584
rect 13971 -1584 14109 1584
rect 14205 -1584 14343 1584
rect 14439 -1584 14577 1584
rect 14673 -1584 14811 1584
rect 14907 -1584 15045 1584
rect 15141 -1584 15279 1584
rect 15375 -1584 15513 1584
rect 15609 -1584 15747 1584
rect 15843 -1584 15981 1584
rect 16077 -1584 16215 1584
rect 16311 -1584 16449 1584
rect 16545 -1584 16683 1584
rect 16779 -1584 16917 1584
rect 17013 -1584 17151 1584
rect 17247 -1584 17385 1584
rect 17481 -1584 17619 1584
rect 17715 -1584 17853 1584
rect 17949 -1584 18087 1584
rect 18183 -1584 18321 1584
rect 18417 -1584 18555 1584
rect 18651 -1584 18789 1584
rect 18885 -1584 19023 1584
rect 19119 -1584 19257 1584
rect 19353 -1584 19491 1584
rect 19587 -1584 19725 1584
rect 19821 -1584 19959 1584
rect 20055 -1584 20193 1584
rect 20289 -1584 20427 1584
rect 20523 -1584 20661 1584
rect 20757 -1584 20895 1584
rect 20991 -1584 21129 1584
rect 21225 -1584 21363 1584
rect 21459 -1584 21597 1584
rect 21693 -1584 21831 1584
rect 21927 -1584 22065 1584
rect 22161 -1584 22299 1584
rect 22395 -1584 22533 1584
rect 22629 -1584 22767 1584
rect 22863 -1584 23001 1584
rect 23097 -1584 23235 1584
rect 23331 -1584 23469 1584
<< locali >>
rect -23599 2112 -23503 2146
rect 23503 2112 23599 2146
rect -23599 2050 -23565 2112
rect 23565 2050 23599 2112
rect -23599 -2112 -23565 -2050
rect 23565 -2112 23599 -2050
rect -23599 -2146 -23503 -2112
rect 23503 -2146 23599 -2112
<< viali >>
rect -23453 1601 -23347 1998
rect -23219 1601 -23113 1998
rect -22985 1601 -22879 1998
rect -22751 1601 -22645 1998
rect -22517 1601 -22411 1998
rect -22283 1601 -22177 1998
rect -22049 1601 -21943 1998
rect -21815 1601 -21709 1998
rect -21581 1601 -21475 1998
rect -21347 1601 -21241 1998
rect -21113 1601 -21007 1998
rect -20879 1601 -20773 1998
rect -20645 1601 -20539 1998
rect -20411 1601 -20305 1998
rect -20177 1601 -20071 1998
rect -19943 1601 -19837 1998
rect -19709 1601 -19603 1998
rect -19475 1601 -19369 1998
rect -19241 1601 -19135 1998
rect -19007 1601 -18901 1998
rect -18773 1601 -18667 1998
rect -18539 1601 -18433 1998
rect -18305 1601 -18199 1998
rect -18071 1601 -17965 1998
rect -17837 1601 -17731 1998
rect -17603 1601 -17497 1998
rect -17369 1601 -17263 1998
rect -17135 1601 -17029 1998
rect -16901 1601 -16795 1998
rect -16667 1601 -16561 1998
rect -16433 1601 -16327 1998
rect -16199 1601 -16093 1998
rect -15965 1601 -15859 1998
rect -15731 1601 -15625 1998
rect -15497 1601 -15391 1998
rect -15263 1601 -15157 1998
rect -15029 1601 -14923 1998
rect -14795 1601 -14689 1998
rect -14561 1601 -14455 1998
rect -14327 1601 -14221 1998
rect -14093 1601 -13987 1998
rect -13859 1601 -13753 1998
rect -13625 1601 -13519 1998
rect -13391 1601 -13285 1998
rect -13157 1601 -13051 1998
rect -12923 1601 -12817 1998
rect -12689 1601 -12583 1998
rect -12455 1601 -12349 1998
rect -12221 1601 -12115 1998
rect -11987 1601 -11881 1998
rect -11753 1601 -11647 1998
rect -11519 1601 -11413 1998
rect -11285 1601 -11179 1998
rect -11051 1601 -10945 1998
rect -10817 1601 -10711 1998
rect -10583 1601 -10477 1998
rect -10349 1601 -10243 1998
rect -10115 1601 -10009 1998
rect -9881 1601 -9775 1998
rect -9647 1601 -9541 1998
rect -9413 1601 -9307 1998
rect -9179 1601 -9073 1998
rect -8945 1601 -8839 1998
rect -8711 1601 -8605 1998
rect -8477 1601 -8371 1998
rect -8243 1601 -8137 1998
rect -8009 1601 -7903 1998
rect -7775 1601 -7669 1998
rect -7541 1601 -7435 1998
rect -7307 1601 -7201 1998
rect -7073 1601 -6967 1998
rect -6839 1601 -6733 1998
rect -6605 1601 -6499 1998
rect -6371 1601 -6265 1998
rect -6137 1601 -6031 1998
rect -5903 1601 -5797 1998
rect -5669 1601 -5563 1998
rect -5435 1601 -5329 1998
rect -5201 1601 -5095 1998
rect -4967 1601 -4861 1998
rect -4733 1601 -4627 1998
rect -4499 1601 -4393 1998
rect -4265 1601 -4159 1998
rect -4031 1601 -3925 1998
rect -3797 1601 -3691 1998
rect -3563 1601 -3457 1998
rect -3329 1601 -3223 1998
rect -3095 1601 -2989 1998
rect -2861 1601 -2755 1998
rect -2627 1601 -2521 1998
rect -2393 1601 -2287 1998
rect -2159 1601 -2053 1998
rect -1925 1601 -1819 1998
rect -1691 1601 -1585 1998
rect -1457 1601 -1351 1998
rect -1223 1601 -1117 1998
rect -989 1601 -883 1998
rect -755 1601 -649 1998
rect -521 1601 -415 1998
rect -287 1601 -181 1998
rect -53 1601 53 1998
rect 181 1601 287 1998
rect 415 1601 521 1998
rect 649 1601 755 1998
rect 883 1601 989 1998
rect 1117 1601 1223 1998
rect 1351 1601 1457 1998
rect 1585 1601 1691 1998
rect 1819 1601 1925 1998
rect 2053 1601 2159 1998
rect 2287 1601 2393 1998
rect 2521 1601 2627 1998
rect 2755 1601 2861 1998
rect 2989 1601 3095 1998
rect 3223 1601 3329 1998
rect 3457 1601 3563 1998
rect 3691 1601 3797 1998
rect 3925 1601 4031 1998
rect 4159 1601 4265 1998
rect 4393 1601 4499 1998
rect 4627 1601 4733 1998
rect 4861 1601 4967 1998
rect 5095 1601 5201 1998
rect 5329 1601 5435 1998
rect 5563 1601 5669 1998
rect 5797 1601 5903 1998
rect 6031 1601 6137 1998
rect 6265 1601 6371 1998
rect 6499 1601 6605 1998
rect 6733 1601 6839 1998
rect 6967 1601 7073 1998
rect 7201 1601 7307 1998
rect 7435 1601 7541 1998
rect 7669 1601 7775 1998
rect 7903 1601 8009 1998
rect 8137 1601 8243 1998
rect 8371 1601 8477 1998
rect 8605 1601 8711 1998
rect 8839 1601 8945 1998
rect 9073 1601 9179 1998
rect 9307 1601 9413 1998
rect 9541 1601 9647 1998
rect 9775 1601 9881 1998
rect 10009 1601 10115 1998
rect 10243 1601 10349 1998
rect 10477 1601 10583 1998
rect 10711 1601 10817 1998
rect 10945 1601 11051 1998
rect 11179 1601 11285 1998
rect 11413 1601 11519 1998
rect 11647 1601 11753 1998
rect 11881 1601 11987 1998
rect 12115 1601 12221 1998
rect 12349 1601 12455 1998
rect 12583 1601 12689 1998
rect 12817 1601 12923 1998
rect 13051 1601 13157 1998
rect 13285 1601 13391 1998
rect 13519 1601 13625 1998
rect 13753 1601 13859 1998
rect 13987 1601 14093 1998
rect 14221 1601 14327 1998
rect 14455 1601 14561 1998
rect 14689 1601 14795 1998
rect 14923 1601 15029 1998
rect 15157 1601 15263 1998
rect 15391 1601 15497 1998
rect 15625 1601 15731 1998
rect 15859 1601 15965 1998
rect 16093 1601 16199 1998
rect 16327 1601 16433 1998
rect 16561 1601 16667 1998
rect 16795 1601 16901 1998
rect 17029 1601 17135 1998
rect 17263 1601 17369 1998
rect 17497 1601 17603 1998
rect 17731 1601 17837 1998
rect 17965 1601 18071 1998
rect 18199 1601 18305 1998
rect 18433 1601 18539 1998
rect 18667 1601 18773 1998
rect 18901 1601 19007 1998
rect 19135 1601 19241 1998
rect 19369 1601 19475 1998
rect 19603 1601 19709 1998
rect 19837 1601 19943 1998
rect 20071 1601 20177 1998
rect 20305 1601 20411 1998
rect 20539 1601 20645 1998
rect 20773 1601 20879 1998
rect 21007 1601 21113 1998
rect 21241 1601 21347 1998
rect 21475 1601 21581 1998
rect 21709 1601 21815 1998
rect 21943 1601 22049 1998
rect 22177 1601 22283 1998
rect 22411 1601 22517 1998
rect 22645 1601 22751 1998
rect 22879 1601 22985 1998
rect 23113 1601 23219 1998
rect 23347 1601 23453 1998
rect -23453 -1998 -23347 -1601
rect -23219 -1998 -23113 -1601
rect -22985 -1998 -22879 -1601
rect -22751 -1998 -22645 -1601
rect -22517 -1998 -22411 -1601
rect -22283 -1998 -22177 -1601
rect -22049 -1998 -21943 -1601
rect -21815 -1998 -21709 -1601
rect -21581 -1998 -21475 -1601
rect -21347 -1998 -21241 -1601
rect -21113 -1998 -21007 -1601
rect -20879 -1998 -20773 -1601
rect -20645 -1998 -20539 -1601
rect -20411 -1998 -20305 -1601
rect -20177 -1998 -20071 -1601
rect -19943 -1998 -19837 -1601
rect -19709 -1998 -19603 -1601
rect -19475 -1998 -19369 -1601
rect -19241 -1998 -19135 -1601
rect -19007 -1998 -18901 -1601
rect -18773 -1998 -18667 -1601
rect -18539 -1998 -18433 -1601
rect -18305 -1998 -18199 -1601
rect -18071 -1998 -17965 -1601
rect -17837 -1998 -17731 -1601
rect -17603 -1998 -17497 -1601
rect -17369 -1998 -17263 -1601
rect -17135 -1998 -17029 -1601
rect -16901 -1998 -16795 -1601
rect -16667 -1998 -16561 -1601
rect -16433 -1998 -16327 -1601
rect -16199 -1998 -16093 -1601
rect -15965 -1998 -15859 -1601
rect -15731 -1998 -15625 -1601
rect -15497 -1998 -15391 -1601
rect -15263 -1998 -15157 -1601
rect -15029 -1998 -14923 -1601
rect -14795 -1998 -14689 -1601
rect -14561 -1998 -14455 -1601
rect -14327 -1998 -14221 -1601
rect -14093 -1998 -13987 -1601
rect -13859 -1998 -13753 -1601
rect -13625 -1998 -13519 -1601
rect -13391 -1998 -13285 -1601
rect -13157 -1998 -13051 -1601
rect -12923 -1998 -12817 -1601
rect -12689 -1998 -12583 -1601
rect -12455 -1998 -12349 -1601
rect -12221 -1998 -12115 -1601
rect -11987 -1998 -11881 -1601
rect -11753 -1998 -11647 -1601
rect -11519 -1998 -11413 -1601
rect -11285 -1998 -11179 -1601
rect -11051 -1998 -10945 -1601
rect -10817 -1998 -10711 -1601
rect -10583 -1998 -10477 -1601
rect -10349 -1998 -10243 -1601
rect -10115 -1998 -10009 -1601
rect -9881 -1998 -9775 -1601
rect -9647 -1998 -9541 -1601
rect -9413 -1998 -9307 -1601
rect -9179 -1998 -9073 -1601
rect -8945 -1998 -8839 -1601
rect -8711 -1998 -8605 -1601
rect -8477 -1998 -8371 -1601
rect -8243 -1998 -8137 -1601
rect -8009 -1998 -7903 -1601
rect -7775 -1998 -7669 -1601
rect -7541 -1998 -7435 -1601
rect -7307 -1998 -7201 -1601
rect -7073 -1998 -6967 -1601
rect -6839 -1998 -6733 -1601
rect -6605 -1998 -6499 -1601
rect -6371 -1998 -6265 -1601
rect -6137 -1998 -6031 -1601
rect -5903 -1998 -5797 -1601
rect -5669 -1998 -5563 -1601
rect -5435 -1998 -5329 -1601
rect -5201 -1998 -5095 -1601
rect -4967 -1998 -4861 -1601
rect -4733 -1998 -4627 -1601
rect -4499 -1998 -4393 -1601
rect -4265 -1998 -4159 -1601
rect -4031 -1998 -3925 -1601
rect -3797 -1998 -3691 -1601
rect -3563 -1998 -3457 -1601
rect -3329 -1998 -3223 -1601
rect -3095 -1998 -2989 -1601
rect -2861 -1998 -2755 -1601
rect -2627 -1998 -2521 -1601
rect -2393 -1998 -2287 -1601
rect -2159 -1998 -2053 -1601
rect -1925 -1998 -1819 -1601
rect -1691 -1998 -1585 -1601
rect -1457 -1998 -1351 -1601
rect -1223 -1998 -1117 -1601
rect -989 -1998 -883 -1601
rect -755 -1998 -649 -1601
rect -521 -1998 -415 -1601
rect -287 -1998 -181 -1601
rect -53 -1998 53 -1601
rect 181 -1998 287 -1601
rect 415 -1998 521 -1601
rect 649 -1998 755 -1601
rect 883 -1998 989 -1601
rect 1117 -1998 1223 -1601
rect 1351 -1998 1457 -1601
rect 1585 -1998 1691 -1601
rect 1819 -1998 1925 -1601
rect 2053 -1998 2159 -1601
rect 2287 -1998 2393 -1601
rect 2521 -1998 2627 -1601
rect 2755 -1998 2861 -1601
rect 2989 -1998 3095 -1601
rect 3223 -1998 3329 -1601
rect 3457 -1998 3563 -1601
rect 3691 -1998 3797 -1601
rect 3925 -1998 4031 -1601
rect 4159 -1998 4265 -1601
rect 4393 -1998 4499 -1601
rect 4627 -1998 4733 -1601
rect 4861 -1998 4967 -1601
rect 5095 -1998 5201 -1601
rect 5329 -1998 5435 -1601
rect 5563 -1998 5669 -1601
rect 5797 -1998 5903 -1601
rect 6031 -1998 6137 -1601
rect 6265 -1998 6371 -1601
rect 6499 -1998 6605 -1601
rect 6733 -1998 6839 -1601
rect 6967 -1998 7073 -1601
rect 7201 -1998 7307 -1601
rect 7435 -1998 7541 -1601
rect 7669 -1998 7775 -1601
rect 7903 -1998 8009 -1601
rect 8137 -1998 8243 -1601
rect 8371 -1998 8477 -1601
rect 8605 -1998 8711 -1601
rect 8839 -1998 8945 -1601
rect 9073 -1998 9179 -1601
rect 9307 -1998 9413 -1601
rect 9541 -1998 9647 -1601
rect 9775 -1998 9881 -1601
rect 10009 -1998 10115 -1601
rect 10243 -1998 10349 -1601
rect 10477 -1998 10583 -1601
rect 10711 -1998 10817 -1601
rect 10945 -1998 11051 -1601
rect 11179 -1998 11285 -1601
rect 11413 -1998 11519 -1601
rect 11647 -1998 11753 -1601
rect 11881 -1998 11987 -1601
rect 12115 -1998 12221 -1601
rect 12349 -1998 12455 -1601
rect 12583 -1998 12689 -1601
rect 12817 -1998 12923 -1601
rect 13051 -1998 13157 -1601
rect 13285 -1998 13391 -1601
rect 13519 -1998 13625 -1601
rect 13753 -1998 13859 -1601
rect 13987 -1998 14093 -1601
rect 14221 -1998 14327 -1601
rect 14455 -1998 14561 -1601
rect 14689 -1998 14795 -1601
rect 14923 -1998 15029 -1601
rect 15157 -1998 15263 -1601
rect 15391 -1998 15497 -1601
rect 15625 -1998 15731 -1601
rect 15859 -1998 15965 -1601
rect 16093 -1998 16199 -1601
rect 16327 -1998 16433 -1601
rect 16561 -1998 16667 -1601
rect 16795 -1998 16901 -1601
rect 17029 -1998 17135 -1601
rect 17263 -1998 17369 -1601
rect 17497 -1998 17603 -1601
rect 17731 -1998 17837 -1601
rect 17965 -1998 18071 -1601
rect 18199 -1998 18305 -1601
rect 18433 -1998 18539 -1601
rect 18667 -1998 18773 -1601
rect 18901 -1998 19007 -1601
rect 19135 -1998 19241 -1601
rect 19369 -1998 19475 -1601
rect 19603 -1998 19709 -1601
rect 19837 -1998 19943 -1601
rect 20071 -1998 20177 -1601
rect 20305 -1998 20411 -1601
rect 20539 -1998 20645 -1601
rect 20773 -1998 20879 -1601
rect 21007 -1998 21113 -1601
rect 21241 -1998 21347 -1601
rect 21475 -1998 21581 -1601
rect 21709 -1998 21815 -1601
rect 21943 -1998 22049 -1601
rect 22177 -1998 22283 -1601
rect 22411 -1998 22517 -1601
rect 22645 -1998 22751 -1601
rect 22879 -1998 22985 -1601
rect 23113 -1998 23219 -1601
rect 23347 -1998 23453 -1601
<< metal1 >>
rect -23459 1998 -23341 2010
rect -23459 1601 -23453 1998
rect -23347 1601 -23341 1998
rect -23459 1589 -23341 1601
rect -23225 1998 -23107 2010
rect -23225 1601 -23219 1998
rect -23113 1601 -23107 1998
rect -23225 1589 -23107 1601
rect -22991 1998 -22873 2010
rect -22991 1601 -22985 1998
rect -22879 1601 -22873 1998
rect -22991 1589 -22873 1601
rect -22757 1998 -22639 2010
rect -22757 1601 -22751 1998
rect -22645 1601 -22639 1998
rect -22757 1589 -22639 1601
rect -22523 1998 -22405 2010
rect -22523 1601 -22517 1998
rect -22411 1601 -22405 1998
rect -22523 1589 -22405 1601
rect -22289 1998 -22171 2010
rect -22289 1601 -22283 1998
rect -22177 1601 -22171 1998
rect -22289 1589 -22171 1601
rect -22055 1998 -21937 2010
rect -22055 1601 -22049 1998
rect -21943 1601 -21937 1998
rect -22055 1589 -21937 1601
rect -21821 1998 -21703 2010
rect -21821 1601 -21815 1998
rect -21709 1601 -21703 1998
rect -21821 1589 -21703 1601
rect -21587 1998 -21469 2010
rect -21587 1601 -21581 1998
rect -21475 1601 -21469 1998
rect -21587 1589 -21469 1601
rect -21353 1998 -21235 2010
rect -21353 1601 -21347 1998
rect -21241 1601 -21235 1998
rect -21353 1589 -21235 1601
rect -21119 1998 -21001 2010
rect -21119 1601 -21113 1998
rect -21007 1601 -21001 1998
rect -21119 1589 -21001 1601
rect -20885 1998 -20767 2010
rect -20885 1601 -20879 1998
rect -20773 1601 -20767 1998
rect -20885 1589 -20767 1601
rect -20651 1998 -20533 2010
rect -20651 1601 -20645 1998
rect -20539 1601 -20533 1998
rect -20651 1589 -20533 1601
rect -20417 1998 -20299 2010
rect -20417 1601 -20411 1998
rect -20305 1601 -20299 1998
rect -20417 1589 -20299 1601
rect -20183 1998 -20065 2010
rect -20183 1601 -20177 1998
rect -20071 1601 -20065 1998
rect -20183 1589 -20065 1601
rect -19949 1998 -19831 2010
rect -19949 1601 -19943 1998
rect -19837 1601 -19831 1998
rect -19949 1589 -19831 1601
rect -19715 1998 -19597 2010
rect -19715 1601 -19709 1998
rect -19603 1601 -19597 1998
rect -19715 1589 -19597 1601
rect -19481 1998 -19363 2010
rect -19481 1601 -19475 1998
rect -19369 1601 -19363 1998
rect -19481 1589 -19363 1601
rect -19247 1998 -19129 2010
rect -19247 1601 -19241 1998
rect -19135 1601 -19129 1998
rect -19247 1589 -19129 1601
rect -19013 1998 -18895 2010
rect -19013 1601 -19007 1998
rect -18901 1601 -18895 1998
rect -19013 1589 -18895 1601
rect -18779 1998 -18661 2010
rect -18779 1601 -18773 1998
rect -18667 1601 -18661 1998
rect -18779 1589 -18661 1601
rect -18545 1998 -18427 2010
rect -18545 1601 -18539 1998
rect -18433 1601 -18427 1998
rect -18545 1589 -18427 1601
rect -18311 1998 -18193 2010
rect -18311 1601 -18305 1998
rect -18199 1601 -18193 1998
rect -18311 1589 -18193 1601
rect -18077 1998 -17959 2010
rect -18077 1601 -18071 1998
rect -17965 1601 -17959 1998
rect -18077 1589 -17959 1601
rect -17843 1998 -17725 2010
rect -17843 1601 -17837 1998
rect -17731 1601 -17725 1998
rect -17843 1589 -17725 1601
rect -17609 1998 -17491 2010
rect -17609 1601 -17603 1998
rect -17497 1601 -17491 1998
rect -17609 1589 -17491 1601
rect -17375 1998 -17257 2010
rect -17375 1601 -17369 1998
rect -17263 1601 -17257 1998
rect -17375 1589 -17257 1601
rect -17141 1998 -17023 2010
rect -17141 1601 -17135 1998
rect -17029 1601 -17023 1998
rect -17141 1589 -17023 1601
rect -16907 1998 -16789 2010
rect -16907 1601 -16901 1998
rect -16795 1601 -16789 1998
rect -16907 1589 -16789 1601
rect -16673 1998 -16555 2010
rect -16673 1601 -16667 1998
rect -16561 1601 -16555 1998
rect -16673 1589 -16555 1601
rect -16439 1998 -16321 2010
rect -16439 1601 -16433 1998
rect -16327 1601 -16321 1998
rect -16439 1589 -16321 1601
rect -16205 1998 -16087 2010
rect -16205 1601 -16199 1998
rect -16093 1601 -16087 1998
rect -16205 1589 -16087 1601
rect -15971 1998 -15853 2010
rect -15971 1601 -15965 1998
rect -15859 1601 -15853 1998
rect -15971 1589 -15853 1601
rect -15737 1998 -15619 2010
rect -15737 1601 -15731 1998
rect -15625 1601 -15619 1998
rect -15737 1589 -15619 1601
rect -15503 1998 -15385 2010
rect -15503 1601 -15497 1998
rect -15391 1601 -15385 1998
rect -15503 1589 -15385 1601
rect -15269 1998 -15151 2010
rect -15269 1601 -15263 1998
rect -15157 1601 -15151 1998
rect -15269 1589 -15151 1601
rect -15035 1998 -14917 2010
rect -15035 1601 -15029 1998
rect -14923 1601 -14917 1998
rect -15035 1589 -14917 1601
rect -14801 1998 -14683 2010
rect -14801 1601 -14795 1998
rect -14689 1601 -14683 1998
rect -14801 1589 -14683 1601
rect -14567 1998 -14449 2010
rect -14567 1601 -14561 1998
rect -14455 1601 -14449 1998
rect -14567 1589 -14449 1601
rect -14333 1998 -14215 2010
rect -14333 1601 -14327 1998
rect -14221 1601 -14215 1998
rect -14333 1589 -14215 1601
rect -14099 1998 -13981 2010
rect -14099 1601 -14093 1998
rect -13987 1601 -13981 1998
rect -14099 1589 -13981 1601
rect -13865 1998 -13747 2010
rect -13865 1601 -13859 1998
rect -13753 1601 -13747 1998
rect -13865 1589 -13747 1601
rect -13631 1998 -13513 2010
rect -13631 1601 -13625 1998
rect -13519 1601 -13513 1998
rect -13631 1589 -13513 1601
rect -13397 1998 -13279 2010
rect -13397 1601 -13391 1998
rect -13285 1601 -13279 1998
rect -13397 1589 -13279 1601
rect -13163 1998 -13045 2010
rect -13163 1601 -13157 1998
rect -13051 1601 -13045 1998
rect -13163 1589 -13045 1601
rect -12929 1998 -12811 2010
rect -12929 1601 -12923 1998
rect -12817 1601 -12811 1998
rect -12929 1589 -12811 1601
rect -12695 1998 -12577 2010
rect -12695 1601 -12689 1998
rect -12583 1601 -12577 1998
rect -12695 1589 -12577 1601
rect -12461 1998 -12343 2010
rect -12461 1601 -12455 1998
rect -12349 1601 -12343 1998
rect -12461 1589 -12343 1601
rect -12227 1998 -12109 2010
rect -12227 1601 -12221 1998
rect -12115 1601 -12109 1998
rect -12227 1589 -12109 1601
rect -11993 1998 -11875 2010
rect -11993 1601 -11987 1998
rect -11881 1601 -11875 1998
rect -11993 1589 -11875 1601
rect -11759 1998 -11641 2010
rect -11759 1601 -11753 1998
rect -11647 1601 -11641 1998
rect -11759 1589 -11641 1601
rect -11525 1998 -11407 2010
rect -11525 1601 -11519 1998
rect -11413 1601 -11407 1998
rect -11525 1589 -11407 1601
rect -11291 1998 -11173 2010
rect -11291 1601 -11285 1998
rect -11179 1601 -11173 1998
rect -11291 1589 -11173 1601
rect -11057 1998 -10939 2010
rect -11057 1601 -11051 1998
rect -10945 1601 -10939 1998
rect -11057 1589 -10939 1601
rect -10823 1998 -10705 2010
rect -10823 1601 -10817 1998
rect -10711 1601 -10705 1998
rect -10823 1589 -10705 1601
rect -10589 1998 -10471 2010
rect -10589 1601 -10583 1998
rect -10477 1601 -10471 1998
rect -10589 1589 -10471 1601
rect -10355 1998 -10237 2010
rect -10355 1601 -10349 1998
rect -10243 1601 -10237 1998
rect -10355 1589 -10237 1601
rect -10121 1998 -10003 2010
rect -10121 1601 -10115 1998
rect -10009 1601 -10003 1998
rect -10121 1589 -10003 1601
rect -9887 1998 -9769 2010
rect -9887 1601 -9881 1998
rect -9775 1601 -9769 1998
rect -9887 1589 -9769 1601
rect -9653 1998 -9535 2010
rect -9653 1601 -9647 1998
rect -9541 1601 -9535 1998
rect -9653 1589 -9535 1601
rect -9419 1998 -9301 2010
rect -9419 1601 -9413 1998
rect -9307 1601 -9301 1998
rect -9419 1589 -9301 1601
rect -9185 1998 -9067 2010
rect -9185 1601 -9179 1998
rect -9073 1601 -9067 1998
rect -9185 1589 -9067 1601
rect -8951 1998 -8833 2010
rect -8951 1601 -8945 1998
rect -8839 1601 -8833 1998
rect -8951 1589 -8833 1601
rect -8717 1998 -8599 2010
rect -8717 1601 -8711 1998
rect -8605 1601 -8599 1998
rect -8717 1589 -8599 1601
rect -8483 1998 -8365 2010
rect -8483 1601 -8477 1998
rect -8371 1601 -8365 1998
rect -8483 1589 -8365 1601
rect -8249 1998 -8131 2010
rect -8249 1601 -8243 1998
rect -8137 1601 -8131 1998
rect -8249 1589 -8131 1601
rect -8015 1998 -7897 2010
rect -8015 1601 -8009 1998
rect -7903 1601 -7897 1998
rect -8015 1589 -7897 1601
rect -7781 1998 -7663 2010
rect -7781 1601 -7775 1998
rect -7669 1601 -7663 1998
rect -7781 1589 -7663 1601
rect -7547 1998 -7429 2010
rect -7547 1601 -7541 1998
rect -7435 1601 -7429 1998
rect -7547 1589 -7429 1601
rect -7313 1998 -7195 2010
rect -7313 1601 -7307 1998
rect -7201 1601 -7195 1998
rect -7313 1589 -7195 1601
rect -7079 1998 -6961 2010
rect -7079 1601 -7073 1998
rect -6967 1601 -6961 1998
rect -7079 1589 -6961 1601
rect -6845 1998 -6727 2010
rect -6845 1601 -6839 1998
rect -6733 1601 -6727 1998
rect -6845 1589 -6727 1601
rect -6611 1998 -6493 2010
rect -6611 1601 -6605 1998
rect -6499 1601 -6493 1998
rect -6611 1589 -6493 1601
rect -6377 1998 -6259 2010
rect -6377 1601 -6371 1998
rect -6265 1601 -6259 1998
rect -6377 1589 -6259 1601
rect -6143 1998 -6025 2010
rect -6143 1601 -6137 1998
rect -6031 1601 -6025 1998
rect -6143 1589 -6025 1601
rect -5909 1998 -5791 2010
rect -5909 1601 -5903 1998
rect -5797 1601 -5791 1998
rect -5909 1589 -5791 1601
rect -5675 1998 -5557 2010
rect -5675 1601 -5669 1998
rect -5563 1601 -5557 1998
rect -5675 1589 -5557 1601
rect -5441 1998 -5323 2010
rect -5441 1601 -5435 1998
rect -5329 1601 -5323 1998
rect -5441 1589 -5323 1601
rect -5207 1998 -5089 2010
rect -5207 1601 -5201 1998
rect -5095 1601 -5089 1998
rect -5207 1589 -5089 1601
rect -4973 1998 -4855 2010
rect -4973 1601 -4967 1998
rect -4861 1601 -4855 1998
rect -4973 1589 -4855 1601
rect -4739 1998 -4621 2010
rect -4739 1601 -4733 1998
rect -4627 1601 -4621 1998
rect -4739 1589 -4621 1601
rect -4505 1998 -4387 2010
rect -4505 1601 -4499 1998
rect -4393 1601 -4387 1998
rect -4505 1589 -4387 1601
rect -4271 1998 -4153 2010
rect -4271 1601 -4265 1998
rect -4159 1601 -4153 1998
rect -4271 1589 -4153 1601
rect -4037 1998 -3919 2010
rect -4037 1601 -4031 1998
rect -3925 1601 -3919 1998
rect -4037 1589 -3919 1601
rect -3803 1998 -3685 2010
rect -3803 1601 -3797 1998
rect -3691 1601 -3685 1998
rect -3803 1589 -3685 1601
rect -3569 1998 -3451 2010
rect -3569 1601 -3563 1998
rect -3457 1601 -3451 1998
rect -3569 1589 -3451 1601
rect -3335 1998 -3217 2010
rect -3335 1601 -3329 1998
rect -3223 1601 -3217 1998
rect -3335 1589 -3217 1601
rect -3101 1998 -2983 2010
rect -3101 1601 -3095 1998
rect -2989 1601 -2983 1998
rect -3101 1589 -2983 1601
rect -2867 1998 -2749 2010
rect -2867 1601 -2861 1998
rect -2755 1601 -2749 1998
rect -2867 1589 -2749 1601
rect -2633 1998 -2515 2010
rect -2633 1601 -2627 1998
rect -2521 1601 -2515 1998
rect -2633 1589 -2515 1601
rect -2399 1998 -2281 2010
rect -2399 1601 -2393 1998
rect -2287 1601 -2281 1998
rect -2399 1589 -2281 1601
rect -2165 1998 -2047 2010
rect -2165 1601 -2159 1998
rect -2053 1601 -2047 1998
rect -2165 1589 -2047 1601
rect -1931 1998 -1813 2010
rect -1931 1601 -1925 1998
rect -1819 1601 -1813 1998
rect -1931 1589 -1813 1601
rect -1697 1998 -1579 2010
rect -1697 1601 -1691 1998
rect -1585 1601 -1579 1998
rect -1697 1589 -1579 1601
rect -1463 1998 -1345 2010
rect -1463 1601 -1457 1998
rect -1351 1601 -1345 1998
rect -1463 1589 -1345 1601
rect -1229 1998 -1111 2010
rect -1229 1601 -1223 1998
rect -1117 1601 -1111 1998
rect -1229 1589 -1111 1601
rect -995 1998 -877 2010
rect -995 1601 -989 1998
rect -883 1601 -877 1998
rect -995 1589 -877 1601
rect -761 1998 -643 2010
rect -761 1601 -755 1998
rect -649 1601 -643 1998
rect -761 1589 -643 1601
rect -527 1998 -409 2010
rect -527 1601 -521 1998
rect -415 1601 -409 1998
rect -527 1589 -409 1601
rect -293 1998 -175 2010
rect -293 1601 -287 1998
rect -181 1601 -175 1998
rect -293 1589 -175 1601
rect -59 1998 59 2010
rect -59 1601 -53 1998
rect 53 1601 59 1998
rect -59 1589 59 1601
rect 175 1998 293 2010
rect 175 1601 181 1998
rect 287 1601 293 1998
rect 175 1589 293 1601
rect 409 1998 527 2010
rect 409 1601 415 1998
rect 521 1601 527 1998
rect 409 1589 527 1601
rect 643 1998 761 2010
rect 643 1601 649 1998
rect 755 1601 761 1998
rect 643 1589 761 1601
rect 877 1998 995 2010
rect 877 1601 883 1998
rect 989 1601 995 1998
rect 877 1589 995 1601
rect 1111 1998 1229 2010
rect 1111 1601 1117 1998
rect 1223 1601 1229 1998
rect 1111 1589 1229 1601
rect 1345 1998 1463 2010
rect 1345 1601 1351 1998
rect 1457 1601 1463 1998
rect 1345 1589 1463 1601
rect 1579 1998 1697 2010
rect 1579 1601 1585 1998
rect 1691 1601 1697 1998
rect 1579 1589 1697 1601
rect 1813 1998 1931 2010
rect 1813 1601 1819 1998
rect 1925 1601 1931 1998
rect 1813 1589 1931 1601
rect 2047 1998 2165 2010
rect 2047 1601 2053 1998
rect 2159 1601 2165 1998
rect 2047 1589 2165 1601
rect 2281 1998 2399 2010
rect 2281 1601 2287 1998
rect 2393 1601 2399 1998
rect 2281 1589 2399 1601
rect 2515 1998 2633 2010
rect 2515 1601 2521 1998
rect 2627 1601 2633 1998
rect 2515 1589 2633 1601
rect 2749 1998 2867 2010
rect 2749 1601 2755 1998
rect 2861 1601 2867 1998
rect 2749 1589 2867 1601
rect 2983 1998 3101 2010
rect 2983 1601 2989 1998
rect 3095 1601 3101 1998
rect 2983 1589 3101 1601
rect 3217 1998 3335 2010
rect 3217 1601 3223 1998
rect 3329 1601 3335 1998
rect 3217 1589 3335 1601
rect 3451 1998 3569 2010
rect 3451 1601 3457 1998
rect 3563 1601 3569 1998
rect 3451 1589 3569 1601
rect 3685 1998 3803 2010
rect 3685 1601 3691 1998
rect 3797 1601 3803 1998
rect 3685 1589 3803 1601
rect 3919 1998 4037 2010
rect 3919 1601 3925 1998
rect 4031 1601 4037 1998
rect 3919 1589 4037 1601
rect 4153 1998 4271 2010
rect 4153 1601 4159 1998
rect 4265 1601 4271 1998
rect 4153 1589 4271 1601
rect 4387 1998 4505 2010
rect 4387 1601 4393 1998
rect 4499 1601 4505 1998
rect 4387 1589 4505 1601
rect 4621 1998 4739 2010
rect 4621 1601 4627 1998
rect 4733 1601 4739 1998
rect 4621 1589 4739 1601
rect 4855 1998 4973 2010
rect 4855 1601 4861 1998
rect 4967 1601 4973 1998
rect 4855 1589 4973 1601
rect 5089 1998 5207 2010
rect 5089 1601 5095 1998
rect 5201 1601 5207 1998
rect 5089 1589 5207 1601
rect 5323 1998 5441 2010
rect 5323 1601 5329 1998
rect 5435 1601 5441 1998
rect 5323 1589 5441 1601
rect 5557 1998 5675 2010
rect 5557 1601 5563 1998
rect 5669 1601 5675 1998
rect 5557 1589 5675 1601
rect 5791 1998 5909 2010
rect 5791 1601 5797 1998
rect 5903 1601 5909 1998
rect 5791 1589 5909 1601
rect 6025 1998 6143 2010
rect 6025 1601 6031 1998
rect 6137 1601 6143 1998
rect 6025 1589 6143 1601
rect 6259 1998 6377 2010
rect 6259 1601 6265 1998
rect 6371 1601 6377 1998
rect 6259 1589 6377 1601
rect 6493 1998 6611 2010
rect 6493 1601 6499 1998
rect 6605 1601 6611 1998
rect 6493 1589 6611 1601
rect 6727 1998 6845 2010
rect 6727 1601 6733 1998
rect 6839 1601 6845 1998
rect 6727 1589 6845 1601
rect 6961 1998 7079 2010
rect 6961 1601 6967 1998
rect 7073 1601 7079 1998
rect 6961 1589 7079 1601
rect 7195 1998 7313 2010
rect 7195 1601 7201 1998
rect 7307 1601 7313 1998
rect 7195 1589 7313 1601
rect 7429 1998 7547 2010
rect 7429 1601 7435 1998
rect 7541 1601 7547 1998
rect 7429 1589 7547 1601
rect 7663 1998 7781 2010
rect 7663 1601 7669 1998
rect 7775 1601 7781 1998
rect 7663 1589 7781 1601
rect 7897 1998 8015 2010
rect 7897 1601 7903 1998
rect 8009 1601 8015 1998
rect 7897 1589 8015 1601
rect 8131 1998 8249 2010
rect 8131 1601 8137 1998
rect 8243 1601 8249 1998
rect 8131 1589 8249 1601
rect 8365 1998 8483 2010
rect 8365 1601 8371 1998
rect 8477 1601 8483 1998
rect 8365 1589 8483 1601
rect 8599 1998 8717 2010
rect 8599 1601 8605 1998
rect 8711 1601 8717 1998
rect 8599 1589 8717 1601
rect 8833 1998 8951 2010
rect 8833 1601 8839 1998
rect 8945 1601 8951 1998
rect 8833 1589 8951 1601
rect 9067 1998 9185 2010
rect 9067 1601 9073 1998
rect 9179 1601 9185 1998
rect 9067 1589 9185 1601
rect 9301 1998 9419 2010
rect 9301 1601 9307 1998
rect 9413 1601 9419 1998
rect 9301 1589 9419 1601
rect 9535 1998 9653 2010
rect 9535 1601 9541 1998
rect 9647 1601 9653 1998
rect 9535 1589 9653 1601
rect 9769 1998 9887 2010
rect 9769 1601 9775 1998
rect 9881 1601 9887 1998
rect 9769 1589 9887 1601
rect 10003 1998 10121 2010
rect 10003 1601 10009 1998
rect 10115 1601 10121 1998
rect 10003 1589 10121 1601
rect 10237 1998 10355 2010
rect 10237 1601 10243 1998
rect 10349 1601 10355 1998
rect 10237 1589 10355 1601
rect 10471 1998 10589 2010
rect 10471 1601 10477 1998
rect 10583 1601 10589 1998
rect 10471 1589 10589 1601
rect 10705 1998 10823 2010
rect 10705 1601 10711 1998
rect 10817 1601 10823 1998
rect 10705 1589 10823 1601
rect 10939 1998 11057 2010
rect 10939 1601 10945 1998
rect 11051 1601 11057 1998
rect 10939 1589 11057 1601
rect 11173 1998 11291 2010
rect 11173 1601 11179 1998
rect 11285 1601 11291 1998
rect 11173 1589 11291 1601
rect 11407 1998 11525 2010
rect 11407 1601 11413 1998
rect 11519 1601 11525 1998
rect 11407 1589 11525 1601
rect 11641 1998 11759 2010
rect 11641 1601 11647 1998
rect 11753 1601 11759 1998
rect 11641 1589 11759 1601
rect 11875 1998 11993 2010
rect 11875 1601 11881 1998
rect 11987 1601 11993 1998
rect 11875 1589 11993 1601
rect 12109 1998 12227 2010
rect 12109 1601 12115 1998
rect 12221 1601 12227 1998
rect 12109 1589 12227 1601
rect 12343 1998 12461 2010
rect 12343 1601 12349 1998
rect 12455 1601 12461 1998
rect 12343 1589 12461 1601
rect 12577 1998 12695 2010
rect 12577 1601 12583 1998
rect 12689 1601 12695 1998
rect 12577 1589 12695 1601
rect 12811 1998 12929 2010
rect 12811 1601 12817 1998
rect 12923 1601 12929 1998
rect 12811 1589 12929 1601
rect 13045 1998 13163 2010
rect 13045 1601 13051 1998
rect 13157 1601 13163 1998
rect 13045 1589 13163 1601
rect 13279 1998 13397 2010
rect 13279 1601 13285 1998
rect 13391 1601 13397 1998
rect 13279 1589 13397 1601
rect 13513 1998 13631 2010
rect 13513 1601 13519 1998
rect 13625 1601 13631 1998
rect 13513 1589 13631 1601
rect 13747 1998 13865 2010
rect 13747 1601 13753 1998
rect 13859 1601 13865 1998
rect 13747 1589 13865 1601
rect 13981 1998 14099 2010
rect 13981 1601 13987 1998
rect 14093 1601 14099 1998
rect 13981 1589 14099 1601
rect 14215 1998 14333 2010
rect 14215 1601 14221 1998
rect 14327 1601 14333 1998
rect 14215 1589 14333 1601
rect 14449 1998 14567 2010
rect 14449 1601 14455 1998
rect 14561 1601 14567 1998
rect 14449 1589 14567 1601
rect 14683 1998 14801 2010
rect 14683 1601 14689 1998
rect 14795 1601 14801 1998
rect 14683 1589 14801 1601
rect 14917 1998 15035 2010
rect 14917 1601 14923 1998
rect 15029 1601 15035 1998
rect 14917 1589 15035 1601
rect 15151 1998 15269 2010
rect 15151 1601 15157 1998
rect 15263 1601 15269 1998
rect 15151 1589 15269 1601
rect 15385 1998 15503 2010
rect 15385 1601 15391 1998
rect 15497 1601 15503 1998
rect 15385 1589 15503 1601
rect 15619 1998 15737 2010
rect 15619 1601 15625 1998
rect 15731 1601 15737 1998
rect 15619 1589 15737 1601
rect 15853 1998 15971 2010
rect 15853 1601 15859 1998
rect 15965 1601 15971 1998
rect 15853 1589 15971 1601
rect 16087 1998 16205 2010
rect 16087 1601 16093 1998
rect 16199 1601 16205 1998
rect 16087 1589 16205 1601
rect 16321 1998 16439 2010
rect 16321 1601 16327 1998
rect 16433 1601 16439 1998
rect 16321 1589 16439 1601
rect 16555 1998 16673 2010
rect 16555 1601 16561 1998
rect 16667 1601 16673 1998
rect 16555 1589 16673 1601
rect 16789 1998 16907 2010
rect 16789 1601 16795 1998
rect 16901 1601 16907 1998
rect 16789 1589 16907 1601
rect 17023 1998 17141 2010
rect 17023 1601 17029 1998
rect 17135 1601 17141 1998
rect 17023 1589 17141 1601
rect 17257 1998 17375 2010
rect 17257 1601 17263 1998
rect 17369 1601 17375 1998
rect 17257 1589 17375 1601
rect 17491 1998 17609 2010
rect 17491 1601 17497 1998
rect 17603 1601 17609 1998
rect 17491 1589 17609 1601
rect 17725 1998 17843 2010
rect 17725 1601 17731 1998
rect 17837 1601 17843 1998
rect 17725 1589 17843 1601
rect 17959 1998 18077 2010
rect 17959 1601 17965 1998
rect 18071 1601 18077 1998
rect 17959 1589 18077 1601
rect 18193 1998 18311 2010
rect 18193 1601 18199 1998
rect 18305 1601 18311 1998
rect 18193 1589 18311 1601
rect 18427 1998 18545 2010
rect 18427 1601 18433 1998
rect 18539 1601 18545 1998
rect 18427 1589 18545 1601
rect 18661 1998 18779 2010
rect 18661 1601 18667 1998
rect 18773 1601 18779 1998
rect 18661 1589 18779 1601
rect 18895 1998 19013 2010
rect 18895 1601 18901 1998
rect 19007 1601 19013 1998
rect 18895 1589 19013 1601
rect 19129 1998 19247 2010
rect 19129 1601 19135 1998
rect 19241 1601 19247 1998
rect 19129 1589 19247 1601
rect 19363 1998 19481 2010
rect 19363 1601 19369 1998
rect 19475 1601 19481 1998
rect 19363 1589 19481 1601
rect 19597 1998 19715 2010
rect 19597 1601 19603 1998
rect 19709 1601 19715 1998
rect 19597 1589 19715 1601
rect 19831 1998 19949 2010
rect 19831 1601 19837 1998
rect 19943 1601 19949 1998
rect 19831 1589 19949 1601
rect 20065 1998 20183 2010
rect 20065 1601 20071 1998
rect 20177 1601 20183 1998
rect 20065 1589 20183 1601
rect 20299 1998 20417 2010
rect 20299 1601 20305 1998
rect 20411 1601 20417 1998
rect 20299 1589 20417 1601
rect 20533 1998 20651 2010
rect 20533 1601 20539 1998
rect 20645 1601 20651 1998
rect 20533 1589 20651 1601
rect 20767 1998 20885 2010
rect 20767 1601 20773 1998
rect 20879 1601 20885 1998
rect 20767 1589 20885 1601
rect 21001 1998 21119 2010
rect 21001 1601 21007 1998
rect 21113 1601 21119 1998
rect 21001 1589 21119 1601
rect 21235 1998 21353 2010
rect 21235 1601 21241 1998
rect 21347 1601 21353 1998
rect 21235 1589 21353 1601
rect 21469 1998 21587 2010
rect 21469 1601 21475 1998
rect 21581 1601 21587 1998
rect 21469 1589 21587 1601
rect 21703 1998 21821 2010
rect 21703 1601 21709 1998
rect 21815 1601 21821 1998
rect 21703 1589 21821 1601
rect 21937 1998 22055 2010
rect 21937 1601 21943 1998
rect 22049 1601 22055 1998
rect 21937 1589 22055 1601
rect 22171 1998 22289 2010
rect 22171 1601 22177 1998
rect 22283 1601 22289 1998
rect 22171 1589 22289 1601
rect 22405 1998 22523 2010
rect 22405 1601 22411 1998
rect 22517 1601 22523 1998
rect 22405 1589 22523 1601
rect 22639 1998 22757 2010
rect 22639 1601 22645 1998
rect 22751 1601 22757 1998
rect 22639 1589 22757 1601
rect 22873 1998 22991 2010
rect 22873 1601 22879 1998
rect 22985 1601 22991 1998
rect 22873 1589 22991 1601
rect 23107 1998 23225 2010
rect 23107 1601 23113 1998
rect 23219 1601 23225 1998
rect 23107 1589 23225 1601
rect 23341 1998 23459 2010
rect 23341 1601 23347 1998
rect 23453 1601 23459 1998
rect 23341 1589 23459 1601
rect -23459 -1601 -23341 -1589
rect -23459 -1998 -23453 -1601
rect -23347 -1998 -23341 -1601
rect -23459 -2010 -23341 -1998
rect -23225 -1601 -23107 -1589
rect -23225 -1998 -23219 -1601
rect -23113 -1998 -23107 -1601
rect -23225 -2010 -23107 -1998
rect -22991 -1601 -22873 -1589
rect -22991 -1998 -22985 -1601
rect -22879 -1998 -22873 -1601
rect -22991 -2010 -22873 -1998
rect -22757 -1601 -22639 -1589
rect -22757 -1998 -22751 -1601
rect -22645 -1998 -22639 -1601
rect -22757 -2010 -22639 -1998
rect -22523 -1601 -22405 -1589
rect -22523 -1998 -22517 -1601
rect -22411 -1998 -22405 -1601
rect -22523 -2010 -22405 -1998
rect -22289 -1601 -22171 -1589
rect -22289 -1998 -22283 -1601
rect -22177 -1998 -22171 -1601
rect -22289 -2010 -22171 -1998
rect -22055 -1601 -21937 -1589
rect -22055 -1998 -22049 -1601
rect -21943 -1998 -21937 -1601
rect -22055 -2010 -21937 -1998
rect -21821 -1601 -21703 -1589
rect -21821 -1998 -21815 -1601
rect -21709 -1998 -21703 -1601
rect -21821 -2010 -21703 -1998
rect -21587 -1601 -21469 -1589
rect -21587 -1998 -21581 -1601
rect -21475 -1998 -21469 -1601
rect -21587 -2010 -21469 -1998
rect -21353 -1601 -21235 -1589
rect -21353 -1998 -21347 -1601
rect -21241 -1998 -21235 -1601
rect -21353 -2010 -21235 -1998
rect -21119 -1601 -21001 -1589
rect -21119 -1998 -21113 -1601
rect -21007 -1998 -21001 -1601
rect -21119 -2010 -21001 -1998
rect -20885 -1601 -20767 -1589
rect -20885 -1998 -20879 -1601
rect -20773 -1998 -20767 -1601
rect -20885 -2010 -20767 -1998
rect -20651 -1601 -20533 -1589
rect -20651 -1998 -20645 -1601
rect -20539 -1998 -20533 -1601
rect -20651 -2010 -20533 -1998
rect -20417 -1601 -20299 -1589
rect -20417 -1998 -20411 -1601
rect -20305 -1998 -20299 -1601
rect -20417 -2010 -20299 -1998
rect -20183 -1601 -20065 -1589
rect -20183 -1998 -20177 -1601
rect -20071 -1998 -20065 -1601
rect -20183 -2010 -20065 -1998
rect -19949 -1601 -19831 -1589
rect -19949 -1998 -19943 -1601
rect -19837 -1998 -19831 -1601
rect -19949 -2010 -19831 -1998
rect -19715 -1601 -19597 -1589
rect -19715 -1998 -19709 -1601
rect -19603 -1998 -19597 -1601
rect -19715 -2010 -19597 -1998
rect -19481 -1601 -19363 -1589
rect -19481 -1998 -19475 -1601
rect -19369 -1998 -19363 -1601
rect -19481 -2010 -19363 -1998
rect -19247 -1601 -19129 -1589
rect -19247 -1998 -19241 -1601
rect -19135 -1998 -19129 -1601
rect -19247 -2010 -19129 -1998
rect -19013 -1601 -18895 -1589
rect -19013 -1998 -19007 -1601
rect -18901 -1998 -18895 -1601
rect -19013 -2010 -18895 -1998
rect -18779 -1601 -18661 -1589
rect -18779 -1998 -18773 -1601
rect -18667 -1998 -18661 -1601
rect -18779 -2010 -18661 -1998
rect -18545 -1601 -18427 -1589
rect -18545 -1998 -18539 -1601
rect -18433 -1998 -18427 -1601
rect -18545 -2010 -18427 -1998
rect -18311 -1601 -18193 -1589
rect -18311 -1998 -18305 -1601
rect -18199 -1998 -18193 -1601
rect -18311 -2010 -18193 -1998
rect -18077 -1601 -17959 -1589
rect -18077 -1998 -18071 -1601
rect -17965 -1998 -17959 -1601
rect -18077 -2010 -17959 -1998
rect -17843 -1601 -17725 -1589
rect -17843 -1998 -17837 -1601
rect -17731 -1998 -17725 -1601
rect -17843 -2010 -17725 -1998
rect -17609 -1601 -17491 -1589
rect -17609 -1998 -17603 -1601
rect -17497 -1998 -17491 -1601
rect -17609 -2010 -17491 -1998
rect -17375 -1601 -17257 -1589
rect -17375 -1998 -17369 -1601
rect -17263 -1998 -17257 -1601
rect -17375 -2010 -17257 -1998
rect -17141 -1601 -17023 -1589
rect -17141 -1998 -17135 -1601
rect -17029 -1998 -17023 -1601
rect -17141 -2010 -17023 -1998
rect -16907 -1601 -16789 -1589
rect -16907 -1998 -16901 -1601
rect -16795 -1998 -16789 -1601
rect -16907 -2010 -16789 -1998
rect -16673 -1601 -16555 -1589
rect -16673 -1998 -16667 -1601
rect -16561 -1998 -16555 -1601
rect -16673 -2010 -16555 -1998
rect -16439 -1601 -16321 -1589
rect -16439 -1998 -16433 -1601
rect -16327 -1998 -16321 -1601
rect -16439 -2010 -16321 -1998
rect -16205 -1601 -16087 -1589
rect -16205 -1998 -16199 -1601
rect -16093 -1998 -16087 -1601
rect -16205 -2010 -16087 -1998
rect -15971 -1601 -15853 -1589
rect -15971 -1998 -15965 -1601
rect -15859 -1998 -15853 -1601
rect -15971 -2010 -15853 -1998
rect -15737 -1601 -15619 -1589
rect -15737 -1998 -15731 -1601
rect -15625 -1998 -15619 -1601
rect -15737 -2010 -15619 -1998
rect -15503 -1601 -15385 -1589
rect -15503 -1998 -15497 -1601
rect -15391 -1998 -15385 -1601
rect -15503 -2010 -15385 -1998
rect -15269 -1601 -15151 -1589
rect -15269 -1998 -15263 -1601
rect -15157 -1998 -15151 -1601
rect -15269 -2010 -15151 -1998
rect -15035 -1601 -14917 -1589
rect -15035 -1998 -15029 -1601
rect -14923 -1998 -14917 -1601
rect -15035 -2010 -14917 -1998
rect -14801 -1601 -14683 -1589
rect -14801 -1998 -14795 -1601
rect -14689 -1998 -14683 -1601
rect -14801 -2010 -14683 -1998
rect -14567 -1601 -14449 -1589
rect -14567 -1998 -14561 -1601
rect -14455 -1998 -14449 -1601
rect -14567 -2010 -14449 -1998
rect -14333 -1601 -14215 -1589
rect -14333 -1998 -14327 -1601
rect -14221 -1998 -14215 -1601
rect -14333 -2010 -14215 -1998
rect -14099 -1601 -13981 -1589
rect -14099 -1998 -14093 -1601
rect -13987 -1998 -13981 -1601
rect -14099 -2010 -13981 -1998
rect -13865 -1601 -13747 -1589
rect -13865 -1998 -13859 -1601
rect -13753 -1998 -13747 -1601
rect -13865 -2010 -13747 -1998
rect -13631 -1601 -13513 -1589
rect -13631 -1998 -13625 -1601
rect -13519 -1998 -13513 -1601
rect -13631 -2010 -13513 -1998
rect -13397 -1601 -13279 -1589
rect -13397 -1998 -13391 -1601
rect -13285 -1998 -13279 -1601
rect -13397 -2010 -13279 -1998
rect -13163 -1601 -13045 -1589
rect -13163 -1998 -13157 -1601
rect -13051 -1998 -13045 -1601
rect -13163 -2010 -13045 -1998
rect -12929 -1601 -12811 -1589
rect -12929 -1998 -12923 -1601
rect -12817 -1998 -12811 -1601
rect -12929 -2010 -12811 -1998
rect -12695 -1601 -12577 -1589
rect -12695 -1998 -12689 -1601
rect -12583 -1998 -12577 -1601
rect -12695 -2010 -12577 -1998
rect -12461 -1601 -12343 -1589
rect -12461 -1998 -12455 -1601
rect -12349 -1998 -12343 -1601
rect -12461 -2010 -12343 -1998
rect -12227 -1601 -12109 -1589
rect -12227 -1998 -12221 -1601
rect -12115 -1998 -12109 -1601
rect -12227 -2010 -12109 -1998
rect -11993 -1601 -11875 -1589
rect -11993 -1998 -11987 -1601
rect -11881 -1998 -11875 -1601
rect -11993 -2010 -11875 -1998
rect -11759 -1601 -11641 -1589
rect -11759 -1998 -11753 -1601
rect -11647 -1998 -11641 -1601
rect -11759 -2010 -11641 -1998
rect -11525 -1601 -11407 -1589
rect -11525 -1998 -11519 -1601
rect -11413 -1998 -11407 -1601
rect -11525 -2010 -11407 -1998
rect -11291 -1601 -11173 -1589
rect -11291 -1998 -11285 -1601
rect -11179 -1998 -11173 -1601
rect -11291 -2010 -11173 -1998
rect -11057 -1601 -10939 -1589
rect -11057 -1998 -11051 -1601
rect -10945 -1998 -10939 -1601
rect -11057 -2010 -10939 -1998
rect -10823 -1601 -10705 -1589
rect -10823 -1998 -10817 -1601
rect -10711 -1998 -10705 -1601
rect -10823 -2010 -10705 -1998
rect -10589 -1601 -10471 -1589
rect -10589 -1998 -10583 -1601
rect -10477 -1998 -10471 -1601
rect -10589 -2010 -10471 -1998
rect -10355 -1601 -10237 -1589
rect -10355 -1998 -10349 -1601
rect -10243 -1998 -10237 -1601
rect -10355 -2010 -10237 -1998
rect -10121 -1601 -10003 -1589
rect -10121 -1998 -10115 -1601
rect -10009 -1998 -10003 -1601
rect -10121 -2010 -10003 -1998
rect -9887 -1601 -9769 -1589
rect -9887 -1998 -9881 -1601
rect -9775 -1998 -9769 -1601
rect -9887 -2010 -9769 -1998
rect -9653 -1601 -9535 -1589
rect -9653 -1998 -9647 -1601
rect -9541 -1998 -9535 -1601
rect -9653 -2010 -9535 -1998
rect -9419 -1601 -9301 -1589
rect -9419 -1998 -9413 -1601
rect -9307 -1998 -9301 -1601
rect -9419 -2010 -9301 -1998
rect -9185 -1601 -9067 -1589
rect -9185 -1998 -9179 -1601
rect -9073 -1998 -9067 -1601
rect -9185 -2010 -9067 -1998
rect -8951 -1601 -8833 -1589
rect -8951 -1998 -8945 -1601
rect -8839 -1998 -8833 -1601
rect -8951 -2010 -8833 -1998
rect -8717 -1601 -8599 -1589
rect -8717 -1998 -8711 -1601
rect -8605 -1998 -8599 -1601
rect -8717 -2010 -8599 -1998
rect -8483 -1601 -8365 -1589
rect -8483 -1998 -8477 -1601
rect -8371 -1998 -8365 -1601
rect -8483 -2010 -8365 -1998
rect -8249 -1601 -8131 -1589
rect -8249 -1998 -8243 -1601
rect -8137 -1998 -8131 -1601
rect -8249 -2010 -8131 -1998
rect -8015 -1601 -7897 -1589
rect -8015 -1998 -8009 -1601
rect -7903 -1998 -7897 -1601
rect -8015 -2010 -7897 -1998
rect -7781 -1601 -7663 -1589
rect -7781 -1998 -7775 -1601
rect -7669 -1998 -7663 -1601
rect -7781 -2010 -7663 -1998
rect -7547 -1601 -7429 -1589
rect -7547 -1998 -7541 -1601
rect -7435 -1998 -7429 -1601
rect -7547 -2010 -7429 -1998
rect -7313 -1601 -7195 -1589
rect -7313 -1998 -7307 -1601
rect -7201 -1998 -7195 -1601
rect -7313 -2010 -7195 -1998
rect -7079 -1601 -6961 -1589
rect -7079 -1998 -7073 -1601
rect -6967 -1998 -6961 -1601
rect -7079 -2010 -6961 -1998
rect -6845 -1601 -6727 -1589
rect -6845 -1998 -6839 -1601
rect -6733 -1998 -6727 -1601
rect -6845 -2010 -6727 -1998
rect -6611 -1601 -6493 -1589
rect -6611 -1998 -6605 -1601
rect -6499 -1998 -6493 -1601
rect -6611 -2010 -6493 -1998
rect -6377 -1601 -6259 -1589
rect -6377 -1998 -6371 -1601
rect -6265 -1998 -6259 -1601
rect -6377 -2010 -6259 -1998
rect -6143 -1601 -6025 -1589
rect -6143 -1998 -6137 -1601
rect -6031 -1998 -6025 -1601
rect -6143 -2010 -6025 -1998
rect -5909 -1601 -5791 -1589
rect -5909 -1998 -5903 -1601
rect -5797 -1998 -5791 -1601
rect -5909 -2010 -5791 -1998
rect -5675 -1601 -5557 -1589
rect -5675 -1998 -5669 -1601
rect -5563 -1998 -5557 -1601
rect -5675 -2010 -5557 -1998
rect -5441 -1601 -5323 -1589
rect -5441 -1998 -5435 -1601
rect -5329 -1998 -5323 -1601
rect -5441 -2010 -5323 -1998
rect -5207 -1601 -5089 -1589
rect -5207 -1998 -5201 -1601
rect -5095 -1998 -5089 -1601
rect -5207 -2010 -5089 -1998
rect -4973 -1601 -4855 -1589
rect -4973 -1998 -4967 -1601
rect -4861 -1998 -4855 -1601
rect -4973 -2010 -4855 -1998
rect -4739 -1601 -4621 -1589
rect -4739 -1998 -4733 -1601
rect -4627 -1998 -4621 -1601
rect -4739 -2010 -4621 -1998
rect -4505 -1601 -4387 -1589
rect -4505 -1998 -4499 -1601
rect -4393 -1998 -4387 -1601
rect -4505 -2010 -4387 -1998
rect -4271 -1601 -4153 -1589
rect -4271 -1998 -4265 -1601
rect -4159 -1998 -4153 -1601
rect -4271 -2010 -4153 -1998
rect -4037 -1601 -3919 -1589
rect -4037 -1998 -4031 -1601
rect -3925 -1998 -3919 -1601
rect -4037 -2010 -3919 -1998
rect -3803 -1601 -3685 -1589
rect -3803 -1998 -3797 -1601
rect -3691 -1998 -3685 -1601
rect -3803 -2010 -3685 -1998
rect -3569 -1601 -3451 -1589
rect -3569 -1998 -3563 -1601
rect -3457 -1998 -3451 -1601
rect -3569 -2010 -3451 -1998
rect -3335 -1601 -3217 -1589
rect -3335 -1998 -3329 -1601
rect -3223 -1998 -3217 -1601
rect -3335 -2010 -3217 -1998
rect -3101 -1601 -2983 -1589
rect -3101 -1998 -3095 -1601
rect -2989 -1998 -2983 -1601
rect -3101 -2010 -2983 -1998
rect -2867 -1601 -2749 -1589
rect -2867 -1998 -2861 -1601
rect -2755 -1998 -2749 -1601
rect -2867 -2010 -2749 -1998
rect -2633 -1601 -2515 -1589
rect -2633 -1998 -2627 -1601
rect -2521 -1998 -2515 -1601
rect -2633 -2010 -2515 -1998
rect -2399 -1601 -2281 -1589
rect -2399 -1998 -2393 -1601
rect -2287 -1998 -2281 -1601
rect -2399 -2010 -2281 -1998
rect -2165 -1601 -2047 -1589
rect -2165 -1998 -2159 -1601
rect -2053 -1998 -2047 -1601
rect -2165 -2010 -2047 -1998
rect -1931 -1601 -1813 -1589
rect -1931 -1998 -1925 -1601
rect -1819 -1998 -1813 -1601
rect -1931 -2010 -1813 -1998
rect -1697 -1601 -1579 -1589
rect -1697 -1998 -1691 -1601
rect -1585 -1998 -1579 -1601
rect -1697 -2010 -1579 -1998
rect -1463 -1601 -1345 -1589
rect -1463 -1998 -1457 -1601
rect -1351 -1998 -1345 -1601
rect -1463 -2010 -1345 -1998
rect -1229 -1601 -1111 -1589
rect -1229 -1998 -1223 -1601
rect -1117 -1998 -1111 -1601
rect -1229 -2010 -1111 -1998
rect -995 -1601 -877 -1589
rect -995 -1998 -989 -1601
rect -883 -1998 -877 -1601
rect -995 -2010 -877 -1998
rect -761 -1601 -643 -1589
rect -761 -1998 -755 -1601
rect -649 -1998 -643 -1601
rect -761 -2010 -643 -1998
rect -527 -1601 -409 -1589
rect -527 -1998 -521 -1601
rect -415 -1998 -409 -1601
rect -527 -2010 -409 -1998
rect -293 -1601 -175 -1589
rect -293 -1998 -287 -1601
rect -181 -1998 -175 -1601
rect -293 -2010 -175 -1998
rect -59 -1601 59 -1589
rect -59 -1998 -53 -1601
rect 53 -1998 59 -1601
rect -59 -2010 59 -1998
rect 175 -1601 293 -1589
rect 175 -1998 181 -1601
rect 287 -1998 293 -1601
rect 175 -2010 293 -1998
rect 409 -1601 527 -1589
rect 409 -1998 415 -1601
rect 521 -1998 527 -1601
rect 409 -2010 527 -1998
rect 643 -1601 761 -1589
rect 643 -1998 649 -1601
rect 755 -1998 761 -1601
rect 643 -2010 761 -1998
rect 877 -1601 995 -1589
rect 877 -1998 883 -1601
rect 989 -1998 995 -1601
rect 877 -2010 995 -1998
rect 1111 -1601 1229 -1589
rect 1111 -1998 1117 -1601
rect 1223 -1998 1229 -1601
rect 1111 -2010 1229 -1998
rect 1345 -1601 1463 -1589
rect 1345 -1998 1351 -1601
rect 1457 -1998 1463 -1601
rect 1345 -2010 1463 -1998
rect 1579 -1601 1697 -1589
rect 1579 -1998 1585 -1601
rect 1691 -1998 1697 -1601
rect 1579 -2010 1697 -1998
rect 1813 -1601 1931 -1589
rect 1813 -1998 1819 -1601
rect 1925 -1998 1931 -1601
rect 1813 -2010 1931 -1998
rect 2047 -1601 2165 -1589
rect 2047 -1998 2053 -1601
rect 2159 -1998 2165 -1601
rect 2047 -2010 2165 -1998
rect 2281 -1601 2399 -1589
rect 2281 -1998 2287 -1601
rect 2393 -1998 2399 -1601
rect 2281 -2010 2399 -1998
rect 2515 -1601 2633 -1589
rect 2515 -1998 2521 -1601
rect 2627 -1998 2633 -1601
rect 2515 -2010 2633 -1998
rect 2749 -1601 2867 -1589
rect 2749 -1998 2755 -1601
rect 2861 -1998 2867 -1601
rect 2749 -2010 2867 -1998
rect 2983 -1601 3101 -1589
rect 2983 -1998 2989 -1601
rect 3095 -1998 3101 -1601
rect 2983 -2010 3101 -1998
rect 3217 -1601 3335 -1589
rect 3217 -1998 3223 -1601
rect 3329 -1998 3335 -1601
rect 3217 -2010 3335 -1998
rect 3451 -1601 3569 -1589
rect 3451 -1998 3457 -1601
rect 3563 -1998 3569 -1601
rect 3451 -2010 3569 -1998
rect 3685 -1601 3803 -1589
rect 3685 -1998 3691 -1601
rect 3797 -1998 3803 -1601
rect 3685 -2010 3803 -1998
rect 3919 -1601 4037 -1589
rect 3919 -1998 3925 -1601
rect 4031 -1998 4037 -1601
rect 3919 -2010 4037 -1998
rect 4153 -1601 4271 -1589
rect 4153 -1998 4159 -1601
rect 4265 -1998 4271 -1601
rect 4153 -2010 4271 -1998
rect 4387 -1601 4505 -1589
rect 4387 -1998 4393 -1601
rect 4499 -1998 4505 -1601
rect 4387 -2010 4505 -1998
rect 4621 -1601 4739 -1589
rect 4621 -1998 4627 -1601
rect 4733 -1998 4739 -1601
rect 4621 -2010 4739 -1998
rect 4855 -1601 4973 -1589
rect 4855 -1998 4861 -1601
rect 4967 -1998 4973 -1601
rect 4855 -2010 4973 -1998
rect 5089 -1601 5207 -1589
rect 5089 -1998 5095 -1601
rect 5201 -1998 5207 -1601
rect 5089 -2010 5207 -1998
rect 5323 -1601 5441 -1589
rect 5323 -1998 5329 -1601
rect 5435 -1998 5441 -1601
rect 5323 -2010 5441 -1998
rect 5557 -1601 5675 -1589
rect 5557 -1998 5563 -1601
rect 5669 -1998 5675 -1601
rect 5557 -2010 5675 -1998
rect 5791 -1601 5909 -1589
rect 5791 -1998 5797 -1601
rect 5903 -1998 5909 -1601
rect 5791 -2010 5909 -1998
rect 6025 -1601 6143 -1589
rect 6025 -1998 6031 -1601
rect 6137 -1998 6143 -1601
rect 6025 -2010 6143 -1998
rect 6259 -1601 6377 -1589
rect 6259 -1998 6265 -1601
rect 6371 -1998 6377 -1601
rect 6259 -2010 6377 -1998
rect 6493 -1601 6611 -1589
rect 6493 -1998 6499 -1601
rect 6605 -1998 6611 -1601
rect 6493 -2010 6611 -1998
rect 6727 -1601 6845 -1589
rect 6727 -1998 6733 -1601
rect 6839 -1998 6845 -1601
rect 6727 -2010 6845 -1998
rect 6961 -1601 7079 -1589
rect 6961 -1998 6967 -1601
rect 7073 -1998 7079 -1601
rect 6961 -2010 7079 -1998
rect 7195 -1601 7313 -1589
rect 7195 -1998 7201 -1601
rect 7307 -1998 7313 -1601
rect 7195 -2010 7313 -1998
rect 7429 -1601 7547 -1589
rect 7429 -1998 7435 -1601
rect 7541 -1998 7547 -1601
rect 7429 -2010 7547 -1998
rect 7663 -1601 7781 -1589
rect 7663 -1998 7669 -1601
rect 7775 -1998 7781 -1601
rect 7663 -2010 7781 -1998
rect 7897 -1601 8015 -1589
rect 7897 -1998 7903 -1601
rect 8009 -1998 8015 -1601
rect 7897 -2010 8015 -1998
rect 8131 -1601 8249 -1589
rect 8131 -1998 8137 -1601
rect 8243 -1998 8249 -1601
rect 8131 -2010 8249 -1998
rect 8365 -1601 8483 -1589
rect 8365 -1998 8371 -1601
rect 8477 -1998 8483 -1601
rect 8365 -2010 8483 -1998
rect 8599 -1601 8717 -1589
rect 8599 -1998 8605 -1601
rect 8711 -1998 8717 -1601
rect 8599 -2010 8717 -1998
rect 8833 -1601 8951 -1589
rect 8833 -1998 8839 -1601
rect 8945 -1998 8951 -1601
rect 8833 -2010 8951 -1998
rect 9067 -1601 9185 -1589
rect 9067 -1998 9073 -1601
rect 9179 -1998 9185 -1601
rect 9067 -2010 9185 -1998
rect 9301 -1601 9419 -1589
rect 9301 -1998 9307 -1601
rect 9413 -1998 9419 -1601
rect 9301 -2010 9419 -1998
rect 9535 -1601 9653 -1589
rect 9535 -1998 9541 -1601
rect 9647 -1998 9653 -1601
rect 9535 -2010 9653 -1998
rect 9769 -1601 9887 -1589
rect 9769 -1998 9775 -1601
rect 9881 -1998 9887 -1601
rect 9769 -2010 9887 -1998
rect 10003 -1601 10121 -1589
rect 10003 -1998 10009 -1601
rect 10115 -1998 10121 -1601
rect 10003 -2010 10121 -1998
rect 10237 -1601 10355 -1589
rect 10237 -1998 10243 -1601
rect 10349 -1998 10355 -1601
rect 10237 -2010 10355 -1998
rect 10471 -1601 10589 -1589
rect 10471 -1998 10477 -1601
rect 10583 -1998 10589 -1601
rect 10471 -2010 10589 -1998
rect 10705 -1601 10823 -1589
rect 10705 -1998 10711 -1601
rect 10817 -1998 10823 -1601
rect 10705 -2010 10823 -1998
rect 10939 -1601 11057 -1589
rect 10939 -1998 10945 -1601
rect 11051 -1998 11057 -1601
rect 10939 -2010 11057 -1998
rect 11173 -1601 11291 -1589
rect 11173 -1998 11179 -1601
rect 11285 -1998 11291 -1601
rect 11173 -2010 11291 -1998
rect 11407 -1601 11525 -1589
rect 11407 -1998 11413 -1601
rect 11519 -1998 11525 -1601
rect 11407 -2010 11525 -1998
rect 11641 -1601 11759 -1589
rect 11641 -1998 11647 -1601
rect 11753 -1998 11759 -1601
rect 11641 -2010 11759 -1998
rect 11875 -1601 11993 -1589
rect 11875 -1998 11881 -1601
rect 11987 -1998 11993 -1601
rect 11875 -2010 11993 -1998
rect 12109 -1601 12227 -1589
rect 12109 -1998 12115 -1601
rect 12221 -1998 12227 -1601
rect 12109 -2010 12227 -1998
rect 12343 -1601 12461 -1589
rect 12343 -1998 12349 -1601
rect 12455 -1998 12461 -1601
rect 12343 -2010 12461 -1998
rect 12577 -1601 12695 -1589
rect 12577 -1998 12583 -1601
rect 12689 -1998 12695 -1601
rect 12577 -2010 12695 -1998
rect 12811 -1601 12929 -1589
rect 12811 -1998 12817 -1601
rect 12923 -1998 12929 -1601
rect 12811 -2010 12929 -1998
rect 13045 -1601 13163 -1589
rect 13045 -1998 13051 -1601
rect 13157 -1998 13163 -1601
rect 13045 -2010 13163 -1998
rect 13279 -1601 13397 -1589
rect 13279 -1998 13285 -1601
rect 13391 -1998 13397 -1601
rect 13279 -2010 13397 -1998
rect 13513 -1601 13631 -1589
rect 13513 -1998 13519 -1601
rect 13625 -1998 13631 -1601
rect 13513 -2010 13631 -1998
rect 13747 -1601 13865 -1589
rect 13747 -1998 13753 -1601
rect 13859 -1998 13865 -1601
rect 13747 -2010 13865 -1998
rect 13981 -1601 14099 -1589
rect 13981 -1998 13987 -1601
rect 14093 -1998 14099 -1601
rect 13981 -2010 14099 -1998
rect 14215 -1601 14333 -1589
rect 14215 -1998 14221 -1601
rect 14327 -1998 14333 -1601
rect 14215 -2010 14333 -1998
rect 14449 -1601 14567 -1589
rect 14449 -1998 14455 -1601
rect 14561 -1998 14567 -1601
rect 14449 -2010 14567 -1998
rect 14683 -1601 14801 -1589
rect 14683 -1998 14689 -1601
rect 14795 -1998 14801 -1601
rect 14683 -2010 14801 -1998
rect 14917 -1601 15035 -1589
rect 14917 -1998 14923 -1601
rect 15029 -1998 15035 -1601
rect 14917 -2010 15035 -1998
rect 15151 -1601 15269 -1589
rect 15151 -1998 15157 -1601
rect 15263 -1998 15269 -1601
rect 15151 -2010 15269 -1998
rect 15385 -1601 15503 -1589
rect 15385 -1998 15391 -1601
rect 15497 -1998 15503 -1601
rect 15385 -2010 15503 -1998
rect 15619 -1601 15737 -1589
rect 15619 -1998 15625 -1601
rect 15731 -1998 15737 -1601
rect 15619 -2010 15737 -1998
rect 15853 -1601 15971 -1589
rect 15853 -1998 15859 -1601
rect 15965 -1998 15971 -1601
rect 15853 -2010 15971 -1998
rect 16087 -1601 16205 -1589
rect 16087 -1998 16093 -1601
rect 16199 -1998 16205 -1601
rect 16087 -2010 16205 -1998
rect 16321 -1601 16439 -1589
rect 16321 -1998 16327 -1601
rect 16433 -1998 16439 -1601
rect 16321 -2010 16439 -1998
rect 16555 -1601 16673 -1589
rect 16555 -1998 16561 -1601
rect 16667 -1998 16673 -1601
rect 16555 -2010 16673 -1998
rect 16789 -1601 16907 -1589
rect 16789 -1998 16795 -1601
rect 16901 -1998 16907 -1601
rect 16789 -2010 16907 -1998
rect 17023 -1601 17141 -1589
rect 17023 -1998 17029 -1601
rect 17135 -1998 17141 -1601
rect 17023 -2010 17141 -1998
rect 17257 -1601 17375 -1589
rect 17257 -1998 17263 -1601
rect 17369 -1998 17375 -1601
rect 17257 -2010 17375 -1998
rect 17491 -1601 17609 -1589
rect 17491 -1998 17497 -1601
rect 17603 -1998 17609 -1601
rect 17491 -2010 17609 -1998
rect 17725 -1601 17843 -1589
rect 17725 -1998 17731 -1601
rect 17837 -1998 17843 -1601
rect 17725 -2010 17843 -1998
rect 17959 -1601 18077 -1589
rect 17959 -1998 17965 -1601
rect 18071 -1998 18077 -1601
rect 17959 -2010 18077 -1998
rect 18193 -1601 18311 -1589
rect 18193 -1998 18199 -1601
rect 18305 -1998 18311 -1601
rect 18193 -2010 18311 -1998
rect 18427 -1601 18545 -1589
rect 18427 -1998 18433 -1601
rect 18539 -1998 18545 -1601
rect 18427 -2010 18545 -1998
rect 18661 -1601 18779 -1589
rect 18661 -1998 18667 -1601
rect 18773 -1998 18779 -1601
rect 18661 -2010 18779 -1998
rect 18895 -1601 19013 -1589
rect 18895 -1998 18901 -1601
rect 19007 -1998 19013 -1601
rect 18895 -2010 19013 -1998
rect 19129 -1601 19247 -1589
rect 19129 -1998 19135 -1601
rect 19241 -1998 19247 -1601
rect 19129 -2010 19247 -1998
rect 19363 -1601 19481 -1589
rect 19363 -1998 19369 -1601
rect 19475 -1998 19481 -1601
rect 19363 -2010 19481 -1998
rect 19597 -1601 19715 -1589
rect 19597 -1998 19603 -1601
rect 19709 -1998 19715 -1601
rect 19597 -2010 19715 -1998
rect 19831 -1601 19949 -1589
rect 19831 -1998 19837 -1601
rect 19943 -1998 19949 -1601
rect 19831 -2010 19949 -1998
rect 20065 -1601 20183 -1589
rect 20065 -1998 20071 -1601
rect 20177 -1998 20183 -1601
rect 20065 -2010 20183 -1998
rect 20299 -1601 20417 -1589
rect 20299 -1998 20305 -1601
rect 20411 -1998 20417 -1601
rect 20299 -2010 20417 -1998
rect 20533 -1601 20651 -1589
rect 20533 -1998 20539 -1601
rect 20645 -1998 20651 -1601
rect 20533 -2010 20651 -1998
rect 20767 -1601 20885 -1589
rect 20767 -1998 20773 -1601
rect 20879 -1998 20885 -1601
rect 20767 -2010 20885 -1998
rect 21001 -1601 21119 -1589
rect 21001 -1998 21007 -1601
rect 21113 -1998 21119 -1601
rect 21001 -2010 21119 -1998
rect 21235 -1601 21353 -1589
rect 21235 -1998 21241 -1601
rect 21347 -1998 21353 -1601
rect 21235 -2010 21353 -1998
rect 21469 -1601 21587 -1589
rect 21469 -1998 21475 -1601
rect 21581 -1998 21587 -1601
rect 21469 -2010 21587 -1998
rect 21703 -1601 21821 -1589
rect 21703 -1998 21709 -1601
rect 21815 -1998 21821 -1601
rect 21703 -2010 21821 -1998
rect 21937 -1601 22055 -1589
rect 21937 -1998 21943 -1601
rect 22049 -1998 22055 -1601
rect 21937 -2010 22055 -1998
rect 22171 -1601 22289 -1589
rect 22171 -1998 22177 -1601
rect 22283 -1998 22289 -1601
rect 22171 -2010 22289 -1998
rect 22405 -1601 22523 -1589
rect 22405 -1998 22411 -1601
rect 22517 -1998 22523 -1601
rect 22405 -2010 22523 -1998
rect 22639 -1601 22757 -1589
rect 22639 -1998 22645 -1601
rect 22751 -1998 22757 -1601
rect 22639 -2010 22757 -1998
rect 22873 -1601 22991 -1589
rect 22873 -1998 22879 -1601
rect 22985 -1998 22991 -1601
rect 22873 -2010 22991 -1998
rect 23107 -1601 23225 -1589
rect 23107 -1998 23113 -1601
rect 23219 -1998 23225 -1601
rect 23107 -2010 23225 -1998
rect 23341 -1601 23459 -1589
rect 23341 -1998 23347 -1601
rect 23453 -1998 23459 -1601
rect 23341 -2010 23459 -1998
<< properties >>
string FIXED_BBOX -23582 -2129 23582 2129
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 16.0 m 1 nx 201 wmin 0.690 lmin 0.50 class resistor rho 319.8 val 7.98k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
