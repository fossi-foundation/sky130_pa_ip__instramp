magic
tech sky130A
magscale 1 2
timestamp 1729623223
<< pwell >>
rect -1446 -2307 1446 2307
<< psubdiff >>
rect -1410 2237 -1314 2271
rect 1314 2237 1410 2271
rect -1410 2175 -1376 2237
rect 1376 2175 1410 2237
rect -1410 -2237 -1376 -2175
rect 1376 -2237 1410 -2175
rect -1410 -2271 -1314 -2237
rect 1314 -2271 1410 -2237
<< psubdiffcont >>
rect -1314 2237 1314 2271
rect -1410 -2175 -1376 2175
rect 1376 -2175 1410 2175
rect -1314 -2271 1314 -2237
<< xpolycontact >>
rect -1280 1709 -1210 2141
rect -1280 -2141 -1210 -1709
rect -1114 1709 -1044 2141
rect -1114 -2141 -1044 -1709
rect -948 1709 -878 2141
rect -948 -2141 -878 -1709
rect -782 1709 -712 2141
rect -782 -2141 -712 -1709
rect -616 1709 -546 2141
rect -616 -2141 -546 -1709
rect -450 1709 -380 2141
rect -450 -2141 -380 -1709
rect -284 1709 -214 2141
rect -284 -2141 -214 -1709
rect -118 1709 -48 2141
rect -118 -2141 -48 -1709
rect 48 1709 118 2141
rect 48 -2141 118 -1709
rect 214 1709 284 2141
rect 214 -2141 284 -1709
rect 380 1709 450 2141
rect 380 -2141 450 -1709
rect 546 1709 616 2141
rect 546 -2141 616 -1709
rect 712 1709 782 2141
rect 712 -2141 782 -1709
rect 878 1709 948 2141
rect 878 -2141 948 -1709
rect 1044 1709 1114 2141
rect 1044 -2141 1114 -1709
rect 1210 1709 1280 2141
rect 1210 -2141 1280 -1709
<< xpolyres >>
rect -1280 -1709 -1210 1709
rect -1114 -1709 -1044 1709
rect -948 -1709 -878 1709
rect -782 -1709 -712 1709
rect -616 -1709 -546 1709
rect -450 -1709 -380 1709
rect -284 -1709 -214 1709
rect -118 -1709 -48 1709
rect 48 -1709 118 1709
rect 214 -1709 284 1709
rect 380 -1709 450 1709
rect 546 -1709 616 1709
rect 712 -1709 782 1709
rect 878 -1709 948 1709
rect 1044 -1709 1114 1709
rect 1210 -1709 1280 1709
<< locali >>
rect -1410 2237 -1314 2271
rect 1314 2237 1410 2271
rect -1410 2175 -1376 2237
rect 1376 2175 1410 2237
rect -1410 -2237 -1376 -2175
rect 1376 -2237 1410 -2175
rect -1410 -2271 -1314 -2237
rect 1314 -2271 1410 -2237
<< viali >>
rect -1264 1726 -1226 2123
rect -1098 1726 -1060 2123
rect -932 1726 -894 2123
rect -766 1726 -728 2123
rect -600 1726 -562 2123
rect -434 1726 -396 2123
rect -268 1726 -230 2123
rect -102 1726 -64 2123
rect 64 1726 102 2123
rect 230 1726 268 2123
rect 396 1726 434 2123
rect 562 1726 600 2123
rect 728 1726 766 2123
rect 894 1726 932 2123
rect 1060 1726 1098 2123
rect 1226 1726 1264 2123
rect -1264 -2123 -1226 -1726
rect -1098 -2123 -1060 -1726
rect -932 -2123 -894 -1726
rect -766 -2123 -728 -1726
rect -600 -2123 -562 -1726
rect -434 -2123 -396 -1726
rect -268 -2123 -230 -1726
rect -102 -2123 -64 -1726
rect 64 -2123 102 -1726
rect 230 -2123 268 -1726
rect 396 -2123 434 -1726
rect 562 -2123 600 -1726
rect 728 -2123 766 -1726
rect 894 -2123 932 -1726
rect 1060 -2123 1098 -1726
rect 1226 -2123 1264 -1726
<< metal1 >>
rect -1270 2123 -1220 2135
rect -1270 1726 -1264 2123
rect -1226 1726 -1220 2123
rect -1270 1714 -1220 1726
rect -1104 2123 -1054 2135
rect -1104 1726 -1098 2123
rect -1060 1726 -1054 2123
rect -1104 1714 -1054 1726
rect -938 2123 -888 2135
rect -938 1726 -932 2123
rect -894 1726 -888 2123
rect -938 1714 -888 1726
rect -772 2123 -722 2135
rect -772 1726 -766 2123
rect -728 1726 -722 2123
rect -772 1714 -722 1726
rect -606 2123 -556 2135
rect -606 1726 -600 2123
rect -562 1726 -556 2123
rect -606 1714 -556 1726
rect -440 2123 -390 2135
rect -440 1726 -434 2123
rect -396 1726 -390 2123
rect -440 1714 -390 1726
rect -274 2123 -224 2135
rect -274 1726 -268 2123
rect -230 1726 -224 2123
rect -274 1714 -224 1726
rect -108 2123 -58 2135
rect -108 1726 -102 2123
rect -64 1726 -58 2123
rect -108 1714 -58 1726
rect 58 2123 108 2135
rect 58 1726 64 2123
rect 102 1726 108 2123
rect 58 1714 108 1726
rect 224 2123 274 2135
rect 224 1726 230 2123
rect 268 1726 274 2123
rect 224 1714 274 1726
rect 390 2123 440 2135
rect 390 1726 396 2123
rect 434 1726 440 2123
rect 390 1714 440 1726
rect 556 2123 606 2135
rect 556 1726 562 2123
rect 600 1726 606 2123
rect 556 1714 606 1726
rect 722 2123 772 2135
rect 722 1726 728 2123
rect 766 1726 772 2123
rect 722 1714 772 1726
rect 888 2123 938 2135
rect 888 1726 894 2123
rect 932 1726 938 2123
rect 888 1714 938 1726
rect 1054 2123 1104 2135
rect 1054 1726 1060 2123
rect 1098 1726 1104 2123
rect 1054 1714 1104 1726
rect 1220 2123 1270 2135
rect 1220 1726 1226 2123
rect 1264 1726 1270 2123
rect 1220 1714 1270 1726
rect -1270 -1726 -1220 -1714
rect -1270 -2123 -1264 -1726
rect -1226 -2123 -1220 -1726
rect -1270 -2135 -1220 -2123
rect -1104 -1726 -1054 -1714
rect -1104 -2123 -1098 -1726
rect -1060 -2123 -1054 -1726
rect -1104 -2135 -1054 -2123
rect -938 -1726 -888 -1714
rect -938 -2123 -932 -1726
rect -894 -2123 -888 -1726
rect -938 -2135 -888 -2123
rect -772 -1726 -722 -1714
rect -772 -2123 -766 -1726
rect -728 -2123 -722 -1726
rect -772 -2135 -722 -2123
rect -606 -1726 -556 -1714
rect -606 -2123 -600 -1726
rect -562 -2123 -556 -1726
rect -606 -2135 -556 -2123
rect -440 -1726 -390 -1714
rect -440 -2123 -434 -1726
rect -396 -2123 -390 -1726
rect -440 -2135 -390 -2123
rect -274 -1726 -224 -1714
rect -274 -2123 -268 -1726
rect -230 -2123 -224 -1726
rect -274 -2135 -224 -2123
rect -108 -1726 -58 -1714
rect -108 -2123 -102 -1726
rect -64 -2123 -58 -1726
rect -108 -2135 -58 -2123
rect 58 -1726 108 -1714
rect 58 -2123 64 -1726
rect 102 -2123 108 -1726
rect 58 -2135 108 -2123
rect 224 -1726 274 -1714
rect 224 -2123 230 -1726
rect 268 -2123 274 -1726
rect 224 -2135 274 -2123
rect 390 -1726 440 -1714
rect 390 -2123 396 -1726
rect 434 -2123 440 -1726
rect 390 -2135 440 -2123
rect 556 -1726 606 -1714
rect 556 -2123 562 -1726
rect 600 -2123 606 -1726
rect 556 -2135 606 -2123
rect 722 -1726 772 -1714
rect 722 -2123 728 -1726
rect 766 -2123 772 -1726
rect 722 -2135 772 -2123
rect 888 -1726 938 -1714
rect 888 -2123 894 -1726
rect 932 -2123 938 -1726
rect 888 -2135 938 -2123
rect 1054 -1726 1104 -1714
rect 1054 -2123 1060 -1726
rect 1098 -2123 1104 -1726
rect 1054 -2135 1104 -2123
rect 1220 -1726 1270 -1714
rect 1220 -2123 1226 -1726
rect 1264 -2123 1270 -1726
rect 1220 -2135 1270 -2123
<< properties >>
string FIXED_BBOX -1393 -2254 1393 2254
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 17.25 m 1 nx 16 wmin 0.350 lmin 0.50 class resistor rho 2000 val 99.646k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
