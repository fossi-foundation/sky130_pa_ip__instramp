magic
tech sky130A
magscale 1 2
timestamp 1729620069
<< pwell >>
rect -9589 -2585 9589 2585
<< mvnmos >>
rect -9361 1327 -9161 2327
rect -8983 1327 -8783 2327
rect -8605 1327 -8405 2327
rect -8227 1327 -8027 2327
rect -7849 1327 -7649 2327
rect -7471 1327 -7271 2327
rect -7093 1327 -6893 2327
rect -6715 1327 -6515 2327
rect -6337 1327 -6137 2327
rect -5959 1327 -5759 2327
rect -5581 1327 -5381 2327
rect -5203 1327 -5003 2327
rect -4825 1327 -4625 2327
rect -4447 1327 -4247 2327
rect -4069 1327 -3869 2327
rect -3691 1327 -3491 2327
rect -3313 1327 -3113 2327
rect -2935 1327 -2735 2327
rect -2557 1327 -2357 2327
rect -2179 1327 -1979 2327
rect -1801 1327 -1601 2327
rect -1423 1327 -1223 2327
rect -1045 1327 -845 2327
rect -667 1327 -467 2327
rect -289 1327 -89 2327
rect 89 1327 289 2327
rect 467 1327 667 2327
rect 845 1327 1045 2327
rect 1223 1327 1423 2327
rect 1601 1327 1801 2327
rect 1979 1327 2179 2327
rect 2357 1327 2557 2327
rect 2735 1327 2935 2327
rect 3113 1327 3313 2327
rect 3491 1327 3691 2327
rect 3869 1327 4069 2327
rect 4247 1327 4447 2327
rect 4625 1327 4825 2327
rect 5003 1327 5203 2327
rect 5381 1327 5581 2327
rect 5759 1327 5959 2327
rect 6137 1327 6337 2327
rect 6515 1327 6715 2327
rect 6893 1327 7093 2327
rect 7271 1327 7471 2327
rect 7649 1327 7849 2327
rect 8027 1327 8227 2327
rect 8405 1327 8605 2327
rect 8783 1327 8983 2327
rect 9161 1327 9361 2327
rect -9361 109 -9161 1109
rect -8983 109 -8783 1109
rect -8605 109 -8405 1109
rect -8227 109 -8027 1109
rect -7849 109 -7649 1109
rect -7471 109 -7271 1109
rect -7093 109 -6893 1109
rect -6715 109 -6515 1109
rect -6337 109 -6137 1109
rect -5959 109 -5759 1109
rect -5581 109 -5381 1109
rect -5203 109 -5003 1109
rect -4825 109 -4625 1109
rect -4447 109 -4247 1109
rect -4069 109 -3869 1109
rect -3691 109 -3491 1109
rect -3313 109 -3113 1109
rect -2935 109 -2735 1109
rect -2557 109 -2357 1109
rect -2179 109 -1979 1109
rect -1801 109 -1601 1109
rect -1423 109 -1223 1109
rect -1045 109 -845 1109
rect -667 109 -467 1109
rect -289 109 -89 1109
rect 89 109 289 1109
rect 467 109 667 1109
rect 845 109 1045 1109
rect 1223 109 1423 1109
rect 1601 109 1801 1109
rect 1979 109 2179 1109
rect 2357 109 2557 1109
rect 2735 109 2935 1109
rect 3113 109 3313 1109
rect 3491 109 3691 1109
rect 3869 109 4069 1109
rect 4247 109 4447 1109
rect 4625 109 4825 1109
rect 5003 109 5203 1109
rect 5381 109 5581 1109
rect 5759 109 5959 1109
rect 6137 109 6337 1109
rect 6515 109 6715 1109
rect 6893 109 7093 1109
rect 7271 109 7471 1109
rect 7649 109 7849 1109
rect 8027 109 8227 1109
rect 8405 109 8605 1109
rect 8783 109 8983 1109
rect 9161 109 9361 1109
rect -9361 -1109 -9161 -109
rect -8983 -1109 -8783 -109
rect -8605 -1109 -8405 -109
rect -8227 -1109 -8027 -109
rect -7849 -1109 -7649 -109
rect -7471 -1109 -7271 -109
rect -7093 -1109 -6893 -109
rect -6715 -1109 -6515 -109
rect -6337 -1109 -6137 -109
rect -5959 -1109 -5759 -109
rect -5581 -1109 -5381 -109
rect -5203 -1109 -5003 -109
rect -4825 -1109 -4625 -109
rect -4447 -1109 -4247 -109
rect -4069 -1109 -3869 -109
rect -3691 -1109 -3491 -109
rect -3313 -1109 -3113 -109
rect -2935 -1109 -2735 -109
rect -2557 -1109 -2357 -109
rect -2179 -1109 -1979 -109
rect -1801 -1109 -1601 -109
rect -1423 -1109 -1223 -109
rect -1045 -1109 -845 -109
rect -667 -1109 -467 -109
rect -289 -1109 -89 -109
rect 89 -1109 289 -109
rect 467 -1109 667 -109
rect 845 -1109 1045 -109
rect 1223 -1109 1423 -109
rect 1601 -1109 1801 -109
rect 1979 -1109 2179 -109
rect 2357 -1109 2557 -109
rect 2735 -1109 2935 -109
rect 3113 -1109 3313 -109
rect 3491 -1109 3691 -109
rect 3869 -1109 4069 -109
rect 4247 -1109 4447 -109
rect 4625 -1109 4825 -109
rect 5003 -1109 5203 -109
rect 5381 -1109 5581 -109
rect 5759 -1109 5959 -109
rect 6137 -1109 6337 -109
rect 6515 -1109 6715 -109
rect 6893 -1109 7093 -109
rect 7271 -1109 7471 -109
rect 7649 -1109 7849 -109
rect 8027 -1109 8227 -109
rect 8405 -1109 8605 -109
rect 8783 -1109 8983 -109
rect 9161 -1109 9361 -109
rect -9361 -2327 -9161 -1327
rect -8983 -2327 -8783 -1327
rect -8605 -2327 -8405 -1327
rect -8227 -2327 -8027 -1327
rect -7849 -2327 -7649 -1327
rect -7471 -2327 -7271 -1327
rect -7093 -2327 -6893 -1327
rect -6715 -2327 -6515 -1327
rect -6337 -2327 -6137 -1327
rect -5959 -2327 -5759 -1327
rect -5581 -2327 -5381 -1327
rect -5203 -2327 -5003 -1327
rect -4825 -2327 -4625 -1327
rect -4447 -2327 -4247 -1327
rect -4069 -2327 -3869 -1327
rect -3691 -2327 -3491 -1327
rect -3313 -2327 -3113 -1327
rect -2935 -2327 -2735 -1327
rect -2557 -2327 -2357 -1327
rect -2179 -2327 -1979 -1327
rect -1801 -2327 -1601 -1327
rect -1423 -2327 -1223 -1327
rect -1045 -2327 -845 -1327
rect -667 -2327 -467 -1327
rect -289 -2327 -89 -1327
rect 89 -2327 289 -1327
rect 467 -2327 667 -1327
rect 845 -2327 1045 -1327
rect 1223 -2327 1423 -1327
rect 1601 -2327 1801 -1327
rect 1979 -2327 2179 -1327
rect 2357 -2327 2557 -1327
rect 2735 -2327 2935 -1327
rect 3113 -2327 3313 -1327
rect 3491 -2327 3691 -1327
rect 3869 -2327 4069 -1327
rect 4247 -2327 4447 -1327
rect 4625 -2327 4825 -1327
rect 5003 -2327 5203 -1327
rect 5381 -2327 5581 -1327
rect 5759 -2327 5959 -1327
rect 6137 -2327 6337 -1327
rect 6515 -2327 6715 -1327
rect 6893 -2327 7093 -1327
rect 7271 -2327 7471 -1327
rect 7649 -2327 7849 -1327
rect 8027 -2327 8227 -1327
rect 8405 -2327 8605 -1327
rect 8783 -2327 8983 -1327
rect 9161 -2327 9361 -1327
<< mvndiff >>
rect -9419 2315 -9361 2327
rect -9419 1339 -9407 2315
rect -9373 1339 -9361 2315
rect -9419 1327 -9361 1339
rect -9161 2315 -9103 2327
rect -9161 1339 -9149 2315
rect -9115 1339 -9103 2315
rect -9161 1327 -9103 1339
rect -9041 2315 -8983 2327
rect -9041 1339 -9029 2315
rect -8995 1339 -8983 2315
rect -9041 1327 -8983 1339
rect -8783 2315 -8725 2327
rect -8783 1339 -8771 2315
rect -8737 1339 -8725 2315
rect -8783 1327 -8725 1339
rect -8663 2315 -8605 2327
rect -8663 1339 -8651 2315
rect -8617 1339 -8605 2315
rect -8663 1327 -8605 1339
rect -8405 2315 -8347 2327
rect -8405 1339 -8393 2315
rect -8359 1339 -8347 2315
rect -8405 1327 -8347 1339
rect -8285 2315 -8227 2327
rect -8285 1339 -8273 2315
rect -8239 1339 -8227 2315
rect -8285 1327 -8227 1339
rect -8027 2315 -7969 2327
rect -8027 1339 -8015 2315
rect -7981 1339 -7969 2315
rect -8027 1327 -7969 1339
rect -7907 2315 -7849 2327
rect -7907 1339 -7895 2315
rect -7861 1339 -7849 2315
rect -7907 1327 -7849 1339
rect -7649 2315 -7591 2327
rect -7649 1339 -7637 2315
rect -7603 1339 -7591 2315
rect -7649 1327 -7591 1339
rect -7529 2315 -7471 2327
rect -7529 1339 -7517 2315
rect -7483 1339 -7471 2315
rect -7529 1327 -7471 1339
rect -7271 2315 -7213 2327
rect -7271 1339 -7259 2315
rect -7225 1339 -7213 2315
rect -7271 1327 -7213 1339
rect -7151 2315 -7093 2327
rect -7151 1339 -7139 2315
rect -7105 1339 -7093 2315
rect -7151 1327 -7093 1339
rect -6893 2315 -6835 2327
rect -6893 1339 -6881 2315
rect -6847 1339 -6835 2315
rect -6893 1327 -6835 1339
rect -6773 2315 -6715 2327
rect -6773 1339 -6761 2315
rect -6727 1339 -6715 2315
rect -6773 1327 -6715 1339
rect -6515 2315 -6457 2327
rect -6515 1339 -6503 2315
rect -6469 1339 -6457 2315
rect -6515 1327 -6457 1339
rect -6395 2315 -6337 2327
rect -6395 1339 -6383 2315
rect -6349 1339 -6337 2315
rect -6395 1327 -6337 1339
rect -6137 2315 -6079 2327
rect -6137 1339 -6125 2315
rect -6091 1339 -6079 2315
rect -6137 1327 -6079 1339
rect -6017 2315 -5959 2327
rect -6017 1339 -6005 2315
rect -5971 1339 -5959 2315
rect -6017 1327 -5959 1339
rect -5759 2315 -5701 2327
rect -5759 1339 -5747 2315
rect -5713 1339 -5701 2315
rect -5759 1327 -5701 1339
rect -5639 2315 -5581 2327
rect -5639 1339 -5627 2315
rect -5593 1339 -5581 2315
rect -5639 1327 -5581 1339
rect -5381 2315 -5323 2327
rect -5381 1339 -5369 2315
rect -5335 1339 -5323 2315
rect -5381 1327 -5323 1339
rect -5261 2315 -5203 2327
rect -5261 1339 -5249 2315
rect -5215 1339 -5203 2315
rect -5261 1327 -5203 1339
rect -5003 2315 -4945 2327
rect -5003 1339 -4991 2315
rect -4957 1339 -4945 2315
rect -5003 1327 -4945 1339
rect -4883 2315 -4825 2327
rect -4883 1339 -4871 2315
rect -4837 1339 -4825 2315
rect -4883 1327 -4825 1339
rect -4625 2315 -4567 2327
rect -4625 1339 -4613 2315
rect -4579 1339 -4567 2315
rect -4625 1327 -4567 1339
rect -4505 2315 -4447 2327
rect -4505 1339 -4493 2315
rect -4459 1339 -4447 2315
rect -4505 1327 -4447 1339
rect -4247 2315 -4189 2327
rect -4247 1339 -4235 2315
rect -4201 1339 -4189 2315
rect -4247 1327 -4189 1339
rect -4127 2315 -4069 2327
rect -4127 1339 -4115 2315
rect -4081 1339 -4069 2315
rect -4127 1327 -4069 1339
rect -3869 2315 -3811 2327
rect -3869 1339 -3857 2315
rect -3823 1339 -3811 2315
rect -3869 1327 -3811 1339
rect -3749 2315 -3691 2327
rect -3749 1339 -3737 2315
rect -3703 1339 -3691 2315
rect -3749 1327 -3691 1339
rect -3491 2315 -3433 2327
rect -3491 1339 -3479 2315
rect -3445 1339 -3433 2315
rect -3491 1327 -3433 1339
rect -3371 2315 -3313 2327
rect -3371 1339 -3359 2315
rect -3325 1339 -3313 2315
rect -3371 1327 -3313 1339
rect -3113 2315 -3055 2327
rect -3113 1339 -3101 2315
rect -3067 1339 -3055 2315
rect -3113 1327 -3055 1339
rect -2993 2315 -2935 2327
rect -2993 1339 -2981 2315
rect -2947 1339 -2935 2315
rect -2993 1327 -2935 1339
rect -2735 2315 -2677 2327
rect -2735 1339 -2723 2315
rect -2689 1339 -2677 2315
rect -2735 1327 -2677 1339
rect -2615 2315 -2557 2327
rect -2615 1339 -2603 2315
rect -2569 1339 -2557 2315
rect -2615 1327 -2557 1339
rect -2357 2315 -2299 2327
rect -2357 1339 -2345 2315
rect -2311 1339 -2299 2315
rect -2357 1327 -2299 1339
rect -2237 2315 -2179 2327
rect -2237 1339 -2225 2315
rect -2191 1339 -2179 2315
rect -2237 1327 -2179 1339
rect -1979 2315 -1921 2327
rect -1979 1339 -1967 2315
rect -1933 1339 -1921 2315
rect -1979 1327 -1921 1339
rect -1859 2315 -1801 2327
rect -1859 1339 -1847 2315
rect -1813 1339 -1801 2315
rect -1859 1327 -1801 1339
rect -1601 2315 -1543 2327
rect -1601 1339 -1589 2315
rect -1555 1339 -1543 2315
rect -1601 1327 -1543 1339
rect -1481 2315 -1423 2327
rect -1481 1339 -1469 2315
rect -1435 1339 -1423 2315
rect -1481 1327 -1423 1339
rect -1223 2315 -1165 2327
rect -1223 1339 -1211 2315
rect -1177 1339 -1165 2315
rect -1223 1327 -1165 1339
rect -1103 2315 -1045 2327
rect -1103 1339 -1091 2315
rect -1057 1339 -1045 2315
rect -1103 1327 -1045 1339
rect -845 2315 -787 2327
rect -845 1339 -833 2315
rect -799 1339 -787 2315
rect -845 1327 -787 1339
rect -725 2315 -667 2327
rect -725 1339 -713 2315
rect -679 1339 -667 2315
rect -725 1327 -667 1339
rect -467 2315 -409 2327
rect -467 1339 -455 2315
rect -421 1339 -409 2315
rect -467 1327 -409 1339
rect -347 2315 -289 2327
rect -347 1339 -335 2315
rect -301 1339 -289 2315
rect -347 1327 -289 1339
rect -89 2315 -31 2327
rect -89 1339 -77 2315
rect -43 1339 -31 2315
rect -89 1327 -31 1339
rect 31 2315 89 2327
rect 31 1339 43 2315
rect 77 1339 89 2315
rect 31 1327 89 1339
rect 289 2315 347 2327
rect 289 1339 301 2315
rect 335 1339 347 2315
rect 289 1327 347 1339
rect 409 2315 467 2327
rect 409 1339 421 2315
rect 455 1339 467 2315
rect 409 1327 467 1339
rect 667 2315 725 2327
rect 667 1339 679 2315
rect 713 1339 725 2315
rect 667 1327 725 1339
rect 787 2315 845 2327
rect 787 1339 799 2315
rect 833 1339 845 2315
rect 787 1327 845 1339
rect 1045 2315 1103 2327
rect 1045 1339 1057 2315
rect 1091 1339 1103 2315
rect 1045 1327 1103 1339
rect 1165 2315 1223 2327
rect 1165 1339 1177 2315
rect 1211 1339 1223 2315
rect 1165 1327 1223 1339
rect 1423 2315 1481 2327
rect 1423 1339 1435 2315
rect 1469 1339 1481 2315
rect 1423 1327 1481 1339
rect 1543 2315 1601 2327
rect 1543 1339 1555 2315
rect 1589 1339 1601 2315
rect 1543 1327 1601 1339
rect 1801 2315 1859 2327
rect 1801 1339 1813 2315
rect 1847 1339 1859 2315
rect 1801 1327 1859 1339
rect 1921 2315 1979 2327
rect 1921 1339 1933 2315
rect 1967 1339 1979 2315
rect 1921 1327 1979 1339
rect 2179 2315 2237 2327
rect 2179 1339 2191 2315
rect 2225 1339 2237 2315
rect 2179 1327 2237 1339
rect 2299 2315 2357 2327
rect 2299 1339 2311 2315
rect 2345 1339 2357 2315
rect 2299 1327 2357 1339
rect 2557 2315 2615 2327
rect 2557 1339 2569 2315
rect 2603 1339 2615 2315
rect 2557 1327 2615 1339
rect 2677 2315 2735 2327
rect 2677 1339 2689 2315
rect 2723 1339 2735 2315
rect 2677 1327 2735 1339
rect 2935 2315 2993 2327
rect 2935 1339 2947 2315
rect 2981 1339 2993 2315
rect 2935 1327 2993 1339
rect 3055 2315 3113 2327
rect 3055 1339 3067 2315
rect 3101 1339 3113 2315
rect 3055 1327 3113 1339
rect 3313 2315 3371 2327
rect 3313 1339 3325 2315
rect 3359 1339 3371 2315
rect 3313 1327 3371 1339
rect 3433 2315 3491 2327
rect 3433 1339 3445 2315
rect 3479 1339 3491 2315
rect 3433 1327 3491 1339
rect 3691 2315 3749 2327
rect 3691 1339 3703 2315
rect 3737 1339 3749 2315
rect 3691 1327 3749 1339
rect 3811 2315 3869 2327
rect 3811 1339 3823 2315
rect 3857 1339 3869 2315
rect 3811 1327 3869 1339
rect 4069 2315 4127 2327
rect 4069 1339 4081 2315
rect 4115 1339 4127 2315
rect 4069 1327 4127 1339
rect 4189 2315 4247 2327
rect 4189 1339 4201 2315
rect 4235 1339 4247 2315
rect 4189 1327 4247 1339
rect 4447 2315 4505 2327
rect 4447 1339 4459 2315
rect 4493 1339 4505 2315
rect 4447 1327 4505 1339
rect 4567 2315 4625 2327
rect 4567 1339 4579 2315
rect 4613 1339 4625 2315
rect 4567 1327 4625 1339
rect 4825 2315 4883 2327
rect 4825 1339 4837 2315
rect 4871 1339 4883 2315
rect 4825 1327 4883 1339
rect 4945 2315 5003 2327
rect 4945 1339 4957 2315
rect 4991 1339 5003 2315
rect 4945 1327 5003 1339
rect 5203 2315 5261 2327
rect 5203 1339 5215 2315
rect 5249 1339 5261 2315
rect 5203 1327 5261 1339
rect 5323 2315 5381 2327
rect 5323 1339 5335 2315
rect 5369 1339 5381 2315
rect 5323 1327 5381 1339
rect 5581 2315 5639 2327
rect 5581 1339 5593 2315
rect 5627 1339 5639 2315
rect 5581 1327 5639 1339
rect 5701 2315 5759 2327
rect 5701 1339 5713 2315
rect 5747 1339 5759 2315
rect 5701 1327 5759 1339
rect 5959 2315 6017 2327
rect 5959 1339 5971 2315
rect 6005 1339 6017 2315
rect 5959 1327 6017 1339
rect 6079 2315 6137 2327
rect 6079 1339 6091 2315
rect 6125 1339 6137 2315
rect 6079 1327 6137 1339
rect 6337 2315 6395 2327
rect 6337 1339 6349 2315
rect 6383 1339 6395 2315
rect 6337 1327 6395 1339
rect 6457 2315 6515 2327
rect 6457 1339 6469 2315
rect 6503 1339 6515 2315
rect 6457 1327 6515 1339
rect 6715 2315 6773 2327
rect 6715 1339 6727 2315
rect 6761 1339 6773 2315
rect 6715 1327 6773 1339
rect 6835 2315 6893 2327
rect 6835 1339 6847 2315
rect 6881 1339 6893 2315
rect 6835 1327 6893 1339
rect 7093 2315 7151 2327
rect 7093 1339 7105 2315
rect 7139 1339 7151 2315
rect 7093 1327 7151 1339
rect 7213 2315 7271 2327
rect 7213 1339 7225 2315
rect 7259 1339 7271 2315
rect 7213 1327 7271 1339
rect 7471 2315 7529 2327
rect 7471 1339 7483 2315
rect 7517 1339 7529 2315
rect 7471 1327 7529 1339
rect 7591 2315 7649 2327
rect 7591 1339 7603 2315
rect 7637 1339 7649 2315
rect 7591 1327 7649 1339
rect 7849 2315 7907 2327
rect 7849 1339 7861 2315
rect 7895 1339 7907 2315
rect 7849 1327 7907 1339
rect 7969 2315 8027 2327
rect 7969 1339 7981 2315
rect 8015 1339 8027 2315
rect 7969 1327 8027 1339
rect 8227 2315 8285 2327
rect 8227 1339 8239 2315
rect 8273 1339 8285 2315
rect 8227 1327 8285 1339
rect 8347 2315 8405 2327
rect 8347 1339 8359 2315
rect 8393 1339 8405 2315
rect 8347 1327 8405 1339
rect 8605 2315 8663 2327
rect 8605 1339 8617 2315
rect 8651 1339 8663 2315
rect 8605 1327 8663 1339
rect 8725 2315 8783 2327
rect 8725 1339 8737 2315
rect 8771 1339 8783 2315
rect 8725 1327 8783 1339
rect 8983 2315 9041 2327
rect 8983 1339 8995 2315
rect 9029 1339 9041 2315
rect 8983 1327 9041 1339
rect 9103 2315 9161 2327
rect 9103 1339 9115 2315
rect 9149 1339 9161 2315
rect 9103 1327 9161 1339
rect 9361 2315 9419 2327
rect 9361 1339 9373 2315
rect 9407 1339 9419 2315
rect 9361 1327 9419 1339
rect -9419 1097 -9361 1109
rect -9419 121 -9407 1097
rect -9373 121 -9361 1097
rect -9419 109 -9361 121
rect -9161 1097 -9103 1109
rect -9161 121 -9149 1097
rect -9115 121 -9103 1097
rect -9161 109 -9103 121
rect -9041 1097 -8983 1109
rect -9041 121 -9029 1097
rect -8995 121 -8983 1097
rect -9041 109 -8983 121
rect -8783 1097 -8725 1109
rect -8783 121 -8771 1097
rect -8737 121 -8725 1097
rect -8783 109 -8725 121
rect -8663 1097 -8605 1109
rect -8663 121 -8651 1097
rect -8617 121 -8605 1097
rect -8663 109 -8605 121
rect -8405 1097 -8347 1109
rect -8405 121 -8393 1097
rect -8359 121 -8347 1097
rect -8405 109 -8347 121
rect -8285 1097 -8227 1109
rect -8285 121 -8273 1097
rect -8239 121 -8227 1097
rect -8285 109 -8227 121
rect -8027 1097 -7969 1109
rect -8027 121 -8015 1097
rect -7981 121 -7969 1097
rect -8027 109 -7969 121
rect -7907 1097 -7849 1109
rect -7907 121 -7895 1097
rect -7861 121 -7849 1097
rect -7907 109 -7849 121
rect -7649 1097 -7591 1109
rect -7649 121 -7637 1097
rect -7603 121 -7591 1097
rect -7649 109 -7591 121
rect -7529 1097 -7471 1109
rect -7529 121 -7517 1097
rect -7483 121 -7471 1097
rect -7529 109 -7471 121
rect -7271 1097 -7213 1109
rect -7271 121 -7259 1097
rect -7225 121 -7213 1097
rect -7271 109 -7213 121
rect -7151 1097 -7093 1109
rect -7151 121 -7139 1097
rect -7105 121 -7093 1097
rect -7151 109 -7093 121
rect -6893 1097 -6835 1109
rect -6893 121 -6881 1097
rect -6847 121 -6835 1097
rect -6893 109 -6835 121
rect -6773 1097 -6715 1109
rect -6773 121 -6761 1097
rect -6727 121 -6715 1097
rect -6773 109 -6715 121
rect -6515 1097 -6457 1109
rect -6515 121 -6503 1097
rect -6469 121 -6457 1097
rect -6515 109 -6457 121
rect -6395 1097 -6337 1109
rect -6395 121 -6383 1097
rect -6349 121 -6337 1097
rect -6395 109 -6337 121
rect -6137 1097 -6079 1109
rect -6137 121 -6125 1097
rect -6091 121 -6079 1097
rect -6137 109 -6079 121
rect -6017 1097 -5959 1109
rect -6017 121 -6005 1097
rect -5971 121 -5959 1097
rect -6017 109 -5959 121
rect -5759 1097 -5701 1109
rect -5759 121 -5747 1097
rect -5713 121 -5701 1097
rect -5759 109 -5701 121
rect -5639 1097 -5581 1109
rect -5639 121 -5627 1097
rect -5593 121 -5581 1097
rect -5639 109 -5581 121
rect -5381 1097 -5323 1109
rect -5381 121 -5369 1097
rect -5335 121 -5323 1097
rect -5381 109 -5323 121
rect -5261 1097 -5203 1109
rect -5261 121 -5249 1097
rect -5215 121 -5203 1097
rect -5261 109 -5203 121
rect -5003 1097 -4945 1109
rect -5003 121 -4991 1097
rect -4957 121 -4945 1097
rect -5003 109 -4945 121
rect -4883 1097 -4825 1109
rect -4883 121 -4871 1097
rect -4837 121 -4825 1097
rect -4883 109 -4825 121
rect -4625 1097 -4567 1109
rect -4625 121 -4613 1097
rect -4579 121 -4567 1097
rect -4625 109 -4567 121
rect -4505 1097 -4447 1109
rect -4505 121 -4493 1097
rect -4459 121 -4447 1097
rect -4505 109 -4447 121
rect -4247 1097 -4189 1109
rect -4247 121 -4235 1097
rect -4201 121 -4189 1097
rect -4247 109 -4189 121
rect -4127 1097 -4069 1109
rect -4127 121 -4115 1097
rect -4081 121 -4069 1097
rect -4127 109 -4069 121
rect -3869 1097 -3811 1109
rect -3869 121 -3857 1097
rect -3823 121 -3811 1097
rect -3869 109 -3811 121
rect -3749 1097 -3691 1109
rect -3749 121 -3737 1097
rect -3703 121 -3691 1097
rect -3749 109 -3691 121
rect -3491 1097 -3433 1109
rect -3491 121 -3479 1097
rect -3445 121 -3433 1097
rect -3491 109 -3433 121
rect -3371 1097 -3313 1109
rect -3371 121 -3359 1097
rect -3325 121 -3313 1097
rect -3371 109 -3313 121
rect -3113 1097 -3055 1109
rect -3113 121 -3101 1097
rect -3067 121 -3055 1097
rect -3113 109 -3055 121
rect -2993 1097 -2935 1109
rect -2993 121 -2981 1097
rect -2947 121 -2935 1097
rect -2993 109 -2935 121
rect -2735 1097 -2677 1109
rect -2735 121 -2723 1097
rect -2689 121 -2677 1097
rect -2735 109 -2677 121
rect -2615 1097 -2557 1109
rect -2615 121 -2603 1097
rect -2569 121 -2557 1097
rect -2615 109 -2557 121
rect -2357 1097 -2299 1109
rect -2357 121 -2345 1097
rect -2311 121 -2299 1097
rect -2357 109 -2299 121
rect -2237 1097 -2179 1109
rect -2237 121 -2225 1097
rect -2191 121 -2179 1097
rect -2237 109 -2179 121
rect -1979 1097 -1921 1109
rect -1979 121 -1967 1097
rect -1933 121 -1921 1097
rect -1979 109 -1921 121
rect -1859 1097 -1801 1109
rect -1859 121 -1847 1097
rect -1813 121 -1801 1097
rect -1859 109 -1801 121
rect -1601 1097 -1543 1109
rect -1601 121 -1589 1097
rect -1555 121 -1543 1097
rect -1601 109 -1543 121
rect -1481 1097 -1423 1109
rect -1481 121 -1469 1097
rect -1435 121 -1423 1097
rect -1481 109 -1423 121
rect -1223 1097 -1165 1109
rect -1223 121 -1211 1097
rect -1177 121 -1165 1097
rect -1223 109 -1165 121
rect -1103 1097 -1045 1109
rect -1103 121 -1091 1097
rect -1057 121 -1045 1097
rect -1103 109 -1045 121
rect -845 1097 -787 1109
rect -845 121 -833 1097
rect -799 121 -787 1097
rect -845 109 -787 121
rect -725 1097 -667 1109
rect -725 121 -713 1097
rect -679 121 -667 1097
rect -725 109 -667 121
rect -467 1097 -409 1109
rect -467 121 -455 1097
rect -421 121 -409 1097
rect -467 109 -409 121
rect -347 1097 -289 1109
rect -347 121 -335 1097
rect -301 121 -289 1097
rect -347 109 -289 121
rect -89 1097 -31 1109
rect -89 121 -77 1097
rect -43 121 -31 1097
rect -89 109 -31 121
rect 31 1097 89 1109
rect 31 121 43 1097
rect 77 121 89 1097
rect 31 109 89 121
rect 289 1097 347 1109
rect 289 121 301 1097
rect 335 121 347 1097
rect 289 109 347 121
rect 409 1097 467 1109
rect 409 121 421 1097
rect 455 121 467 1097
rect 409 109 467 121
rect 667 1097 725 1109
rect 667 121 679 1097
rect 713 121 725 1097
rect 667 109 725 121
rect 787 1097 845 1109
rect 787 121 799 1097
rect 833 121 845 1097
rect 787 109 845 121
rect 1045 1097 1103 1109
rect 1045 121 1057 1097
rect 1091 121 1103 1097
rect 1045 109 1103 121
rect 1165 1097 1223 1109
rect 1165 121 1177 1097
rect 1211 121 1223 1097
rect 1165 109 1223 121
rect 1423 1097 1481 1109
rect 1423 121 1435 1097
rect 1469 121 1481 1097
rect 1423 109 1481 121
rect 1543 1097 1601 1109
rect 1543 121 1555 1097
rect 1589 121 1601 1097
rect 1543 109 1601 121
rect 1801 1097 1859 1109
rect 1801 121 1813 1097
rect 1847 121 1859 1097
rect 1801 109 1859 121
rect 1921 1097 1979 1109
rect 1921 121 1933 1097
rect 1967 121 1979 1097
rect 1921 109 1979 121
rect 2179 1097 2237 1109
rect 2179 121 2191 1097
rect 2225 121 2237 1097
rect 2179 109 2237 121
rect 2299 1097 2357 1109
rect 2299 121 2311 1097
rect 2345 121 2357 1097
rect 2299 109 2357 121
rect 2557 1097 2615 1109
rect 2557 121 2569 1097
rect 2603 121 2615 1097
rect 2557 109 2615 121
rect 2677 1097 2735 1109
rect 2677 121 2689 1097
rect 2723 121 2735 1097
rect 2677 109 2735 121
rect 2935 1097 2993 1109
rect 2935 121 2947 1097
rect 2981 121 2993 1097
rect 2935 109 2993 121
rect 3055 1097 3113 1109
rect 3055 121 3067 1097
rect 3101 121 3113 1097
rect 3055 109 3113 121
rect 3313 1097 3371 1109
rect 3313 121 3325 1097
rect 3359 121 3371 1097
rect 3313 109 3371 121
rect 3433 1097 3491 1109
rect 3433 121 3445 1097
rect 3479 121 3491 1097
rect 3433 109 3491 121
rect 3691 1097 3749 1109
rect 3691 121 3703 1097
rect 3737 121 3749 1097
rect 3691 109 3749 121
rect 3811 1097 3869 1109
rect 3811 121 3823 1097
rect 3857 121 3869 1097
rect 3811 109 3869 121
rect 4069 1097 4127 1109
rect 4069 121 4081 1097
rect 4115 121 4127 1097
rect 4069 109 4127 121
rect 4189 1097 4247 1109
rect 4189 121 4201 1097
rect 4235 121 4247 1097
rect 4189 109 4247 121
rect 4447 1097 4505 1109
rect 4447 121 4459 1097
rect 4493 121 4505 1097
rect 4447 109 4505 121
rect 4567 1097 4625 1109
rect 4567 121 4579 1097
rect 4613 121 4625 1097
rect 4567 109 4625 121
rect 4825 1097 4883 1109
rect 4825 121 4837 1097
rect 4871 121 4883 1097
rect 4825 109 4883 121
rect 4945 1097 5003 1109
rect 4945 121 4957 1097
rect 4991 121 5003 1097
rect 4945 109 5003 121
rect 5203 1097 5261 1109
rect 5203 121 5215 1097
rect 5249 121 5261 1097
rect 5203 109 5261 121
rect 5323 1097 5381 1109
rect 5323 121 5335 1097
rect 5369 121 5381 1097
rect 5323 109 5381 121
rect 5581 1097 5639 1109
rect 5581 121 5593 1097
rect 5627 121 5639 1097
rect 5581 109 5639 121
rect 5701 1097 5759 1109
rect 5701 121 5713 1097
rect 5747 121 5759 1097
rect 5701 109 5759 121
rect 5959 1097 6017 1109
rect 5959 121 5971 1097
rect 6005 121 6017 1097
rect 5959 109 6017 121
rect 6079 1097 6137 1109
rect 6079 121 6091 1097
rect 6125 121 6137 1097
rect 6079 109 6137 121
rect 6337 1097 6395 1109
rect 6337 121 6349 1097
rect 6383 121 6395 1097
rect 6337 109 6395 121
rect 6457 1097 6515 1109
rect 6457 121 6469 1097
rect 6503 121 6515 1097
rect 6457 109 6515 121
rect 6715 1097 6773 1109
rect 6715 121 6727 1097
rect 6761 121 6773 1097
rect 6715 109 6773 121
rect 6835 1097 6893 1109
rect 6835 121 6847 1097
rect 6881 121 6893 1097
rect 6835 109 6893 121
rect 7093 1097 7151 1109
rect 7093 121 7105 1097
rect 7139 121 7151 1097
rect 7093 109 7151 121
rect 7213 1097 7271 1109
rect 7213 121 7225 1097
rect 7259 121 7271 1097
rect 7213 109 7271 121
rect 7471 1097 7529 1109
rect 7471 121 7483 1097
rect 7517 121 7529 1097
rect 7471 109 7529 121
rect 7591 1097 7649 1109
rect 7591 121 7603 1097
rect 7637 121 7649 1097
rect 7591 109 7649 121
rect 7849 1097 7907 1109
rect 7849 121 7861 1097
rect 7895 121 7907 1097
rect 7849 109 7907 121
rect 7969 1097 8027 1109
rect 7969 121 7981 1097
rect 8015 121 8027 1097
rect 7969 109 8027 121
rect 8227 1097 8285 1109
rect 8227 121 8239 1097
rect 8273 121 8285 1097
rect 8227 109 8285 121
rect 8347 1097 8405 1109
rect 8347 121 8359 1097
rect 8393 121 8405 1097
rect 8347 109 8405 121
rect 8605 1097 8663 1109
rect 8605 121 8617 1097
rect 8651 121 8663 1097
rect 8605 109 8663 121
rect 8725 1097 8783 1109
rect 8725 121 8737 1097
rect 8771 121 8783 1097
rect 8725 109 8783 121
rect 8983 1097 9041 1109
rect 8983 121 8995 1097
rect 9029 121 9041 1097
rect 8983 109 9041 121
rect 9103 1097 9161 1109
rect 9103 121 9115 1097
rect 9149 121 9161 1097
rect 9103 109 9161 121
rect 9361 1097 9419 1109
rect 9361 121 9373 1097
rect 9407 121 9419 1097
rect 9361 109 9419 121
rect -9419 -121 -9361 -109
rect -9419 -1097 -9407 -121
rect -9373 -1097 -9361 -121
rect -9419 -1109 -9361 -1097
rect -9161 -121 -9103 -109
rect -9161 -1097 -9149 -121
rect -9115 -1097 -9103 -121
rect -9161 -1109 -9103 -1097
rect -9041 -121 -8983 -109
rect -9041 -1097 -9029 -121
rect -8995 -1097 -8983 -121
rect -9041 -1109 -8983 -1097
rect -8783 -121 -8725 -109
rect -8783 -1097 -8771 -121
rect -8737 -1097 -8725 -121
rect -8783 -1109 -8725 -1097
rect -8663 -121 -8605 -109
rect -8663 -1097 -8651 -121
rect -8617 -1097 -8605 -121
rect -8663 -1109 -8605 -1097
rect -8405 -121 -8347 -109
rect -8405 -1097 -8393 -121
rect -8359 -1097 -8347 -121
rect -8405 -1109 -8347 -1097
rect -8285 -121 -8227 -109
rect -8285 -1097 -8273 -121
rect -8239 -1097 -8227 -121
rect -8285 -1109 -8227 -1097
rect -8027 -121 -7969 -109
rect -8027 -1097 -8015 -121
rect -7981 -1097 -7969 -121
rect -8027 -1109 -7969 -1097
rect -7907 -121 -7849 -109
rect -7907 -1097 -7895 -121
rect -7861 -1097 -7849 -121
rect -7907 -1109 -7849 -1097
rect -7649 -121 -7591 -109
rect -7649 -1097 -7637 -121
rect -7603 -1097 -7591 -121
rect -7649 -1109 -7591 -1097
rect -7529 -121 -7471 -109
rect -7529 -1097 -7517 -121
rect -7483 -1097 -7471 -121
rect -7529 -1109 -7471 -1097
rect -7271 -121 -7213 -109
rect -7271 -1097 -7259 -121
rect -7225 -1097 -7213 -121
rect -7271 -1109 -7213 -1097
rect -7151 -121 -7093 -109
rect -7151 -1097 -7139 -121
rect -7105 -1097 -7093 -121
rect -7151 -1109 -7093 -1097
rect -6893 -121 -6835 -109
rect -6893 -1097 -6881 -121
rect -6847 -1097 -6835 -121
rect -6893 -1109 -6835 -1097
rect -6773 -121 -6715 -109
rect -6773 -1097 -6761 -121
rect -6727 -1097 -6715 -121
rect -6773 -1109 -6715 -1097
rect -6515 -121 -6457 -109
rect -6515 -1097 -6503 -121
rect -6469 -1097 -6457 -121
rect -6515 -1109 -6457 -1097
rect -6395 -121 -6337 -109
rect -6395 -1097 -6383 -121
rect -6349 -1097 -6337 -121
rect -6395 -1109 -6337 -1097
rect -6137 -121 -6079 -109
rect -6137 -1097 -6125 -121
rect -6091 -1097 -6079 -121
rect -6137 -1109 -6079 -1097
rect -6017 -121 -5959 -109
rect -6017 -1097 -6005 -121
rect -5971 -1097 -5959 -121
rect -6017 -1109 -5959 -1097
rect -5759 -121 -5701 -109
rect -5759 -1097 -5747 -121
rect -5713 -1097 -5701 -121
rect -5759 -1109 -5701 -1097
rect -5639 -121 -5581 -109
rect -5639 -1097 -5627 -121
rect -5593 -1097 -5581 -121
rect -5639 -1109 -5581 -1097
rect -5381 -121 -5323 -109
rect -5381 -1097 -5369 -121
rect -5335 -1097 -5323 -121
rect -5381 -1109 -5323 -1097
rect -5261 -121 -5203 -109
rect -5261 -1097 -5249 -121
rect -5215 -1097 -5203 -121
rect -5261 -1109 -5203 -1097
rect -5003 -121 -4945 -109
rect -5003 -1097 -4991 -121
rect -4957 -1097 -4945 -121
rect -5003 -1109 -4945 -1097
rect -4883 -121 -4825 -109
rect -4883 -1097 -4871 -121
rect -4837 -1097 -4825 -121
rect -4883 -1109 -4825 -1097
rect -4625 -121 -4567 -109
rect -4625 -1097 -4613 -121
rect -4579 -1097 -4567 -121
rect -4625 -1109 -4567 -1097
rect -4505 -121 -4447 -109
rect -4505 -1097 -4493 -121
rect -4459 -1097 -4447 -121
rect -4505 -1109 -4447 -1097
rect -4247 -121 -4189 -109
rect -4247 -1097 -4235 -121
rect -4201 -1097 -4189 -121
rect -4247 -1109 -4189 -1097
rect -4127 -121 -4069 -109
rect -4127 -1097 -4115 -121
rect -4081 -1097 -4069 -121
rect -4127 -1109 -4069 -1097
rect -3869 -121 -3811 -109
rect -3869 -1097 -3857 -121
rect -3823 -1097 -3811 -121
rect -3869 -1109 -3811 -1097
rect -3749 -121 -3691 -109
rect -3749 -1097 -3737 -121
rect -3703 -1097 -3691 -121
rect -3749 -1109 -3691 -1097
rect -3491 -121 -3433 -109
rect -3491 -1097 -3479 -121
rect -3445 -1097 -3433 -121
rect -3491 -1109 -3433 -1097
rect -3371 -121 -3313 -109
rect -3371 -1097 -3359 -121
rect -3325 -1097 -3313 -121
rect -3371 -1109 -3313 -1097
rect -3113 -121 -3055 -109
rect -3113 -1097 -3101 -121
rect -3067 -1097 -3055 -121
rect -3113 -1109 -3055 -1097
rect -2993 -121 -2935 -109
rect -2993 -1097 -2981 -121
rect -2947 -1097 -2935 -121
rect -2993 -1109 -2935 -1097
rect -2735 -121 -2677 -109
rect -2735 -1097 -2723 -121
rect -2689 -1097 -2677 -121
rect -2735 -1109 -2677 -1097
rect -2615 -121 -2557 -109
rect -2615 -1097 -2603 -121
rect -2569 -1097 -2557 -121
rect -2615 -1109 -2557 -1097
rect -2357 -121 -2299 -109
rect -2357 -1097 -2345 -121
rect -2311 -1097 -2299 -121
rect -2357 -1109 -2299 -1097
rect -2237 -121 -2179 -109
rect -2237 -1097 -2225 -121
rect -2191 -1097 -2179 -121
rect -2237 -1109 -2179 -1097
rect -1979 -121 -1921 -109
rect -1979 -1097 -1967 -121
rect -1933 -1097 -1921 -121
rect -1979 -1109 -1921 -1097
rect -1859 -121 -1801 -109
rect -1859 -1097 -1847 -121
rect -1813 -1097 -1801 -121
rect -1859 -1109 -1801 -1097
rect -1601 -121 -1543 -109
rect -1601 -1097 -1589 -121
rect -1555 -1097 -1543 -121
rect -1601 -1109 -1543 -1097
rect -1481 -121 -1423 -109
rect -1481 -1097 -1469 -121
rect -1435 -1097 -1423 -121
rect -1481 -1109 -1423 -1097
rect -1223 -121 -1165 -109
rect -1223 -1097 -1211 -121
rect -1177 -1097 -1165 -121
rect -1223 -1109 -1165 -1097
rect -1103 -121 -1045 -109
rect -1103 -1097 -1091 -121
rect -1057 -1097 -1045 -121
rect -1103 -1109 -1045 -1097
rect -845 -121 -787 -109
rect -845 -1097 -833 -121
rect -799 -1097 -787 -121
rect -845 -1109 -787 -1097
rect -725 -121 -667 -109
rect -725 -1097 -713 -121
rect -679 -1097 -667 -121
rect -725 -1109 -667 -1097
rect -467 -121 -409 -109
rect -467 -1097 -455 -121
rect -421 -1097 -409 -121
rect -467 -1109 -409 -1097
rect -347 -121 -289 -109
rect -347 -1097 -335 -121
rect -301 -1097 -289 -121
rect -347 -1109 -289 -1097
rect -89 -121 -31 -109
rect -89 -1097 -77 -121
rect -43 -1097 -31 -121
rect -89 -1109 -31 -1097
rect 31 -121 89 -109
rect 31 -1097 43 -121
rect 77 -1097 89 -121
rect 31 -1109 89 -1097
rect 289 -121 347 -109
rect 289 -1097 301 -121
rect 335 -1097 347 -121
rect 289 -1109 347 -1097
rect 409 -121 467 -109
rect 409 -1097 421 -121
rect 455 -1097 467 -121
rect 409 -1109 467 -1097
rect 667 -121 725 -109
rect 667 -1097 679 -121
rect 713 -1097 725 -121
rect 667 -1109 725 -1097
rect 787 -121 845 -109
rect 787 -1097 799 -121
rect 833 -1097 845 -121
rect 787 -1109 845 -1097
rect 1045 -121 1103 -109
rect 1045 -1097 1057 -121
rect 1091 -1097 1103 -121
rect 1045 -1109 1103 -1097
rect 1165 -121 1223 -109
rect 1165 -1097 1177 -121
rect 1211 -1097 1223 -121
rect 1165 -1109 1223 -1097
rect 1423 -121 1481 -109
rect 1423 -1097 1435 -121
rect 1469 -1097 1481 -121
rect 1423 -1109 1481 -1097
rect 1543 -121 1601 -109
rect 1543 -1097 1555 -121
rect 1589 -1097 1601 -121
rect 1543 -1109 1601 -1097
rect 1801 -121 1859 -109
rect 1801 -1097 1813 -121
rect 1847 -1097 1859 -121
rect 1801 -1109 1859 -1097
rect 1921 -121 1979 -109
rect 1921 -1097 1933 -121
rect 1967 -1097 1979 -121
rect 1921 -1109 1979 -1097
rect 2179 -121 2237 -109
rect 2179 -1097 2191 -121
rect 2225 -1097 2237 -121
rect 2179 -1109 2237 -1097
rect 2299 -121 2357 -109
rect 2299 -1097 2311 -121
rect 2345 -1097 2357 -121
rect 2299 -1109 2357 -1097
rect 2557 -121 2615 -109
rect 2557 -1097 2569 -121
rect 2603 -1097 2615 -121
rect 2557 -1109 2615 -1097
rect 2677 -121 2735 -109
rect 2677 -1097 2689 -121
rect 2723 -1097 2735 -121
rect 2677 -1109 2735 -1097
rect 2935 -121 2993 -109
rect 2935 -1097 2947 -121
rect 2981 -1097 2993 -121
rect 2935 -1109 2993 -1097
rect 3055 -121 3113 -109
rect 3055 -1097 3067 -121
rect 3101 -1097 3113 -121
rect 3055 -1109 3113 -1097
rect 3313 -121 3371 -109
rect 3313 -1097 3325 -121
rect 3359 -1097 3371 -121
rect 3313 -1109 3371 -1097
rect 3433 -121 3491 -109
rect 3433 -1097 3445 -121
rect 3479 -1097 3491 -121
rect 3433 -1109 3491 -1097
rect 3691 -121 3749 -109
rect 3691 -1097 3703 -121
rect 3737 -1097 3749 -121
rect 3691 -1109 3749 -1097
rect 3811 -121 3869 -109
rect 3811 -1097 3823 -121
rect 3857 -1097 3869 -121
rect 3811 -1109 3869 -1097
rect 4069 -121 4127 -109
rect 4069 -1097 4081 -121
rect 4115 -1097 4127 -121
rect 4069 -1109 4127 -1097
rect 4189 -121 4247 -109
rect 4189 -1097 4201 -121
rect 4235 -1097 4247 -121
rect 4189 -1109 4247 -1097
rect 4447 -121 4505 -109
rect 4447 -1097 4459 -121
rect 4493 -1097 4505 -121
rect 4447 -1109 4505 -1097
rect 4567 -121 4625 -109
rect 4567 -1097 4579 -121
rect 4613 -1097 4625 -121
rect 4567 -1109 4625 -1097
rect 4825 -121 4883 -109
rect 4825 -1097 4837 -121
rect 4871 -1097 4883 -121
rect 4825 -1109 4883 -1097
rect 4945 -121 5003 -109
rect 4945 -1097 4957 -121
rect 4991 -1097 5003 -121
rect 4945 -1109 5003 -1097
rect 5203 -121 5261 -109
rect 5203 -1097 5215 -121
rect 5249 -1097 5261 -121
rect 5203 -1109 5261 -1097
rect 5323 -121 5381 -109
rect 5323 -1097 5335 -121
rect 5369 -1097 5381 -121
rect 5323 -1109 5381 -1097
rect 5581 -121 5639 -109
rect 5581 -1097 5593 -121
rect 5627 -1097 5639 -121
rect 5581 -1109 5639 -1097
rect 5701 -121 5759 -109
rect 5701 -1097 5713 -121
rect 5747 -1097 5759 -121
rect 5701 -1109 5759 -1097
rect 5959 -121 6017 -109
rect 5959 -1097 5971 -121
rect 6005 -1097 6017 -121
rect 5959 -1109 6017 -1097
rect 6079 -121 6137 -109
rect 6079 -1097 6091 -121
rect 6125 -1097 6137 -121
rect 6079 -1109 6137 -1097
rect 6337 -121 6395 -109
rect 6337 -1097 6349 -121
rect 6383 -1097 6395 -121
rect 6337 -1109 6395 -1097
rect 6457 -121 6515 -109
rect 6457 -1097 6469 -121
rect 6503 -1097 6515 -121
rect 6457 -1109 6515 -1097
rect 6715 -121 6773 -109
rect 6715 -1097 6727 -121
rect 6761 -1097 6773 -121
rect 6715 -1109 6773 -1097
rect 6835 -121 6893 -109
rect 6835 -1097 6847 -121
rect 6881 -1097 6893 -121
rect 6835 -1109 6893 -1097
rect 7093 -121 7151 -109
rect 7093 -1097 7105 -121
rect 7139 -1097 7151 -121
rect 7093 -1109 7151 -1097
rect 7213 -121 7271 -109
rect 7213 -1097 7225 -121
rect 7259 -1097 7271 -121
rect 7213 -1109 7271 -1097
rect 7471 -121 7529 -109
rect 7471 -1097 7483 -121
rect 7517 -1097 7529 -121
rect 7471 -1109 7529 -1097
rect 7591 -121 7649 -109
rect 7591 -1097 7603 -121
rect 7637 -1097 7649 -121
rect 7591 -1109 7649 -1097
rect 7849 -121 7907 -109
rect 7849 -1097 7861 -121
rect 7895 -1097 7907 -121
rect 7849 -1109 7907 -1097
rect 7969 -121 8027 -109
rect 7969 -1097 7981 -121
rect 8015 -1097 8027 -121
rect 7969 -1109 8027 -1097
rect 8227 -121 8285 -109
rect 8227 -1097 8239 -121
rect 8273 -1097 8285 -121
rect 8227 -1109 8285 -1097
rect 8347 -121 8405 -109
rect 8347 -1097 8359 -121
rect 8393 -1097 8405 -121
rect 8347 -1109 8405 -1097
rect 8605 -121 8663 -109
rect 8605 -1097 8617 -121
rect 8651 -1097 8663 -121
rect 8605 -1109 8663 -1097
rect 8725 -121 8783 -109
rect 8725 -1097 8737 -121
rect 8771 -1097 8783 -121
rect 8725 -1109 8783 -1097
rect 8983 -121 9041 -109
rect 8983 -1097 8995 -121
rect 9029 -1097 9041 -121
rect 8983 -1109 9041 -1097
rect 9103 -121 9161 -109
rect 9103 -1097 9115 -121
rect 9149 -1097 9161 -121
rect 9103 -1109 9161 -1097
rect 9361 -121 9419 -109
rect 9361 -1097 9373 -121
rect 9407 -1097 9419 -121
rect 9361 -1109 9419 -1097
rect -9419 -1339 -9361 -1327
rect -9419 -2315 -9407 -1339
rect -9373 -2315 -9361 -1339
rect -9419 -2327 -9361 -2315
rect -9161 -1339 -9103 -1327
rect -9161 -2315 -9149 -1339
rect -9115 -2315 -9103 -1339
rect -9161 -2327 -9103 -2315
rect -9041 -1339 -8983 -1327
rect -9041 -2315 -9029 -1339
rect -8995 -2315 -8983 -1339
rect -9041 -2327 -8983 -2315
rect -8783 -1339 -8725 -1327
rect -8783 -2315 -8771 -1339
rect -8737 -2315 -8725 -1339
rect -8783 -2327 -8725 -2315
rect -8663 -1339 -8605 -1327
rect -8663 -2315 -8651 -1339
rect -8617 -2315 -8605 -1339
rect -8663 -2327 -8605 -2315
rect -8405 -1339 -8347 -1327
rect -8405 -2315 -8393 -1339
rect -8359 -2315 -8347 -1339
rect -8405 -2327 -8347 -2315
rect -8285 -1339 -8227 -1327
rect -8285 -2315 -8273 -1339
rect -8239 -2315 -8227 -1339
rect -8285 -2327 -8227 -2315
rect -8027 -1339 -7969 -1327
rect -8027 -2315 -8015 -1339
rect -7981 -2315 -7969 -1339
rect -8027 -2327 -7969 -2315
rect -7907 -1339 -7849 -1327
rect -7907 -2315 -7895 -1339
rect -7861 -2315 -7849 -1339
rect -7907 -2327 -7849 -2315
rect -7649 -1339 -7591 -1327
rect -7649 -2315 -7637 -1339
rect -7603 -2315 -7591 -1339
rect -7649 -2327 -7591 -2315
rect -7529 -1339 -7471 -1327
rect -7529 -2315 -7517 -1339
rect -7483 -2315 -7471 -1339
rect -7529 -2327 -7471 -2315
rect -7271 -1339 -7213 -1327
rect -7271 -2315 -7259 -1339
rect -7225 -2315 -7213 -1339
rect -7271 -2327 -7213 -2315
rect -7151 -1339 -7093 -1327
rect -7151 -2315 -7139 -1339
rect -7105 -2315 -7093 -1339
rect -7151 -2327 -7093 -2315
rect -6893 -1339 -6835 -1327
rect -6893 -2315 -6881 -1339
rect -6847 -2315 -6835 -1339
rect -6893 -2327 -6835 -2315
rect -6773 -1339 -6715 -1327
rect -6773 -2315 -6761 -1339
rect -6727 -2315 -6715 -1339
rect -6773 -2327 -6715 -2315
rect -6515 -1339 -6457 -1327
rect -6515 -2315 -6503 -1339
rect -6469 -2315 -6457 -1339
rect -6515 -2327 -6457 -2315
rect -6395 -1339 -6337 -1327
rect -6395 -2315 -6383 -1339
rect -6349 -2315 -6337 -1339
rect -6395 -2327 -6337 -2315
rect -6137 -1339 -6079 -1327
rect -6137 -2315 -6125 -1339
rect -6091 -2315 -6079 -1339
rect -6137 -2327 -6079 -2315
rect -6017 -1339 -5959 -1327
rect -6017 -2315 -6005 -1339
rect -5971 -2315 -5959 -1339
rect -6017 -2327 -5959 -2315
rect -5759 -1339 -5701 -1327
rect -5759 -2315 -5747 -1339
rect -5713 -2315 -5701 -1339
rect -5759 -2327 -5701 -2315
rect -5639 -1339 -5581 -1327
rect -5639 -2315 -5627 -1339
rect -5593 -2315 -5581 -1339
rect -5639 -2327 -5581 -2315
rect -5381 -1339 -5323 -1327
rect -5381 -2315 -5369 -1339
rect -5335 -2315 -5323 -1339
rect -5381 -2327 -5323 -2315
rect -5261 -1339 -5203 -1327
rect -5261 -2315 -5249 -1339
rect -5215 -2315 -5203 -1339
rect -5261 -2327 -5203 -2315
rect -5003 -1339 -4945 -1327
rect -5003 -2315 -4991 -1339
rect -4957 -2315 -4945 -1339
rect -5003 -2327 -4945 -2315
rect -4883 -1339 -4825 -1327
rect -4883 -2315 -4871 -1339
rect -4837 -2315 -4825 -1339
rect -4883 -2327 -4825 -2315
rect -4625 -1339 -4567 -1327
rect -4625 -2315 -4613 -1339
rect -4579 -2315 -4567 -1339
rect -4625 -2327 -4567 -2315
rect -4505 -1339 -4447 -1327
rect -4505 -2315 -4493 -1339
rect -4459 -2315 -4447 -1339
rect -4505 -2327 -4447 -2315
rect -4247 -1339 -4189 -1327
rect -4247 -2315 -4235 -1339
rect -4201 -2315 -4189 -1339
rect -4247 -2327 -4189 -2315
rect -4127 -1339 -4069 -1327
rect -4127 -2315 -4115 -1339
rect -4081 -2315 -4069 -1339
rect -4127 -2327 -4069 -2315
rect -3869 -1339 -3811 -1327
rect -3869 -2315 -3857 -1339
rect -3823 -2315 -3811 -1339
rect -3869 -2327 -3811 -2315
rect -3749 -1339 -3691 -1327
rect -3749 -2315 -3737 -1339
rect -3703 -2315 -3691 -1339
rect -3749 -2327 -3691 -2315
rect -3491 -1339 -3433 -1327
rect -3491 -2315 -3479 -1339
rect -3445 -2315 -3433 -1339
rect -3491 -2327 -3433 -2315
rect -3371 -1339 -3313 -1327
rect -3371 -2315 -3359 -1339
rect -3325 -2315 -3313 -1339
rect -3371 -2327 -3313 -2315
rect -3113 -1339 -3055 -1327
rect -3113 -2315 -3101 -1339
rect -3067 -2315 -3055 -1339
rect -3113 -2327 -3055 -2315
rect -2993 -1339 -2935 -1327
rect -2993 -2315 -2981 -1339
rect -2947 -2315 -2935 -1339
rect -2993 -2327 -2935 -2315
rect -2735 -1339 -2677 -1327
rect -2735 -2315 -2723 -1339
rect -2689 -2315 -2677 -1339
rect -2735 -2327 -2677 -2315
rect -2615 -1339 -2557 -1327
rect -2615 -2315 -2603 -1339
rect -2569 -2315 -2557 -1339
rect -2615 -2327 -2557 -2315
rect -2357 -1339 -2299 -1327
rect -2357 -2315 -2345 -1339
rect -2311 -2315 -2299 -1339
rect -2357 -2327 -2299 -2315
rect -2237 -1339 -2179 -1327
rect -2237 -2315 -2225 -1339
rect -2191 -2315 -2179 -1339
rect -2237 -2327 -2179 -2315
rect -1979 -1339 -1921 -1327
rect -1979 -2315 -1967 -1339
rect -1933 -2315 -1921 -1339
rect -1979 -2327 -1921 -2315
rect -1859 -1339 -1801 -1327
rect -1859 -2315 -1847 -1339
rect -1813 -2315 -1801 -1339
rect -1859 -2327 -1801 -2315
rect -1601 -1339 -1543 -1327
rect -1601 -2315 -1589 -1339
rect -1555 -2315 -1543 -1339
rect -1601 -2327 -1543 -2315
rect -1481 -1339 -1423 -1327
rect -1481 -2315 -1469 -1339
rect -1435 -2315 -1423 -1339
rect -1481 -2327 -1423 -2315
rect -1223 -1339 -1165 -1327
rect -1223 -2315 -1211 -1339
rect -1177 -2315 -1165 -1339
rect -1223 -2327 -1165 -2315
rect -1103 -1339 -1045 -1327
rect -1103 -2315 -1091 -1339
rect -1057 -2315 -1045 -1339
rect -1103 -2327 -1045 -2315
rect -845 -1339 -787 -1327
rect -845 -2315 -833 -1339
rect -799 -2315 -787 -1339
rect -845 -2327 -787 -2315
rect -725 -1339 -667 -1327
rect -725 -2315 -713 -1339
rect -679 -2315 -667 -1339
rect -725 -2327 -667 -2315
rect -467 -1339 -409 -1327
rect -467 -2315 -455 -1339
rect -421 -2315 -409 -1339
rect -467 -2327 -409 -2315
rect -347 -1339 -289 -1327
rect -347 -2315 -335 -1339
rect -301 -2315 -289 -1339
rect -347 -2327 -289 -2315
rect -89 -1339 -31 -1327
rect -89 -2315 -77 -1339
rect -43 -2315 -31 -1339
rect -89 -2327 -31 -2315
rect 31 -1339 89 -1327
rect 31 -2315 43 -1339
rect 77 -2315 89 -1339
rect 31 -2327 89 -2315
rect 289 -1339 347 -1327
rect 289 -2315 301 -1339
rect 335 -2315 347 -1339
rect 289 -2327 347 -2315
rect 409 -1339 467 -1327
rect 409 -2315 421 -1339
rect 455 -2315 467 -1339
rect 409 -2327 467 -2315
rect 667 -1339 725 -1327
rect 667 -2315 679 -1339
rect 713 -2315 725 -1339
rect 667 -2327 725 -2315
rect 787 -1339 845 -1327
rect 787 -2315 799 -1339
rect 833 -2315 845 -1339
rect 787 -2327 845 -2315
rect 1045 -1339 1103 -1327
rect 1045 -2315 1057 -1339
rect 1091 -2315 1103 -1339
rect 1045 -2327 1103 -2315
rect 1165 -1339 1223 -1327
rect 1165 -2315 1177 -1339
rect 1211 -2315 1223 -1339
rect 1165 -2327 1223 -2315
rect 1423 -1339 1481 -1327
rect 1423 -2315 1435 -1339
rect 1469 -2315 1481 -1339
rect 1423 -2327 1481 -2315
rect 1543 -1339 1601 -1327
rect 1543 -2315 1555 -1339
rect 1589 -2315 1601 -1339
rect 1543 -2327 1601 -2315
rect 1801 -1339 1859 -1327
rect 1801 -2315 1813 -1339
rect 1847 -2315 1859 -1339
rect 1801 -2327 1859 -2315
rect 1921 -1339 1979 -1327
rect 1921 -2315 1933 -1339
rect 1967 -2315 1979 -1339
rect 1921 -2327 1979 -2315
rect 2179 -1339 2237 -1327
rect 2179 -2315 2191 -1339
rect 2225 -2315 2237 -1339
rect 2179 -2327 2237 -2315
rect 2299 -1339 2357 -1327
rect 2299 -2315 2311 -1339
rect 2345 -2315 2357 -1339
rect 2299 -2327 2357 -2315
rect 2557 -1339 2615 -1327
rect 2557 -2315 2569 -1339
rect 2603 -2315 2615 -1339
rect 2557 -2327 2615 -2315
rect 2677 -1339 2735 -1327
rect 2677 -2315 2689 -1339
rect 2723 -2315 2735 -1339
rect 2677 -2327 2735 -2315
rect 2935 -1339 2993 -1327
rect 2935 -2315 2947 -1339
rect 2981 -2315 2993 -1339
rect 2935 -2327 2993 -2315
rect 3055 -1339 3113 -1327
rect 3055 -2315 3067 -1339
rect 3101 -2315 3113 -1339
rect 3055 -2327 3113 -2315
rect 3313 -1339 3371 -1327
rect 3313 -2315 3325 -1339
rect 3359 -2315 3371 -1339
rect 3313 -2327 3371 -2315
rect 3433 -1339 3491 -1327
rect 3433 -2315 3445 -1339
rect 3479 -2315 3491 -1339
rect 3433 -2327 3491 -2315
rect 3691 -1339 3749 -1327
rect 3691 -2315 3703 -1339
rect 3737 -2315 3749 -1339
rect 3691 -2327 3749 -2315
rect 3811 -1339 3869 -1327
rect 3811 -2315 3823 -1339
rect 3857 -2315 3869 -1339
rect 3811 -2327 3869 -2315
rect 4069 -1339 4127 -1327
rect 4069 -2315 4081 -1339
rect 4115 -2315 4127 -1339
rect 4069 -2327 4127 -2315
rect 4189 -1339 4247 -1327
rect 4189 -2315 4201 -1339
rect 4235 -2315 4247 -1339
rect 4189 -2327 4247 -2315
rect 4447 -1339 4505 -1327
rect 4447 -2315 4459 -1339
rect 4493 -2315 4505 -1339
rect 4447 -2327 4505 -2315
rect 4567 -1339 4625 -1327
rect 4567 -2315 4579 -1339
rect 4613 -2315 4625 -1339
rect 4567 -2327 4625 -2315
rect 4825 -1339 4883 -1327
rect 4825 -2315 4837 -1339
rect 4871 -2315 4883 -1339
rect 4825 -2327 4883 -2315
rect 4945 -1339 5003 -1327
rect 4945 -2315 4957 -1339
rect 4991 -2315 5003 -1339
rect 4945 -2327 5003 -2315
rect 5203 -1339 5261 -1327
rect 5203 -2315 5215 -1339
rect 5249 -2315 5261 -1339
rect 5203 -2327 5261 -2315
rect 5323 -1339 5381 -1327
rect 5323 -2315 5335 -1339
rect 5369 -2315 5381 -1339
rect 5323 -2327 5381 -2315
rect 5581 -1339 5639 -1327
rect 5581 -2315 5593 -1339
rect 5627 -2315 5639 -1339
rect 5581 -2327 5639 -2315
rect 5701 -1339 5759 -1327
rect 5701 -2315 5713 -1339
rect 5747 -2315 5759 -1339
rect 5701 -2327 5759 -2315
rect 5959 -1339 6017 -1327
rect 5959 -2315 5971 -1339
rect 6005 -2315 6017 -1339
rect 5959 -2327 6017 -2315
rect 6079 -1339 6137 -1327
rect 6079 -2315 6091 -1339
rect 6125 -2315 6137 -1339
rect 6079 -2327 6137 -2315
rect 6337 -1339 6395 -1327
rect 6337 -2315 6349 -1339
rect 6383 -2315 6395 -1339
rect 6337 -2327 6395 -2315
rect 6457 -1339 6515 -1327
rect 6457 -2315 6469 -1339
rect 6503 -2315 6515 -1339
rect 6457 -2327 6515 -2315
rect 6715 -1339 6773 -1327
rect 6715 -2315 6727 -1339
rect 6761 -2315 6773 -1339
rect 6715 -2327 6773 -2315
rect 6835 -1339 6893 -1327
rect 6835 -2315 6847 -1339
rect 6881 -2315 6893 -1339
rect 6835 -2327 6893 -2315
rect 7093 -1339 7151 -1327
rect 7093 -2315 7105 -1339
rect 7139 -2315 7151 -1339
rect 7093 -2327 7151 -2315
rect 7213 -1339 7271 -1327
rect 7213 -2315 7225 -1339
rect 7259 -2315 7271 -1339
rect 7213 -2327 7271 -2315
rect 7471 -1339 7529 -1327
rect 7471 -2315 7483 -1339
rect 7517 -2315 7529 -1339
rect 7471 -2327 7529 -2315
rect 7591 -1339 7649 -1327
rect 7591 -2315 7603 -1339
rect 7637 -2315 7649 -1339
rect 7591 -2327 7649 -2315
rect 7849 -1339 7907 -1327
rect 7849 -2315 7861 -1339
rect 7895 -2315 7907 -1339
rect 7849 -2327 7907 -2315
rect 7969 -1339 8027 -1327
rect 7969 -2315 7981 -1339
rect 8015 -2315 8027 -1339
rect 7969 -2327 8027 -2315
rect 8227 -1339 8285 -1327
rect 8227 -2315 8239 -1339
rect 8273 -2315 8285 -1339
rect 8227 -2327 8285 -2315
rect 8347 -1339 8405 -1327
rect 8347 -2315 8359 -1339
rect 8393 -2315 8405 -1339
rect 8347 -2327 8405 -2315
rect 8605 -1339 8663 -1327
rect 8605 -2315 8617 -1339
rect 8651 -2315 8663 -1339
rect 8605 -2327 8663 -2315
rect 8725 -1339 8783 -1327
rect 8725 -2315 8737 -1339
rect 8771 -2315 8783 -1339
rect 8725 -2327 8783 -2315
rect 8983 -1339 9041 -1327
rect 8983 -2315 8995 -1339
rect 9029 -2315 9041 -1339
rect 8983 -2327 9041 -2315
rect 9103 -1339 9161 -1327
rect 9103 -2315 9115 -1339
rect 9149 -2315 9161 -1339
rect 9103 -2327 9161 -2315
rect 9361 -1339 9419 -1327
rect 9361 -2315 9373 -1339
rect 9407 -2315 9419 -1339
rect 9361 -2327 9419 -2315
<< mvndiffc >>
rect -9407 1339 -9373 2315
rect -9149 1339 -9115 2315
rect -9029 1339 -8995 2315
rect -8771 1339 -8737 2315
rect -8651 1339 -8617 2315
rect -8393 1339 -8359 2315
rect -8273 1339 -8239 2315
rect -8015 1339 -7981 2315
rect -7895 1339 -7861 2315
rect -7637 1339 -7603 2315
rect -7517 1339 -7483 2315
rect -7259 1339 -7225 2315
rect -7139 1339 -7105 2315
rect -6881 1339 -6847 2315
rect -6761 1339 -6727 2315
rect -6503 1339 -6469 2315
rect -6383 1339 -6349 2315
rect -6125 1339 -6091 2315
rect -6005 1339 -5971 2315
rect -5747 1339 -5713 2315
rect -5627 1339 -5593 2315
rect -5369 1339 -5335 2315
rect -5249 1339 -5215 2315
rect -4991 1339 -4957 2315
rect -4871 1339 -4837 2315
rect -4613 1339 -4579 2315
rect -4493 1339 -4459 2315
rect -4235 1339 -4201 2315
rect -4115 1339 -4081 2315
rect -3857 1339 -3823 2315
rect -3737 1339 -3703 2315
rect -3479 1339 -3445 2315
rect -3359 1339 -3325 2315
rect -3101 1339 -3067 2315
rect -2981 1339 -2947 2315
rect -2723 1339 -2689 2315
rect -2603 1339 -2569 2315
rect -2345 1339 -2311 2315
rect -2225 1339 -2191 2315
rect -1967 1339 -1933 2315
rect -1847 1339 -1813 2315
rect -1589 1339 -1555 2315
rect -1469 1339 -1435 2315
rect -1211 1339 -1177 2315
rect -1091 1339 -1057 2315
rect -833 1339 -799 2315
rect -713 1339 -679 2315
rect -455 1339 -421 2315
rect -335 1339 -301 2315
rect -77 1339 -43 2315
rect 43 1339 77 2315
rect 301 1339 335 2315
rect 421 1339 455 2315
rect 679 1339 713 2315
rect 799 1339 833 2315
rect 1057 1339 1091 2315
rect 1177 1339 1211 2315
rect 1435 1339 1469 2315
rect 1555 1339 1589 2315
rect 1813 1339 1847 2315
rect 1933 1339 1967 2315
rect 2191 1339 2225 2315
rect 2311 1339 2345 2315
rect 2569 1339 2603 2315
rect 2689 1339 2723 2315
rect 2947 1339 2981 2315
rect 3067 1339 3101 2315
rect 3325 1339 3359 2315
rect 3445 1339 3479 2315
rect 3703 1339 3737 2315
rect 3823 1339 3857 2315
rect 4081 1339 4115 2315
rect 4201 1339 4235 2315
rect 4459 1339 4493 2315
rect 4579 1339 4613 2315
rect 4837 1339 4871 2315
rect 4957 1339 4991 2315
rect 5215 1339 5249 2315
rect 5335 1339 5369 2315
rect 5593 1339 5627 2315
rect 5713 1339 5747 2315
rect 5971 1339 6005 2315
rect 6091 1339 6125 2315
rect 6349 1339 6383 2315
rect 6469 1339 6503 2315
rect 6727 1339 6761 2315
rect 6847 1339 6881 2315
rect 7105 1339 7139 2315
rect 7225 1339 7259 2315
rect 7483 1339 7517 2315
rect 7603 1339 7637 2315
rect 7861 1339 7895 2315
rect 7981 1339 8015 2315
rect 8239 1339 8273 2315
rect 8359 1339 8393 2315
rect 8617 1339 8651 2315
rect 8737 1339 8771 2315
rect 8995 1339 9029 2315
rect 9115 1339 9149 2315
rect 9373 1339 9407 2315
rect -9407 121 -9373 1097
rect -9149 121 -9115 1097
rect -9029 121 -8995 1097
rect -8771 121 -8737 1097
rect -8651 121 -8617 1097
rect -8393 121 -8359 1097
rect -8273 121 -8239 1097
rect -8015 121 -7981 1097
rect -7895 121 -7861 1097
rect -7637 121 -7603 1097
rect -7517 121 -7483 1097
rect -7259 121 -7225 1097
rect -7139 121 -7105 1097
rect -6881 121 -6847 1097
rect -6761 121 -6727 1097
rect -6503 121 -6469 1097
rect -6383 121 -6349 1097
rect -6125 121 -6091 1097
rect -6005 121 -5971 1097
rect -5747 121 -5713 1097
rect -5627 121 -5593 1097
rect -5369 121 -5335 1097
rect -5249 121 -5215 1097
rect -4991 121 -4957 1097
rect -4871 121 -4837 1097
rect -4613 121 -4579 1097
rect -4493 121 -4459 1097
rect -4235 121 -4201 1097
rect -4115 121 -4081 1097
rect -3857 121 -3823 1097
rect -3737 121 -3703 1097
rect -3479 121 -3445 1097
rect -3359 121 -3325 1097
rect -3101 121 -3067 1097
rect -2981 121 -2947 1097
rect -2723 121 -2689 1097
rect -2603 121 -2569 1097
rect -2345 121 -2311 1097
rect -2225 121 -2191 1097
rect -1967 121 -1933 1097
rect -1847 121 -1813 1097
rect -1589 121 -1555 1097
rect -1469 121 -1435 1097
rect -1211 121 -1177 1097
rect -1091 121 -1057 1097
rect -833 121 -799 1097
rect -713 121 -679 1097
rect -455 121 -421 1097
rect -335 121 -301 1097
rect -77 121 -43 1097
rect 43 121 77 1097
rect 301 121 335 1097
rect 421 121 455 1097
rect 679 121 713 1097
rect 799 121 833 1097
rect 1057 121 1091 1097
rect 1177 121 1211 1097
rect 1435 121 1469 1097
rect 1555 121 1589 1097
rect 1813 121 1847 1097
rect 1933 121 1967 1097
rect 2191 121 2225 1097
rect 2311 121 2345 1097
rect 2569 121 2603 1097
rect 2689 121 2723 1097
rect 2947 121 2981 1097
rect 3067 121 3101 1097
rect 3325 121 3359 1097
rect 3445 121 3479 1097
rect 3703 121 3737 1097
rect 3823 121 3857 1097
rect 4081 121 4115 1097
rect 4201 121 4235 1097
rect 4459 121 4493 1097
rect 4579 121 4613 1097
rect 4837 121 4871 1097
rect 4957 121 4991 1097
rect 5215 121 5249 1097
rect 5335 121 5369 1097
rect 5593 121 5627 1097
rect 5713 121 5747 1097
rect 5971 121 6005 1097
rect 6091 121 6125 1097
rect 6349 121 6383 1097
rect 6469 121 6503 1097
rect 6727 121 6761 1097
rect 6847 121 6881 1097
rect 7105 121 7139 1097
rect 7225 121 7259 1097
rect 7483 121 7517 1097
rect 7603 121 7637 1097
rect 7861 121 7895 1097
rect 7981 121 8015 1097
rect 8239 121 8273 1097
rect 8359 121 8393 1097
rect 8617 121 8651 1097
rect 8737 121 8771 1097
rect 8995 121 9029 1097
rect 9115 121 9149 1097
rect 9373 121 9407 1097
rect -9407 -1097 -9373 -121
rect -9149 -1097 -9115 -121
rect -9029 -1097 -8995 -121
rect -8771 -1097 -8737 -121
rect -8651 -1097 -8617 -121
rect -8393 -1097 -8359 -121
rect -8273 -1097 -8239 -121
rect -8015 -1097 -7981 -121
rect -7895 -1097 -7861 -121
rect -7637 -1097 -7603 -121
rect -7517 -1097 -7483 -121
rect -7259 -1097 -7225 -121
rect -7139 -1097 -7105 -121
rect -6881 -1097 -6847 -121
rect -6761 -1097 -6727 -121
rect -6503 -1097 -6469 -121
rect -6383 -1097 -6349 -121
rect -6125 -1097 -6091 -121
rect -6005 -1097 -5971 -121
rect -5747 -1097 -5713 -121
rect -5627 -1097 -5593 -121
rect -5369 -1097 -5335 -121
rect -5249 -1097 -5215 -121
rect -4991 -1097 -4957 -121
rect -4871 -1097 -4837 -121
rect -4613 -1097 -4579 -121
rect -4493 -1097 -4459 -121
rect -4235 -1097 -4201 -121
rect -4115 -1097 -4081 -121
rect -3857 -1097 -3823 -121
rect -3737 -1097 -3703 -121
rect -3479 -1097 -3445 -121
rect -3359 -1097 -3325 -121
rect -3101 -1097 -3067 -121
rect -2981 -1097 -2947 -121
rect -2723 -1097 -2689 -121
rect -2603 -1097 -2569 -121
rect -2345 -1097 -2311 -121
rect -2225 -1097 -2191 -121
rect -1967 -1097 -1933 -121
rect -1847 -1097 -1813 -121
rect -1589 -1097 -1555 -121
rect -1469 -1097 -1435 -121
rect -1211 -1097 -1177 -121
rect -1091 -1097 -1057 -121
rect -833 -1097 -799 -121
rect -713 -1097 -679 -121
rect -455 -1097 -421 -121
rect -335 -1097 -301 -121
rect -77 -1097 -43 -121
rect 43 -1097 77 -121
rect 301 -1097 335 -121
rect 421 -1097 455 -121
rect 679 -1097 713 -121
rect 799 -1097 833 -121
rect 1057 -1097 1091 -121
rect 1177 -1097 1211 -121
rect 1435 -1097 1469 -121
rect 1555 -1097 1589 -121
rect 1813 -1097 1847 -121
rect 1933 -1097 1967 -121
rect 2191 -1097 2225 -121
rect 2311 -1097 2345 -121
rect 2569 -1097 2603 -121
rect 2689 -1097 2723 -121
rect 2947 -1097 2981 -121
rect 3067 -1097 3101 -121
rect 3325 -1097 3359 -121
rect 3445 -1097 3479 -121
rect 3703 -1097 3737 -121
rect 3823 -1097 3857 -121
rect 4081 -1097 4115 -121
rect 4201 -1097 4235 -121
rect 4459 -1097 4493 -121
rect 4579 -1097 4613 -121
rect 4837 -1097 4871 -121
rect 4957 -1097 4991 -121
rect 5215 -1097 5249 -121
rect 5335 -1097 5369 -121
rect 5593 -1097 5627 -121
rect 5713 -1097 5747 -121
rect 5971 -1097 6005 -121
rect 6091 -1097 6125 -121
rect 6349 -1097 6383 -121
rect 6469 -1097 6503 -121
rect 6727 -1097 6761 -121
rect 6847 -1097 6881 -121
rect 7105 -1097 7139 -121
rect 7225 -1097 7259 -121
rect 7483 -1097 7517 -121
rect 7603 -1097 7637 -121
rect 7861 -1097 7895 -121
rect 7981 -1097 8015 -121
rect 8239 -1097 8273 -121
rect 8359 -1097 8393 -121
rect 8617 -1097 8651 -121
rect 8737 -1097 8771 -121
rect 8995 -1097 9029 -121
rect 9115 -1097 9149 -121
rect 9373 -1097 9407 -121
rect -9407 -2315 -9373 -1339
rect -9149 -2315 -9115 -1339
rect -9029 -2315 -8995 -1339
rect -8771 -2315 -8737 -1339
rect -8651 -2315 -8617 -1339
rect -8393 -2315 -8359 -1339
rect -8273 -2315 -8239 -1339
rect -8015 -2315 -7981 -1339
rect -7895 -2315 -7861 -1339
rect -7637 -2315 -7603 -1339
rect -7517 -2315 -7483 -1339
rect -7259 -2315 -7225 -1339
rect -7139 -2315 -7105 -1339
rect -6881 -2315 -6847 -1339
rect -6761 -2315 -6727 -1339
rect -6503 -2315 -6469 -1339
rect -6383 -2315 -6349 -1339
rect -6125 -2315 -6091 -1339
rect -6005 -2315 -5971 -1339
rect -5747 -2315 -5713 -1339
rect -5627 -2315 -5593 -1339
rect -5369 -2315 -5335 -1339
rect -5249 -2315 -5215 -1339
rect -4991 -2315 -4957 -1339
rect -4871 -2315 -4837 -1339
rect -4613 -2315 -4579 -1339
rect -4493 -2315 -4459 -1339
rect -4235 -2315 -4201 -1339
rect -4115 -2315 -4081 -1339
rect -3857 -2315 -3823 -1339
rect -3737 -2315 -3703 -1339
rect -3479 -2315 -3445 -1339
rect -3359 -2315 -3325 -1339
rect -3101 -2315 -3067 -1339
rect -2981 -2315 -2947 -1339
rect -2723 -2315 -2689 -1339
rect -2603 -2315 -2569 -1339
rect -2345 -2315 -2311 -1339
rect -2225 -2315 -2191 -1339
rect -1967 -2315 -1933 -1339
rect -1847 -2315 -1813 -1339
rect -1589 -2315 -1555 -1339
rect -1469 -2315 -1435 -1339
rect -1211 -2315 -1177 -1339
rect -1091 -2315 -1057 -1339
rect -833 -2315 -799 -1339
rect -713 -2315 -679 -1339
rect -455 -2315 -421 -1339
rect -335 -2315 -301 -1339
rect -77 -2315 -43 -1339
rect 43 -2315 77 -1339
rect 301 -2315 335 -1339
rect 421 -2315 455 -1339
rect 679 -2315 713 -1339
rect 799 -2315 833 -1339
rect 1057 -2315 1091 -1339
rect 1177 -2315 1211 -1339
rect 1435 -2315 1469 -1339
rect 1555 -2315 1589 -1339
rect 1813 -2315 1847 -1339
rect 1933 -2315 1967 -1339
rect 2191 -2315 2225 -1339
rect 2311 -2315 2345 -1339
rect 2569 -2315 2603 -1339
rect 2689 -2315 2723 -1339
rect 2947 -2315 2981 -1339
rect 3067 -2315 3101 -1339
rect 3325 -2315 3359 -1339
rect 3445 -2315 3479 -1339
rect 3703 -2315 3737 -1339
rect 3823 -2315 3857 -1339
rect 4081 -2315 4115 -1339
rect 4201 -2315 4235 -1339
rect 4459 -2315 4493 -1339
rect 4579 -2315 4613 -1339
rect 4837 -2315 4871 -1339
rect 4957 -2315 4991 -1339
rect 5215 -2315 5249 -1339
rect 5335 -2315 5369 -1339
rect 5593 -2315 5627 -1339
rect 5713 -2315 5747 -1339
rect 5971 -2315 6005 -1339
rect 6091 -2315 6125 -1339
rect 6349 -2315 6383 -1339
rect 6469 -2315 6503 -1339
rect 6727 -2315 6761 -1339
rect 6847 -2315 6881 -1339
rect 7105 -2315 7139 -1339
rect 7225 -2315 7259 -1339
rect 7483 -2315 7517 -1339
rect 7603 -2315 7637 -1339
rect 7861 -2315 7895 -1339
rect 7981 -2315 8015 -1339
rect 8239 -2315 8273 -1339
rect 8359 -2315 8393 -1339
rect 8617 -2315 8651 -1339
rect 8737 -2315 8771 -1339
rect 8995 -2315 9029 -1339
rect 9115 -2315 9149 -1339
rect 9373 -2315 9407 -1339
<< mvpsubdiff >>
rect -9553 2537 9553 2549
rect -9553 2503 -9445 2537
rect 9445 2503 9553 2537
rect -9553 2491 9553 2503
rect -9553 2441 -9495 2491
rect -9553 -2441 -9541 2441
rect -9507 -2441 -9495 2441
rect 9495 2441 9553 2491
rect -9553 -2491 -9495 -2441
rect 9495 -2441 9507 2441
rect 9541 -2441 9553 2441
rect 9495 -2491 9553 -2441
rect -9553 -2503 9553 -2491
rect -9553 -2537 -9445 -2503
rect 9445 -2537 9553 -2503
rect -9553 -2549 9553 -2537
<< mvpsubdiffcont >>
rect -9445 2503 9445 2537
rect -9541 -2441 -9507 2441
rect 9507 -2441 9541 2441
rect -9445 -2537 9445 -2503
<< poly >>
rect -9361 2399 -9161 2415
rect -9361 2365 -9345 2399
rect -9177 2365 -9161 2399
rect -9361 2327 -9161 2365
rect -8983 2399 -8783 2415
rect -8983 2365 -8967 2399
rect -8799 2365 -8783 2399
rect -8983 2327 -8783 2365
rect -8605 2399 -8405 2415
rect -8605 2365 -8589 2399
rect -8421 2365 -8405 2399
rect -8605 2327 -8405 2365
rect -8227 2399 -8027 2415
rect -8227 2365 -8211 2399
rect -8043 2365 -8027 2399
rect -8227 2327 -8027 2365
rect -7849 2399 -7649 2415
rect -7849 2365 -7833 2399
rect -7665 2365 -7649 2399
rect -7849 2327 -7649 2365
rect -7471 2399 -7271 2415
rect -7471 2365 -7455 2399
rect -7287 2365 -7271 2399
rect -7471 2327 -7271 2365
rect -7093 2399 -6893 2415
rect -7093 2365 -7077 2399
rect -6909 2365 -6893 2399
rect -7093 2327 -6893 2365
rect -6715 2399 -6515 2415
rect -6715 2365 -6699 2399
rect -6531 2365 -6515 2399
rect -6715 2327 -6515 2365
rect -6337 2399 -6137 2415
rect -6337 2365 -6321 2399
rect -6153 2365 -6137 2399
rect -6337 2327 -6137 2365
rect -5959 2399 -5759 2415
rect -5959 2365 -5943 2399
rect -5775 2365 -5759 2399
rect -5959 2327 -5759 2365
rect -5581 2399 -5381 2415
rect -5581 2365 -5565 2399
rect -5397 2365 -5381 2399
rect -5581 2327 -5381 2365
rect -5203 2399 -5003 2415
rect -5203 2365 -5187 2399
rect -5019 2365 -5003 2399
rect -5203 2327 -5003 2365
rect -4825 2399 -4625 2415
rect -4825 2365 -4809 2399
rect -4641 2365 -4625 2399
rect -4825 2327 -4625 2365
rect -4447 2399 -4247 2415
rect -4447 2365 -4431 2399
rect -4263 2365 -4247 2399
rect -4447 2327 -4247 2365
rect -4069 2399 -3869 2415
rect -4069 2365 -4053 2399
rect -3885 2365 -3869 2399
rect -4069 2327 -3869 2365
rect -3691 2399 -3491 2415
rect -3691 2365 -3675 2399
rect -3507 2365 -3491 2399
rect -3691 2327 -3491 2365
rect -3313 2399 -3113 2415
rect -3313 2365 -3297 2399
rect -3129 2365 -3113 2399
rect -3313 2327 -3113 2365
rect -2935 2399 -2735 2415
rect -2935 2365 -2919 2399
rect -2751 2365 -2735 2399
rect -2935 2327 -2735 2365
rect -2557 2399 -2357 2415
rect -2557 2365 -2541 2399
rect -2373 2365 -2357 2399
rect -2557 2327 -2357 2365
rect -2179 2399 -1979 2415
rect -2179 2365 -2163 2399
rect -1995 2365 -1979 2399
rect -2179 2327 -1979 2365
rect -1801 2399 -1601 2415
rect -1801 2365 -1785 2399
rect -1617 2365 -1601 2399
rect -1801 2327 -1601 2365
rect -1423 2399 -1223 2415
rect -1423 2365 -1407 2399
rect -1239 2365 -1223 2399
rect -1423 2327 -1223 2365
rect -1045 2399 -845 2415
rect -1045 2365 -1029 2399
rect -861 2365 -845 2399
rect -1045 2327 -845 2365
rect -667 2399 -467 2415
rect -667 2365 -651 2399
rect -483 2365 -467 2399
rect -667 2327 -467 2365
rect -289 2399 -89 2415
rect -289 2365 -273 2399
rect -105 2365 -89 2399
rect -289 2327 -89 2365
rect 89 2399 289 2415
rect 89 2365 105 2399
rect 273 2365 289 2399
rect 89 2327 289 2365
rect 467 2399 667 2415
rect 467 2365 483 2399
rect 651 2365 667 2399
rect 467 2327 667 2365
rect 845 2399 1045 2415
rect 845 2365 861 2399
rect 1029 2365 1045 2399
rect 845 2327 1045 2365
rect 1223 2399 1423 2415
rect 1223 2365 1239 2399
rect 1407 2365 1423 2399
rect 1223 2327 1423 2365
rect 1601 2399 1801 2415
rect 1601 2365 1617 2399
rect 1785 2365 1801 2399
rect 1601 2327 1801 2365
rect 1979 2399 2179 2415
rect 1979 2365 1995 2399
rect 2163 2365 2179 2399
rect 1979 2327 2179 2365
rect 2357 2399 2557 2415
rect 2357 2365 2373 2399
rect 2541 2365 2557 2399
rect 2357 2327 2557 2365
rect 2735 2399 2935 2415
rect 2735 2365 2751 2399
rect 2919 2365 2935 2399
rect 2735 2327 2935 2365
rect 3113 2399 3313 2415
rect 3113 2365 3129 2399
rect 3297 2365 3313 2399
rect 3113 2327 3313 2365
rect 3491 2399 3691 2415
rect 3491 2365 3507 2399
rect 3675 2365 3691 2399
rect 3491 2327 3691 2365
rect 3869 2399 4069 2415
rect 3869 2365 3885 2399
rect 4053 2365 4069 2399
rect 3869 2327 4069 2365
rect 4247 2399 4447 2415
rect 4247 2365 4263 2399
rect 4431 2365 4447 2399
rect 4247 2327 4447 2365
rect 4625 2399 4825 2415
rect 4625 2365 4641 2399
rect 4809 2365 4825 2399
rect 4625 2327 4825 2365
rect 5003 2399 5203 2415
rect 5003 2365 5019 2399
rect 5187 2365 5203 2399
rect 5003 2327 5203 2365
rect 5381 2399 5581 2415
rect 5381 2365 5397 2399
rect 5565 2365 5581 2399
rect 5381 2327 5581 2365
rect 5759 2399 5959 2415
rect 5759 2365 5775 2399
rect 5943 2365 5959 2399
rect 5759 2327 5959 2365
rect 6137 2399 6337 2415
rect 6137 2365 6153 2399
rect 6321 2365 6337 2399
rect 6137 2327 6337 2365
rect 6515 2399 6715 2415
rect 6515 2365 6531 2399
rect 6699 2365 6715 2399
rect 6515 2327 6715 2365
rect 6893 2399 7093 2415
rect 6893 2365 6909 2399
rect 7077 2365 7093 2399
rect 6893 2327 7093 2365
rect 7271 2399 7471 2415
rect 7271 2365 7287 2399
rect 7455 2365 7471 2399
rect 7271 2327 7471 2365
rect 7649 2399 7849 2415
rect 7649 2365 7665 2399
rect 7833 2365 7849 2399
rect 7649 2327 7849 2365
rect 8027 2399 8227 2415
rect 8027 2365 8043 2399
rect 8211 2365 8227 2399
rect 8027 2327 8227 2365
rect 8405 2399 8605 2415
rect 8405 2365 8421 2399
rect 8589 2365 8605 2399
rect 8405 2327 8605 2365
rect 8783 2399 8983 2415
rect 8783 2365 8799 2399
rect 8967 2365 8983 2399
rect 8783 2327 8983 2365
rect 9161 2399 9361 2415
rect 9161 2365 9177 2399
rect 9345 2365 9361 2399
rect 9161 2327 9361 2365
rect -9361 1289 -9161 1327
rect -9361 1255 -9345 1289
rect -9177 1255 -9161 1289
rect -9361 1239 -9161 1255
rect -8983 1289 -8783 1327
rect -8983 1255 -8967 1289
rect -8799 1255 -8783 1289
rect -8983 1239 -8783 1255
rect -8605 1289 -8405 1327
rect -8605 1255 -8589 1289
rect -8421 1255 -8405 1289
rect -8605 1239 -8405 1255
rect -8227 1289 -8027 1327
rect -8227 1255 -8211 1289
rect -8043 1255 -8027 1289
rect -8227 1239 -8027 1255
rect -7849 1289 -7649 1327
rect -7849 1255 -7833 1289
rect -7665 1255 -7649 1289
rect -7849 1239 -7649 1255
rect -7471 1289 -7271 1327
rect -7471 1255 -7455 1289
rect -7287 1255 -7271 1289
rect -7471 1239 -7271 1255
rect -7093 1289 -6893 1327
rect -7093 1255 -7077 1289
rect -6909 1255 -6893 1289
rect -7093 1239 -6893 1255
rect -6715 1289 -6515 1327
rect -6715 1255 -6699 1289
rect -6531 1255 -6515 1289
rect -6715 1239 -6515 1255
rect -6337 1289 -6137 1327
rect -6337 1255 -6321 1289
rect -6153 1255 -6137 1289
rect -6337 1239 -6137 1255
rect -5959 1289 -5759 1327
rect -5959 1255 -5943 1289
rect -5775 1255 -5759 1289
rect -5959 1239 -5759 1255
rect -5581 1289 -5381 1327
rect -5581 1255 -5565 1289
rect -5397 1255 -5381 1289
rect -5581 1239 -5381 1255
rect -5203 1289 -5003 1327
rect -5203 1255 -5187 1289
rect -5019 1255 -5003 1289
rect -5203 1239 -5003 1255
rect -4825 1289 -4625 1327
rect -4825 1255 -4809 1289
rect -4641 1255 -4625 1289
rect -4825 1239 -4625 1255
rect -4447 1289 -4247 1327
rect -4447 1255 -4431 1289
rect -4263 1255 -4247 1289
rect -4447 1239 -4247 1255
rect -4069 1289 -3869 1327
rect -4069 1255 -4053 1289
rect -3885 1255 -3869 1289
rect -4069 1239 -3869 1255
rect -3691 1289 -3491 1327
rect -3691 1255 -3675 1289
rect -3507 1255 -3491 1289
rect -3691 1239 -3491 1255
rect -3313 1289 -3113 1327
rect -3313 1255 -3297 1289
rect -3129 1255 -3113 1289
rect -3313 1239 -3113 1255
rect -2935 1289 -2735 1327
rect -2935 1255 -2919 1289
rect -2751 1255 -2735 1289
rect -2935 1239 -2735 1255
rect -2557 1289 -2357 1327
rect -2557 1255 -2541 1289
rect -2373 1255 -2357 1289
rect -2557 1239 -2357 1255
rect -2179 1289 -1979 1327
rect -2179 1255 -2163 1289
rect -1995 1255 -1979 1289
rect -2179 1239 -1979 1255
rect -1801 1289 -1601 1327
rect -1801 1255 -1785 1289
rect -1617 1255 -1601 1289
rect -1801 1239 -1601 1255
rect -1423 1289 -1223 1327
rect -1423 1255 -1407 1289
rect -1239 1255 -1223 1289
rect -1423 1239 -1223 1255
rect -1045 1289 -845 1327
rect -1045 1255 -1029 1289
rect -861 1255 -845 1289
rect -1045 1239 -845 1255
rect -667 1289 -467 1327
rect -667 1255 -651 1289
rect -483 1255 -467 1289
rect -667 1239 -467 1255
rect -289 1289 -89 1327
rect -289 1255 -273 1289
rect -105 1255 -89 1289
rect -289 1239 -89 1255
rect 89 1289 289 1327
rect 89 1255 105 1289
rect 273 1255 289 1289
rect 89 1239 289 1255
rect 467 1289 667 1327
rect 467 1255 483 1289
rect 651 1255 667 1289
rect 467 1239 667 1255
rect 845 1289 1045 1327
rect 845 1255 861 1289
rect 1029 1255 1045 1289
rect 845 1239 1045 1255
rect 1223 1289 1423 1327
rect 1223 1255 1239 1289
rect 1407 1255 1423 1289
rect 1223 1239 1423 1255
rect 1601 1289 1801 1327
rect 1601 1255 1617 1289
rect 1785 1255 1801 1289
rect 1601 1239 1801 1255
rect 1979 1289 2179 1327
rect 1979 1255 1995 1289
rect 2163 1255 2179 1289
rect 1979 1239 2179 1255
rect 2357 1289 2557 1327
rect 2357 1255 2373 1289
rect 2541 1255 2557 1289
rect 2357 1239 2557 1255
rect 2735 1289 2935 1327
rect 2735 1255 2751 1289
rect 2919 1255 2935 1289
rect 2735 1239 2935 1255
rect 3113 1289 3313 1327
rect 3113 1255 3129 1289
rect 3297 1255 3313 1289
rect 3113 1239 3313 1255
rect 3491 1289 3691 1327
rect 3491 1255 3507 1289
rect 3675 1255 3691 1289
rect 3491 1239 3691 1255
rect 3869 1289 4069 1327
rect 3869 1255 3885 1289
rect 4053 1255 4069 1289
rect 3869 1239 4069 1255
rect 4247 1289 4447 1327
rect 4247 1255 4263 1289
rect 4431 1255 4447 1289
rect 4247 1239 4447 1255
rect 4625 1289 4825 1327
rect 4625 1255 4641 1289
rect 4809 1255 4825 1289
rect 4625 1239 4825 1255
rect 5003 1289 5203 1327
rect 5003 1255 5019 1289
rect 5187 1255 5203 1289
rect 5003 1239 5203 1255
rect 5381 1289 5581 1327
rect 5381 1255 5397 1289
rect 5565 1255 5581 1289
rect 5381 1239 5581 1255
rect 5759 1289 5959 1327
rect 5759 1255 5775 1289
rect 5943 1255 5959 1289
rect 5759 1239 5959 1255
rect 6137 1289 6337 1327
rect 6137 1255 6153 1289
rect 6321 1255 6337 1289
rect 6137 1239 6337 1255
rect 6515 1289 6715 1327
rect 6515 1255 6531 1289
rect 6699 1255 6715 1289
rect 6515 1239 6715 1255
rect 6893 1289 7093 1327
rect 6893 1255 6909 1289
rect 7077 1255 7093 1289
rect 6893 1239 7093 1255
rect 7271 1289 7471 1327
rect 7271 1255 7287 1289
rect 7455 1255 7471 1289
rect 7271 1239 7471 1255
rect 7649 1289 7849 1327
rect 7649 1255 7665 1289
rect 7833 1255 7849 1289
rect 7649 1239 7849 1255
rect 8027 1289 8227 1327
rect 8027 1255 8043 1289
rect 8211 1255 8227 1289
rect 8027 1239 8227 1255
rect 8405 1289 8605 1327
rect 8405 1255 8421 1289
rect 8589 1255 8605 1289
rect 8405 1239 8605 1255
rect 8783 1289 8983 1327
rect 8783 1255 8799 1289
rect 8967 1255 8983 1289
rect 8783 1239 8983 1255
rect 9161 1289 9361 1327
rect 9161 1255 9177 1289
rect 9345 1255 9361 1289
rect 9161 1239 9361 1255
rect -9361 1181 -9161 1197
rect -9361 1147 -9345 1181
rect -9177 1147 -9161 1181
rect -9361 1109 -9161 1147
rect -8983 1181 -8783 1197
rect -8983 1147 -8967 1181
rect -8799 1147 -8783 1181
rect -8983 1109 -8783 1147
rect -8605 1181 -8405 1197
rect -8605 1147 -8589 1181
rect -8421 1147 -8405 1181
rect -8605 1109 -8405 1147
rect -8227 1181 -8027 1197
rect -8227 1147 -8211 1181
rect -8043 1147 -8027 1181
rect -8227 1109 -8027 1147
rect -7849 1181 -7649 1197
rect -7849 1147 -7833 1181
rect -7665 1147 -7649 1181
rect -7849 1109 -7649 1147
rect -7471 1181 -7271 1197
rect -7471 1147 -7455 1181
rect -7287 1147 -7271 1181
rect -7471 1109 -7271 1147
rect -7093 1181 -6893 1197
rect -7093 1147 -7077 1181
rect -6909 1147 -6893 1181
rect -7093 1109 -6893 1147
rect -6715 1181 -6515 1197
rect -6715 1147 -6699 1181
rect -6531 1147 -6515 1181
rect -6715 1109 -6515 1147
rect -6337 1181 -6137 1197
rect -6337 1147 -6321 1181
rect -6153 1147 -6137 1181
rect -6337 1109 -6137 1147
rect -5959 1181 -5759 1197
rect -5959 1147 -5943 1181
rect -5775 1147 -5759 1181
rect -5959 1109 -5759 1147
rect -5581 1181 -5381 1197
rect -5581 1147 -5565 1181
rect -5397 1147 -5381 1181
rect -5581 1109 -5381 1147
rect -5203 1181 -5003 1197
rect -5203 1147 -5187 1181
rect -5019 1147 -5003 1181
rect -5203 1109 -5003 1147
rect -4825 1181 -4625 1197
rect -4825 1147 -4809 1181
rect -4641 1147 -4625 1181
rect -4825 1109 -4625 1147
rect -4447 1181 -4247 1197
rect -4447 1147 -4431 1181
rect -4263 1147 -4247 1181
rect -4447 1109 -4247 1147
rect -4069 1181 -3869 1197
rect -4069 1147 -4053 1181
rect -3885 1147 -3869 1181
rect -4069 1109 -3869 1147
rect -3691 1181 -3491 1197
rect -3691 1147 -3675 1181
rect -3507 1147 -3491 1181
rect -3691 1109 -3491 1147
rect -3313 1181 -3113 1197
rect -3313 1147 -3297 1181
rect -3129 1147 -3113 1181
rect -3313 1109 -3113 1147
rect -2935 1181 -2735 1197
rect -2935 1147 -2919 1181
rect -2751 1147 -2735 1181
rect -2935 1109 -2735 1147
rect -2557 1181 -2357 1197
rect -2557 1147 -2541 1181
rect -2373 1147 -2357 1181
rect -2557 1109 -2357 1147
rect -2179 1181 -1979 1197
rect -2179 1147 -2163 1181
rect -1995 1147 -1979 1181
rect -2179 1109 -1979 1147
rect -1801 1181 -1601 1197
rect -1801 1147 -1785 1181
rect -1617 1147 -1601 1181
rect -1801 1109 -1601 1147
rect -1423 1181 -1223 1197
rect -1423 1147 -1407 1181
rect -1239 1147 -1223 1181
rect -1423 1109 -1223 1147
rect -1045 1181 -845 1197
rect -1045 1147 -1029 1181
rect -861 1147 -845 1181
rect -1045 1109 -845 1147
rect -667 1181 -467 1197
rect -667 1147 -651 1181
rect -483 1147 -467 1181
rect -667 1109 -467 1147
rect -289 1181 -89 1197
rect -289 1147 -273 1181
rect -105 1147 -89 1181
rect -289 1109 -89 1147
rect 89 1181 289 1197
rect 89 1147 105 1181
rect 273 1147 289 1181
rect 89 1109 289 1147
rect 467 1181 667 1197
rect 467 1147 483 1181
rect 651 1147 667 1181
rect 467 1109 667 1147
rect 845 1181 1045 1197
rect 845 1147 861 1181
rect 1029 1147 1045 1181
rect 845 1109 1045 1147
rect 1223 1181 1423 1197
rect 1223 1147 1239 1181
rect 1407 1147 1423 1181
rect 1223 1109 1423 1147
rect 1601 1181 1801 1197
rect 1601 1147 1617 1181
rect 1785 1147 1801 1181
rect 1601 1109 1801 1147
rect 1979 1181 2179 1197
rect 1979 1147 1995 1181
rect 2163 1147 2179 1181
rect 1979 1109 2179 1147
rect 2357 1181 2557 1197
rect 2357 1147 2373 1181
rect 2541 1147 2557 1181
rect 2357 1109 2557 1147
rect 2735 1181 2935 1197
rect 2735 1147 2751 1181
rect 2919 1147 2935 1181
rect 2735 1109 2935 1147
rect 3113 1181 3313 1197
rect 3113 1147 3129 1181
rect 3297 1147 3313 1181
rect 3113 1109 3313 1147
rect 3491 1181 3691 1197
rect 3491 1147 3507 1181
rect 3675 1147 3691 1181
rect 3491 1109 3691 1147
rect 3869 1181 4069 1197
rect 3869 1147 3885 1181
rect 4053 1147 4069 1181
rect 3869 1109 4069 1147
rect 4247 1181 4447 1197
rect 4247 1147 4263 1181
rect 4431 1147 4447 1181
rect 4247 1109 4447 1147
rect 4625 1181 4825 1197
rect 4625 1147 4641 1181
rect 4809 1147 4825 1181
rect 4625 1109 4825 1147
rect 5003 1181 5203 1197
rect 5003 1147 5019 1181
rect 5187 1147 5203 1181
rect 5003 1109 5203 1147
rect 5381 1181 5581 1197
rect 5381 1147 5397 1181
rect 5565 1147 5581 1181
rect 5381 1109 5581 1147
rect 5759 1181 5959 1197
rect 5759 1147 5775 1181
rect 5943 1147 5959 1181
rect 5759 1109 5959 1147
rect 6137 1181 6337 1197
rect 6137 1147 6153 1181
rect 6321 1147 6337 1181
rect 6137 1109 6337 1147
rect 6515 1181 6715 1197
rect 6515 1147 6531 1181
rect 6699 1147 6715 1181
rect 6515 1109 6715 1147
rect 6893 1181 7093 1197
rect 6893 1147 6909 1181
rect 7077 1147 7093 1181
rect 6893 1109 7093 1147
rect 7271 1181 7471 1197
rect 7271 1147 7287 1181
rect 7455 1147 7471 1181
rect 7271 1109 7471 1147
rect 7649 1181 7849 1197
rect 7649 1147 7665 1181
rect 7833 1147 7849 1181
rect 7649 1109 7849 1147
rect 8027 1181 8227 1197
rect 8027 1147 8043 1181
rect 8211 1147 8227 1181
rect 8027 1109 8227 1147
rect 8405 1181 8605 1197
rect 8405 1147 8421 1181
rect 8589 1147 8605 1181
rect 8405 1109 8605 1147
rect 8783 1181 8983 1197
rect 8783 1147 8799 1181
rect 8967 1147 8983 1181
rect 8783 1109 8983 1147
rect 9161 1181 9361 1197
rect 9161 1147 9177 1181
rect 9345 1147 9361 1181
rect 9161 1109 9361 1147
rect -9361 71 -9161 109
rect -9361 37 -9345 71
rect -9177 37 -9161 71
rect -9361 21 -9161 37
rect -8983 71 -8783 109
rect -8983 37 -8967 71
rect -8799 37 -8783 71
rect -8983 21 -8783 37
rect -8605 71 -8405 109
rect -8605 37 -8589 71
rect -8421 37 -8405 71
rect -8605 21 -8405 37
rect -8227 71 -8027 109
rect -8227 37 -8211 71
rect -8043 37 -8027 71
rect -8227 21 -8027 37
rect -7849 71 -7649 109
rect -7849 37 -7833 71
rect -7665 37 -7649 71
rect -7849 21 -7649 37
rect -7471 71 -7271 109
rect -7471 37 -7455 71
rect -7287 37 -7271 71
rect -7471 21 -7271 37
rect -7093 71 -6893 109
rect -7093 37 -7077 71
rect -6909 37 -6893 71
rect -7093 21 -6893 37
rect -6715 71 -6515 109
rect -6715 37 -6699 71
rect -6531 37 -6515 71
rect -6715 21 -6515 37
rect -6337 71 -6137 109
rect -6337 37 -6321 71
rect -6153 37 -6137 71
rect -6337 21 -6137 37
rect -5959 71 -5759 109
rect -5959 37 -5943 71
rect -5775 37 -5759 71
rect -5959 21 -5759 37
rect -5581 71 -5381 109
rect -5581 37 -5565 71
rect -5397 37 -5381 71
rect -5581 21 -5381 37
rect -5203 71 -5003 109
rect -5203 37 -5187 71
rect -5019 37 -5003 71
rect -5203 21 -5003 37
rect -4825 71 -4625 109
rect -4825 37 -4809 71
rect -4641 37 -4625 71
rect -4825 21 -4625 37
rect -4447 71 -4247 109
rect -4447 37 -4431 71
rect -4263 37 -4247 71
rect -4447 21 -4247 37
rect -4069 71 -3869 109
rect -4069 37 -4053 71
rect -3885 37 -3869 71
rect -4069 21 -3869 37
rect -3691 71 -3491 109
rect -3691 37 -3675 71
rect -3507 37 -3491 71
rect -3691 21 -3491 37
rect -3313 71 -3113 109
rect -3313 37 -3297 71
rect -3129 37 -3113 71
rect -3313 21 -3113 37
rect -2935 71 -2735 109
rect -2935 37 -2919 71
rect -2751 37 -2735 71
rect -2935 21 -2735 37
rect -2557 71 -2357 109
rect -2557 37 -2541 71
rect -2373 37 -2357 71
rect -2557 21 -2357 37
rect -2179 71 -1979 109
rect -2179 37 -2163 71
rect -1995 37 -1979 71
rect -2179 21 -1979 37
rect -1801 71 -1601 109
rect -1801 37 -1785 71
rect -1617 37 -1601 71
rect -1801 21 -1601 37
rect -1423 71 -1223 109
rect -1423 37 -1407 71
rect -1239 37 -1223 71
rect -1423 21 -1223 37
rect -1045 71 -845 109
rect -1045 37 -1029 71
rect -861 37 -845 71
rect -1045 21 -845 37
rect -667 71 -467 109
rect -667 37 -651 71
rect -483 37 -467 71
rect -667 21 -467 37
rect -289 71 -89 109
rect -289 37 -273 71
rect -105 37 -89 71
rect -289 21 -89 37
rect 89 71 289 109
rect 89 37 105 71
rect 273 37 289 71
rect 89 21 289 37
rect 467 71 667 109
rect 467 37 483 71
rect 651 37 667 71
rect 467 21 667 37
rect 845 71 1045 109
rect 845 37 861 71
rect 1029 37 1045 71
rect 845 21 1045 37
rect 1223 71 1423 109
rect 1223 37 1239 71
rect 1407 37 1423 71
rect 1223 21 1423 37
rect 1601 71 1801 109
rect 1601 37 1617 71
rect 1785 37 1801 71
rect 1601 21 1801 37
rect 1979 71 2179 109
rect 1979 37 1995 71
rect 2163 37 2179 71
rect 1979 21 2179 37
rect 2357 71 2557 109
rect 2357 37 2373 71
rect 2541 37 2557 71
rect 2357 21 2557 37
rect 2735 71 2935 109
rect 2735 37 2751 71
rect 2919 37 2935 71
rect 2735 21 2935 37
rect 3113 71 3313 109
rect 3113 37 3129 71
rect 3297 37 3313 71
rect 3113 21 3313 37
rect 3491 71 3691 109
rect 3491 37 3507 71
rect 3675 37 3691 71
rect 3491 21 3691 37
rect 3869 71 4069 109
rect 3869 37 3885 71
rect 4053 37 4069 71
rect 3869 21 4069 37
rect 4247 71 4447 109
rect 4247 37 4263 71
rect 4431 37 4447 71
rect 4247 21 4447 37
rect 4625 71 4825 109
rect 4625 37 4641 71
rect 4809 37 4825 71
rect 4625 21 4825 37
rect 5003 71 5203 109
rect 5003 37 5019 71
rect 5187 37 5203 71
rect 5003 21 5203 37
rect 5381 71 5581 109
rect 5381 37 5397 71
rect 5565 37 5581 71
rect 5381 21 5581 37
rect 5759 71 5959 109
rect 5759 37 5775 71
rect 5943 37 5959 71
rect 5759 21 5959 37
rect 6137 71 6337 109
rect 6137 37 6153 71
rect 6321 37 6337 71
rect 6137 21 6337 37
rect 6515 71 6715 109
rect 6515 37 6531 71
rect 6699 37 6715 71
rect 6515 21 6715 37
rect 6893 71 7093 109
rect 6893 37 6909 71
rect 7077 37 7093 71
rect 6893 21 7093 37
rect 7271 71 7471 109
rect 7271 37 7287 71
rect 7455 37 7471 71
rect 7271 21 7471 37
rect 7649 71 7849 109
rect 7649 37 7665 71
rect 7833 37 7849 71
rect 7649 21 7849 37
rect 8027 71 8227 109
rect 8027 37 8043 71
rect 8211 37 8227 71
rect 8027 21 8227 37
rect 8405 71 8605 109
rect 8405 37 8421 71
rect 8589 37 8605 71
rect 8405 21 8605 37
rect 8783 71 8983 109
rect 8783 37 8799 71
rect 8967 37 8983 71
rect 8783 21 8983 37
rect 9161 71 9361 109
rect 9161 37 9177 71
rect 9345 37 9361 71
rect 9161 21 9361 37
rect -9361 -37 -9161 -21
rect -9361 -71 -9345 -37
rect -9177 -71 -9161 -37
rect -9361 -109 -9161 -71
rect -8983 -37 -8783 -21
rect -8983 -71 -8967 -37
rect -8799 -71 -8783 -37
rect -8983 -109 -8783 -71
rect -8605 -37 -8405 -21
rect -8605 -71 -8589 -37
rect -8421 -71 -8405 -37
rect -8605 -109 -8405 -71
rect -8227 -37 -8027 -21
rect -8227 -71 -8211 -37
rect -8043 -71 -8027 -37
rect -8227 -109 -8027 -71
rect -7849 -37 -7649 -21
rect -7849 -71 -7833 -37
rect -7665 -71 -7649 -37
rect -7849 -109 -7649 -71
rect -7471 -37 -7271 -21
rect -7471 -71 -7455 -37
rect -7287 -71 -7271 -37
rect -7471 -109 -7271 -71
rect -7093 -37 -6893 -21
rect -7093 -71 -7077 -37
rect -6909 -71 -6893 -37
rect -7093 -109 -6893 -71
rect -6715 -37 -6515 -21
rect -6715 -71 -6699 -37
rect -6531 -71 -6515 -37
rect -6715 -109 -6515 -71
rect -6337 -37 -6137 -21
rect -6337 -71 -6321 -37
rect -6153 -71 -6137 -37
rect -6337 -109 -6137 -71
rect -5959 -37 -5759 -21
rect -5959 -71 -5943 -37
rect -5775 -71 -5759 -37
rect -5959 -109 -5759 -71
rect -5581 -37 -5381 -21
rect -5581 -71 -5565 -37
rect -5397 -71 -5381 -37
rect -5581 -109 -5381 -71
rect -5203 -37 -5003 -21
rect -5203 -71 -5187 -37
rect -5019 -71 -5003 -37
rect -5203 -109 -5003 -71
rect -4825 -37 -4625 -21
rect -4825 -71 -4809 -37
rect -4641 -71 -4625 -37
rect -4825 -109 -4625 -71
rect -4447 -37 -4247 -21
rect -4447 -71 -4431 -37
rect -4263 -71 -4247 -37
rect -4447 -109 -4247 -71
rect -4069 -37 -3869 -21
rect -4069 -71 -4053 -37
rect -3885 -71 -3869 -37
rect -4069 -109 -3869 -71
rect -3691 -37 -3491 -21
rect -3691 -71 -3675 -37
rect -3507 -71 -3491 -37
rect -3691 -109 -3491 -71
rect -3313 -37 -3113 -21
rect -3313 -71 -3297 -37
rect -3129 -71 -3113 -37
rect -3313 -109 -3113 -71
rect -2935 -37 -2735 -21
rect -2935 -71 -2919 -37
rect -2751 -71 -2735 -37
rect -2935 -109 -2735 -71
rect -2557 -37 -2357 -21
rect -2557 -71 -2541 -37
rect -2373 -71 -2357 -37
rect -2557 -109 -2357 -71
rect -2179 -37 -1979 -21
rect -2179 -71 -2163 -37
rect -1995 -71 -1979 -37
rect -2179 -109 -1979 -71
rect -1801 -37 -1601 -21
rect -1801 -71 -1785 -37
rect -1617 -71 -1601 -37
rect -1801 -109 -1601 -71
rect -1423 -37 -1223 -21
rect -1423 -71 -1407 -37
rect -1239 -71 -1223 -37
rect -1423 -109 -1223 -71
rect -1045 -37 -845 -21
rect -1045 -71 -1029 -37
rect -861 -71 -845 -37
rect -1045 -109 -845 -71
rect -667 -37 -467 -21
rect -667 -71 -651 -37
rect -483 -71 -467 -37
rect -667 -109 -467 -71
rect -289 -37 -89 -21
rect -289 -71 -273 -37
rect -105 -71 -89 -37
rect -289 -109 -89 -71
rect 89 -37 289 -21
rect 89 -71 105 -37
rect 273 -71 289 -37
rect 89 -109 289 -71
rect 467 -37 667 -21
rect 467 -71 483 -37
rect 651 -71 667 -37
rect 467 -109 667 -71
rect 845 -37 1045 -21
rect 845 -71 861 -37
rect 1029 -71 1045 -37
rect 845 -109 1045 -71
rect 1223 -37 1423 -21
rect 1223 -71 1239 -37
rect 1407 -71 1423 -37
rect 1223 -109 1423 -71
rect 1601 -37 1801 -21
rect 1601 -71 1617 -37
rect 1785 -71 1801 -37
rect 1601 -109 1801 -71
rect 1979 -37 2179 -21
rect 1979 -71 1995 -37
rect 2163 -71 2179 -37
rect 1979 -109 2179 -71
rect 2357 -37 2557 -21
rect 2357 -71 2373 -37
rect 2541 -71 2557 -37
rect 2357 -109 2557 -71
rect 2735 -37 2935 -21
rect 2735 -71 2751 -37
rect 2919 -71 2935 -37
rect 2735 -109 2935 -71
rect 3113 -37 3313 -21
rect 3113 -71 3129 -37
rect 3297 -71 3313 -37
rect 3113 -109 3313 -71
rect 3491 -37 3691 -21
rect 3491 -71 3507 -37
rect 3675 -71 3691 -37
rect 3491 -109 3691 -71
rect 3869 -37 4069 -21
rect 3869 -71 3885 -37
rect 4053 -71 4069 -37
rect 3869 -109 4069 -71
rect 4247 -37 4447 -21
rect 4247 -71 4263 -37
rect 4431 -71 4447 -37
rect 4247 -109 4447 -71
rect 4625 -37 4825 -21
rect 4625 -71 4641 -37
rect 4809 -71 4825 -37
rect 4625 -109 4825 -71
rect 5003 -37 5203 -21
rect 5003 -71 5019 -37
rect 5187 -71 5203 -37
rect 5003 -109 5203 -71
rect 5381 -37 5581 -21
rect 5381 -71 5397 -37
rect 5565 -71 5581 -37
rect 5381 -109 5581 -71
rect 5759 -37 5959 -21
rect 5759 -71 5775 -37
rect 5943 -71 5959 -37
rect 5759 -109 5959 -71
rect 6137 -37 6337 -21
rect 6137 -71 6153 -37
rect 6321 -71 6337 -37
rect 6137 -109 6337 -71
rect 6515 -37 6715 -21
rect 6515 -71 6531 -37
rect 6699 -71 6715 -37
rect 6515 -109 6715 -71
rect 6893 -37 7093 -21
rect 6893 -71 6909 -37
rect 7077 -71 7093 -37
rect 6893 -109 7093 -71
rect 7271 -37 7471 -21
rect 7271 -71 7287 -37
rect 7455 -71 7471 -37
rect 7271 -109 7471 -71
rect 7649 -37 7849 -21
rect 7649 -71 7665 -37
rect 7833 -71 7849 -37
rect 7649 -109 7849 -71
rect 8027 -37 8227 -21
rect 8027 -71 8043 -37
rect 8211 -71 8227 -37
rect 8027 -109 8227 -71
rect 8405 -37 8605 -21
rect 8405 -71 8421 -37
rect 8589 -71 8605 -37
rect 8405 -109 8605 -71
rect 8783 -37 8983 -21
rect 8783 -71 8799 -37
rect 8967 -71 8983 -37
rect 8783 -109 8983 -71
rect 9161 -37 9361 -21
rect 9161 -71 9177 -37
rect 9345 -71 9361 -37
rect 9161 -109 9361 -71
rect -9361 -1147 -9161 -1109
rect -9361 -1181 -9345 -1147
rect -9177 -1181 -9161 -1147
rect -9361 -1197 -9161 -1181
rect -8983 -1147 -8783 -1109
rect -8983 -1181 -8967 -1147
rect -8799 -1181 -8783 -1147
rect -8983 -1197 -8783 -1181
rect -8605 -1147 -8405 -1109
rect -8605 -1181 -8589 -1147
rect -8421 -1181 -8405 -1147
rect -8605 -1197 -8405 -1181
rect -8227 -1147 -8027 -1109
rect -8227 -1181 -8211 -1147
rect -8043 -1181 -8027 -1147
rect -8227 -1197 -8027 -1181
rect -7849 -1147 -7649 -1109
rect -7849 -1181 -7833 -1147
rect -7665 -1181 -7649 -1147
rect -7849 -1197 -7649 -1181
rect -7471 -1147 -7271 -1109
rect -7471 -1181 -7455 -1147
rect -7287 -1181 -7271 -1147
rect -7471 -1197 -7271 -1181
rect -7093 -1147 -6893 -1109
rect -7093 -1181 -7077 -1147
rect -6909 -1181 -6893 -1147
rect -7093 -1197 -6893 -1181
rect -6715 -1147 -6515 -1109
rect -6715 -1181 -6699 -1147
rect -6531 -1181 -6515 -1147
rect -6715 -1197 -6515 -1181
rect -6337 -1147 -6137 -1109
rect -6337 -1181 -6321 -1147
rect -6153 -1181 -6137 -1147
rect -6337 -1197 -6137 -1181
rect -5959 -1147 -5759 -1109
rect -5959 -1181 -5943 -1147
rect -5775 -1181 -5759 -1147
rect -5959 -1197 -5759 -1181
rect -5581 -1147 -5381 -1109
rect -5581 -1181 -5565 -1147
rect -5397 -1181 -5381 -1147
rect -5581 -1197 -5381 -1181
rect -5203 -1147 -5003 -1109
rect -5203 -1181 -5187 -1147
rect -5019 -1181 -5003 -1147
rect -5203 -1197 -5003 -1181
rect -4825 -1147 -4625 -1109
rect -4825 -1181 -4809 -1147
rect -4641 -1181 -4625 -1147
rect -4825 -1197 -4625 -1181
rect -4447 -1147 -4247 -1109
rect -4447 -1181 -4431 -1147
rect -4263 -1181 -4247 -1147
rect -4447 -1197 -4247 -1181
rect -4069 -1147 -3869 -1109
rect -4069 -1181 -4053 -1147
rect -3885 -1181 -3869 -1147
rect -4069 -1197 -3869 -1181
rect -3691 -1147 -3491 -1109
rect -3691 -1181 -3675 -1147
rect -3507 -1181 -3491 -1147
rect -3691 -1197 -3491 -1181
rect -3313 -1147 -3113 -1109
rect -3313 -1181 -3297 -1147
rect -3129 -1181 -3113 -1147
rect -3313 -1197 -3113 -1181
rect -2935 -1147 -2735 -1109
rect -2935 -1181 -2919 -1147
rect -2751 -1181 -2735 -1147
rect -2935 -1197 -2735 -1181
rect -2557 -1147 -2357 -1109
rect -2557 -1181 -2541 -1147
rect -2373 -1181 -2357 -1147
rect -2557 -1197 -2357 -1181
rect -2179 -1147 -1979 -1109
rect -2179 -1181 -2163 -1147
rect -1995 -1181 -1979 -1147
rect -2179 -1197 -1979 -1181
rect -1801 -1147 -1601 -1109
rect -1801 -1181 -1785 -1147
rect -1617 -1181 -1601 -1147
rect -1801 -1197 -1601 -1181
rect -1423 -1147 -1223 -1109
rect -1423 -1181 -1407 -1147
rect -1239 -1181 -1223 -1147
rect -1423 -1197 -1223 -1181
rect -1045 -1147 -845 -1109
rect -1045 -1181 -1029 -1147
rect -861 -1181 -845 -1147
rect -1045 -1197 -845 -1181
rect -667 -1147 -467 -1109
rect -667 -1181 -651 -1147
rect -483 -1181 -467 -1147
rect -667 -1197 -467 -1181
rect -289 -1147 -89 -1109
rect -289 -1181 -273 -1147
rect -105 -1181 -89 -1147
rect -289 -1197 -89 -1181
rect 89 -1147 289 -1109
rect 89 -1181 105 -1147
rect 273 -1181 289 -1147
rect 89 -1197 289 -1181
rect 467 -1147 667 -1109
rect 467 -1181 483 -1147
rect 651 -1181 667 -1147
rect 467 -1197 667 -1181
rect 845 -1147 1045 -1109
rect 845 -1181 861 -1147
rect 1029 -1181 1045 -1147
rect 845 -1197 1045 -1181
rect 1223 -1147 1423 -1109
rect 1223 -1181 1239 -1147
rect 1407 -1181 1423 -1147
rect 1223 -1197 1423 -1181
rect 1601 -1147 1801 -1109
rect 1601 -1181 1617 -1147
rect 1785 -1181 1801 -1147
rect 1601 -1197 1801 -1181
rect 1979 -1147 2179 -1109
rect 1979 -1181 1995 -1147
rect 2163 -1181 2179 -1147
rect 1979 -1197 2179 -1181
rect 2357 -1147 2557 -1109
rect 2357 -1181 2373 -1147
rect 2541 -1181 2557 -1147
rect 2357 -1197 2557 -1181
rect 2735 -1147 2935 -1109
rect 2735 -1181 2751 -1147
rect 2919 -1181 2935 -1147
rect 2735 -1197 2935 -1181
rect 3113 -1147 3313 -1109
rect 3113 -1181 3129 -1147
rect 3297 -1181 3313 -1147
rect 3113 -1197 3313 -1181
rect 3491 -1147 3691 -1109
rect 3491 -1181 3507 -1147
rect 3675 -1181 3691 -1147
rect 3491 -1197 3691 -1181
rect 3869 -1147 4069 -1109
rect 3869 -1181 3885 -1147
rect 4053 -1181 4069 -1147
rect 3869 -1197 4069 -1181
rect 4247 -1147 4447 -1109
rect 4247 -1181 4263 -1147
rect 4431 -1181 4447 -1147
rect 4247 -1197 4447 -1181
rect 4625 -1147 4825 -1109
rect 4625 -1181 4641 -1147
rect 4809 -1181 4825 -1147
rect 4625 -1197 4825 -1181
rect 5003 -1147 5203 -1109
rect 5003 -1181 5019 -1147
rect 5187 -1181 5203 -1147
rect 5003 -1197 5203 -1181
rect 5381 -1147 5581 -1109
rect 5381 -1181 5397 -1147
rect 5565 -1181 5581 -1147
rect 5381 -1197 5581 -1181
rect 5759 -1147 5959 -1109
rect 5759 -1181 5775 -1147
rect 5943 -1181 5959 -1147
rect 5759 -1197 5959 -1181
rect 6137 -1147 6337 -1109
rect 6137 -1181 6153 -1147
rect 6321 -1181 6337 -1147
rect 6137 -1197 6337 -1181
rect 6515 -1147 6715 -1109
rect 6515 -1181 6531 -1147
rect 6699 -1181 6715 -1147
rect 6515 -1197 6715 -1181
rect 6893 -1147 7093 -1109
rect 6893 -1181 6909 -1147
rect 7077 -1181 7093 -1147
rect 6893 -1197 7093 -1181
rect 7271 -1147 7471 -1109
rect 7271 -1181 7287 -1147
rect 7455 -1181 7471 -1147
rect 7271 -1197 7471 -1181
rect 7649 -1147 7849 -1109
rect 7649 -1181 7665 -1147
rect 7833 -1181 7849 -1147
rect 7649 -1197 7849 -1181
rect 8027 -1147 8227 -1109
rect 8027 -1181 8043 -1147
rect 8211 -1181 8227 -1147
rect 8027 -1197 8227 -1181
rect 8405 -1147 8605 -1109
rect 8405 -1181 8421 -1147
rect 8589 -1181 8605 -1147
rect 8405 -1197 8605 -1181
rect 8783 -1147 8983 -1109
rect 8783 -1181 8799 -1147
rect 8967 -1181 8983 -1147
rect 8783 -1197 8983 -1181
rect 9161 -1147 9361 -1109
rect 9161 -1181 9177 -1147
rect 9345 -1181 9361 -1147
rect 9161 -1197 9361 -1181
rect -9361 -1255 -9161 -1239
rect -9361 -1289 -9345 -1255
rect -9177 -1289 -9161 -1255
rect -9361 -1327 -9161 -1289
rect -8983 -1255 -8783 -1239
rect -8983 -1289 -8967 -1255
rect -8799 -1289 -8783 -1255
rect -8983 -1327 -8783 -1289
rect -8605 -1255 -8405 -1239
rect -8605 -1289 -8589 -1255
rect -8421 -1289 -8405 -1255
rect -8605 -1327 -8405 -1289
rect -8227 -1255 -8027 -1239
rect -8227 -1289 -8211 -1255
rect -8043 -1289 -8027 -1255
rect -8227 -1327 -8027 -1289
rect -7849 -1255 -7649 -1239
rect -7849 -1289 -7833 -1255
rect -7665 -1289 -7649 -1255
rect -7849 -1327 -7649 -1289
rect -7471 -1255 -7271 -1239
rect -7471 -1289 -7455 -1255
rect -7287 -1289 -7271 -1255
rect -7471 -1327 -7271 -1289
rect -7093 -1255 -6893 -1239
rect -7093 -1289 -7077 -1255
rect -6909 -1289 -6893 -1255
rect -7093 -1327 -6893 -1289
rect -6715 -1255 -6515 -1239
rect -6715 -1289 -6699 -1255
rect -6531 -1289 -6515 -1255
rect -6715 -1327 -6515 -1289
rect -6337 -1255 -6137 -1239
rect -6337 -1289 -6321 -1255
rect -6153 -1289 -6137 -1255
rect -6337 -1327 -6137 -1289
rect -5959 -1255 -5759 -1239
rect -5959 -1289 -5943 -1255
rect -5775 -1289 -5759 -1255
rect -5959 -1327 -5759 -1289
rect -5581 -1255 -5381 -1239
rect -5581 -1289 -5565 -1255
rect -5397 -1289 -5381 -1255
rect -5581 -1327 -5381 -1289
rect -5203 -1255 -5003 -1239
rect -5203 -1289 -5187 -1255
rect -5019 -1289 -5003 -1255
rect -5203 -1327 -5003 -1289
rect -4825 -1255 -4625 -1239
rect -4825 -1289 -4809 -1255
rect -4641 -1289 -4625 -1255
rect -4825 -1327 -4625 -1289
rect -4447 -1255 -4247 -1239
rect -4447 -1289 -4431 -1255
rect -4263 -1289 -4247 -1255
rect -4447 -1327 -4247 -1289
rect -4069 -1255 -3869 -1239
rect -4069 -1289 -4053 -1255
rect -3885 -1289 -3869 -1255
rect -4069 -1327 -3869 -1289
rect -3691 -1255 -3491 -1239
rect -3691 -1289 -3675 -1255
rect -3507 -1289 -3491 -1255
rect -3691 -1327 -3491 -1289
rect -3313 -1255 -3113 -1239
rect -3313 -1289 -3297 -1255
rect -3129 -1289 -3113 -1255
rect -3313 -1327 -3113 -1289
rect -2935 -1255 -2735 -1239
rect -2935 -1289 -2919 -1255
rect -2751 -1289 -2735 -1255
rect -2935 -1327 -2735 -1289
rect -2557 -1255 -2357 -1239
rect -2557 -1289 -2541 -1255
rect -2373 -1289 -2357 -1255
rect -2557 -1327 -2357 -1289
rect -2179 -1255 -1979 -1239
rect -2179 -1289 -2163 -1255
rect -1995 -1289 -1979 -1255
rect -2179 -1327 -1979 -1289
rect -1801 -1255 -1601 -1239
rect -1801 -1289 -1785 -1255
rect -1617 -1289 -1601 -1255
rect -1801 -1327 -1601 -1289
rect -1423 -1255 -1223 -1239
rect -1423 -1289 -1407 -1255
rect -1239 -1289 -1223 -1255
rect -1423 -1327 -1223 -1289
rect -1045 -1255 -845 -1239
rect -1045 -1289 -1029 -1255
rect -861 -1289 -845 -1255
rect -1045 -1327 -845 -1289
rect -667 -1255 -467 -1239
rect -667 -1289 -651 -1255
rect -483 -1289 -467 -1255
rect -667 -1327 -467 -1289
rect -289 -1255 -89 -1239
rect -289 -1289 -273 -1255
rect -105 -1289 -89 -1255
rect -289 -1327 -89 -1289
rect 89 -1255 289 -1239
rect 89 -1289 105 -1255
rect 273 -1289 289 -1255
rect 89 -1327 289 -1289
rect 467 -1255 667 -1239
rect 467 -1289 483 -1255
rect 651 -1289 667 -1255
rect 467 -1327 667 -1289
rect 845 -1255 1045 -1239
rect 845 -1289 861 -1255
rect 1029 -1289 1045 -1255
rect 845 -1327 1045 -1289
rect 1223 -1255 1423 -1239
rect 1223 -1289 1239 -1255
rect 1407 -1289 1423 -1255
rect 1223 -1327 1423 -1289
rect 1601 -1255 1801 -1239
rect 1601 -1289 1617 -1255
rect 1785 -1289 1801 -1255
rect 1601 -1327 1801 -1289
rect 1979 -1255 2179 -1239
rect 1979 -1289 1995 -1255
rect 2163 -1289 2179 -1255
rect 1979 -1327 2179 -1289
rect 2357 -1255 2557 -1239
rect 2357 -1289 2373 -1255
rect 2541 -1289 2557 -1255
rect 2357 -1327 2557 -1289
rect 2735 -1255 2935 -1239
rect 2735 -1289 2751 -1255
rect 2919 -1289 2935 -1255
rect 2735 -1327 2935 -1289
rect 3113 -1255 3313 -1239
rect 3113 -1289 3129 -1255
rect 3297 -1289 3313 -1255
rect 3113 -1327 3313 -1289
rect 3491 -1255 3691 -1239
rect 3491 -1289 3507 -1255
rect 3675 -1289 3691 -1255
rect 3491 -1327 3691 -1289
rect 3869 -1255 4069 -1239
rect 3869 -1289 3885 -1255
rect 4053 -1289 4069 -1255
rect 3869 -1327 4069 -1289
rect 4247 -1255 4447 -1239
rect 4247 -1289 4263 -1255
rect 4431 -1289 4447 -1255
rect 4247 -1327 4447 -1289
rect 4625 -1255 4825 -1239
rect 4625 -1289 4641 -1255
rect 4809 -1289 4825 -1255
rect 4625 -1327 4825 -1289
rect 5003 -1255 5203 -1239
rect 5003 -1289 5019 -1255
rect 5187 -1289 5203 -1255
rect 5003 -1327 5203 -1289
rect 5381 -1255 5581 -1239
rect 5381 -1289 5397 -1255
rect 5565 -1289 5581 -1255
rect 5381 -1327 5581 -1289
rect 5759 -1255 5959 -1239
rect 5759 -1289 5775 -1255
rect 5943 -1289 5959 -1255
rect 5759 -1327 5959 -1289
rect 6137 -1255 6337 -1239
rect 6137 -1289 6153 -1255
rect 6321 -1289 6337 -1255
rect 6137 -1327 6337 -1289
rect 6515 -1255 6715 -1239
rect 6515 -1289 6531 -1255
rect 6699 -1289 6715 -1255
rect 6515 -1327 6715 -1289
rect 6893 -1255 7093 -1239
rect 6893 -1289 6909 -1255
rect 7077 -1289 7093 -1255
rect 6893 -1327 7093 -1289
rect 7271 -1255 7471 -1239
rect 7271 -1289 7287 -1255
rect 7455 -1289 7471 -1255
rect 7271 -1327 7471 -1289
rect 7649 -1255 7849 -1239
rect 7649 -1289 7665 -1255
rect 7833 -1289 7849 -1255
rect 7649 -1327 7849 -1289
rect 8027 -1255 8227 -1239
rect 8027 -1289 8043 -1255
rect 8211 -1289 8227 -1255
rect 8027 -1327 8227 -1289
rect 8405 -1255 8605 -1239
rect 8405 -1289 8421 -1255
rect 8589 -1289 8605 -1255
rect 8405 -1327 8605 -1289
rect 8783 -1255 8983 -1239
rect 8783 -1289 8799 -1255
rect 8967 -1289 8983 -1255
rect 8783 -1327 8983 -1289
rect 9161 -1255 9361 -1239
rect 9161 -1289 9177 -1255
rect 9345 -1289 9361 -1255
rect 9161 -1327 9361 -1289
rect -9361 -2365 -9161 -2327
rect -9361 -2399 -9345 -2365
rect -9177 -2399 -9161 -2365
rect -9361 -2415 -9161 -2399
rect -8983 -2365 -8783 -2327
rect -8983 -2399 -8967 -2365
rect -8799 -2399 -8783 -2365
rect -8983 -2415 -8783 -2399
rect -8605 -2365 -8405 -2327
rect -8605 -2399 -8589 -2365
rect -8421 -2399 -8405 -2365
rect -8605 -2415 -8405 -2399
rect -8227 -2365 -8027 -2327
rect -8227 -2399 -8211 -2365
rect -8043 -2399 -8027 -2365
rect -8227 -2415 -8027 -2399
rect -7849 -2365 -7649 -2327
rect -7849 -2399 -7833 -2365
rect -7665 -2399 -7649 -2365
rect -7849 -2415 -7649 -2399
rect -7471 -2365 -7271 -2327
rect -7471 -2399 -7455 -2365
rect -7287 -2399 -7271 -2365
rect -7471 -2415 -7271 -2399
rect -7093 -2365 -6893 -2327
rect -7093 -2399 -7077 -2365
rect -6909 -2399 -6893 -2365
rect -7093 -2415 -6893 -2399
rect -6715 -2365 -6515 -2327
rect -6715 -2399 -6699 -2365
rect -6531 -2399 -6515 -2365
rect -6715 -2415 -6515 -2399
rect -6337 -2365 -6137 -2327
rect -6337 -2399 -6321 -2365
rect -6153 -2399 -6137 -2365
rect -6337 -2415 -6137 -2399
rect -5959 -2365 -5759 -2327
rect -5959 -2399 -5943 -2365
rect -5775 -2399 -5759 -2365
rect -5959 -2415 -5759 -2399
rect -5581 -2365 -5381 -2327
rect -5581 -2399 -5565 -2365
rect -5397 -2399 -5381 -2365
rect -5581 -2415 -5381 -2399
rect -5203 -2365 -5003 -2327
rect -5203 -2399 -5187 -2365
rect -5019 -2399 -5003 -2365
rect -5203 -2415 -5003 -2399
rect -4825 -2365 -4625 -2327
rect -4825 -2399 -4809 -2365
rect -4641 -2399 -4625 -2365
rect -4825 -2415 -4625 -2399
rect -4447 -2365 -4247 -2327
rect -4447 -2399 -4431 -2365
rect -4263 -2399 -4247 -2365
rect -4447 -2415 -4247 -2399
rect -4069 -2365 -3869 -2327
rect -4069 -2399 -4053 -2365
rect -3885 -2399 -3869 -2365
rect -4069 -2415 -3869 -2399
rect -3691 -2365 -3491 -2327
rect -3691 -2399 -3675 -2365
rect -3507 -2399 -3491 -2365
rect -3691 -2415 -3491 -2399
rect -3313 -2365 -3113 -2327
rect -3313 -2399 -3297 -2365
rect -3129 -2399 -3113 -2365
rect -3313 -2415 -3113 -2399
rect -2935 -2365 -2735 -2327
rect -2935 -2399 -2919 -2365
rect -2751 -2399 -2735 -2365
rect -2935 -2415 -2735 -2399
rect -2557 -2365 -2357 -2327
rect -2557 -2399 -2541 -2365
rect -2373 -2399 -2357 -2365
rect -2557 -2415 -2357 -2399
rect -2179 -2365 -1979 -2327
rect -2179 -2399 -2163 -2365
rect -1995 -2399 -1979 -2365
rect -2179 -2415 -1979 -2399
rect -1801 -2365 -1601 -2327
rect -1801 -2399 -1785 -2365
rect -1617 -2399 -1601 -2365
rect -1801 -2415 -1601 -2399
rect -1423 -2365 -1223 -2327
rect -1423 -2399 -1407 -2365
rect -1239 -2399 -1223 -2365
rect -1423 -2415 -1223 -2399
rect -1045 -2365 -845 -2327
rect -1045 -2399 -1029 -2365
rect -861 -2399 -845 -2365
rect -1045 -2415 -845 -2399
rect -667 -2365 -467 -2327
rect -667 -2399 -651 -2365
rect -483 -2399 -467 -2365
rect -667 -2415 -467 -2399
rect -289 -2365 -89 -2327
rect -289 -2399 -273 -2365
rect -105 -2399 -89 -2365
rect -289 -2415 -89 -2399
rect 89 -2365 289 -2327
rect 89 -2399 105 -2365
rect 273 -2399 289 -2365
rect 89 -2415 289 -2399
rect 467 -2365 667 -2327
rect 467 -2399 483 -2365
rect 651 -2399 667 -2365
rect 467 -2415 667 -2399
rect 845 -2365 1045 -2327
rect 845 -2399 861 -2365
rect 1029 -2399 1045 -2365
rect 845 -2415 1045 -2399
rect 1223 -2365 1423 -2327
rect 1223 -2399 1239 -2365
rect 1407 -2399 1423 -2365
rect 1223 -2415 1423 -2399
rect 1601 -2365 1801 -2327
rect 1601 -2399 1617 -2365
rect 1785 -2399 1801 -2365
rect 1601 -2415 1801 -2399
rect 1979 -2365 2179 -2327
rect 1979 -2399 1995 -2365
rect 2163 -2399 2179 -2365
rect 1979 -2415 2179 -2399
rect 2357 -2365 2557 -2327
rect 2357 -2399 2373 -2365
rect 2541 -2399 2557 -2365
rect 2357 -2415 2557 -2399
rect 2735 -2365 2935 -2327
rect 2735 -2399 2751 -2365
rect 2919 -2399 2935 -2365
rect 2735 -2415 2935 -2399
rect 3113 -2365 3313 -2327
rect 3113 -2399 3129 -2365
rect 3297 -2399 3313 -2365
rect 3113 -2415 3313 -2399
rect 3491 -2365 3691 -2327
rect 3491 -2399 3507 -2365
rect 3675 -2399 3691 -2365
rect 3491 -2415 3691 -2399
rect 3869 -2365 4069 -2327
rect 3869 -2399 3885 -2365
rect 4053 -2399 4069 -2365
rect 3869 -2415 4069 -2399
rect 4247 -2365 4447 -2327
rect 4247 -2399 4263 -2365
rect 4431 -2399 4447 -2365
rect 4247 -2415 4447 -2399
rect 4625 -2365 4825 -2327
rect 4625 -2399 4641 -2365
rect 4809 -2399 4825 -2365
rect 4625 -2415 4825 -2399
rect 5003 -2365 5203 -2327
rect 5003 -2399 5019 -2365
rect 5187 -2399 5203 -2365
rect 5003 -2415 5203 -2399
rect 5381 -2365 5581 -2327
rect 5381 -2399 5397 -2365
rect 5565 -2399 5581 -2365
rect 5381 -2415 5581 -2399
rect 5759 -2365 5959 -2327
rect 5759 -2399 5775 -2365
rect 5943 -2399 5959 -2365
rect 5759 -2415 5959 -2399
rect 6137 -2365 6337 -2327
rect 6137 -2399 6153 -2365
rect 6321 -2399 6337 -2365
rect 6137 -2415 6337 -2399
rect 6515 -2365 6715 -2327
rect 6515 -2399 6531 -2365
rect 6699 -2399 6715 -2365
rect 6515 -2415 6715 -2399
rect 6893 -2365 7093 -2327
rect 6893 -2399 6909 -2365
rect 7077 -2399 7093 -2365
rect 6893 -2415 7093 -2399
rect 7271 -2365 7471 -2327
rect 7271 -2399 7287 -2365
rect 7455 -2399 7471 -2365
rect 7271 -2415 7471 -2399
rect 7649 -2365 7849 -2327
rect 7649 -2399 7665 -2365
rect 7833 -2399 7849 -2365
rect 7649 -2415 7849 -2399
rect 8027 -2365 8227 -2327
rect 8027 -2399 8043 -2365
rect 8211 -2399 8227 -2365
rect 8027 -2415 8227 -2399
rect 8405 -2365 8605 -2327
rect 8405 -2399 8421 -2365
rect 8589 -2399 8605 -2365
rect 8405 -2415 8605 -2399
rect 8783 -2365 8983 -2327
rect 8783 -2399 8799 -2365
rect 8967 -2399 8983 -2365
rect 8783 -2415 8983 -2399
rect 9161 -2365 9361 -2327
rect 9161 -2399 9177 -2365
rect 9345 -2399 9361 -2365
rect 9161 -2415 9361 -2399
<< polycont >>
rect -9345 2365 -9177 2399
rect -8967 2365 -8799 2399
rect -8589 2365 -8421 2399
rect -8211 2365 -8043 2399
rect -7833 2365 -7665 2399
rect -7455 2365 -7287 2399
rect -7077 2365 -6909 2399
rect -6699 2365 -6531 2399
rect -6321 2365 -6153 2399
rect -5943 2365 -5775 2399
rect -5565 2365 -5397 2399
rect -5187 2365 -5019 2399
rect -4809 2365 -4641 2399
rect -4431 2365 -4263 2399
rect -4053 2365 -3885 2399
rect -3675 2365 -3507 2399
rect -3297 2365 -3129 2399
rect -2919 2365 -2751 2399
rect -2541 2365 -2373 2399
rect -2163 2365 -1995 2399
rect -1785 2365 -1617 2399
rect -1407 2365 -1239 2399
rect -1029 2365 -861 2399
rect -651 2365 -483 2399
rect -273 2365 -105 2399
rect 105 2365 273 2399
rect 483 2365 651 2399
rect 861 2365 1029 2399
rect 1239 2365 1407 2399
rect 1617 2365 1785 2399
rect 1995 2365 2163 2399
rect 2373 2365 2541 2399
rect 2751 2365 2919 2399
rect 3129 2365 3297 2399
rect 3507 2365 3675 2399
rect 3885 2365 4053 2399
rect 4263 2365 4431 2399
rect 4641 2365 4809 2399
rect 5019 2365 5187 2399
rect 5397 2365 5565 2399
rect 5775 2365 5943 2399
rect 6153 2365 6321 2399
rect 6531 2365 6699 2399
rect 6909 2365 7077 2399
rect 7287 2365 7455 2399
rect 7665 2365 7833 2399
rect 8043 2365 8211 2399
rect 8421 2365 8589 2399
rect 8799 2365 8967 2399
rect 9177 2365 9345 2399
rect -9345 1255 -9177 1289
rect -8967 1255 -8799 1289
rect -8589 1255 -8421 1289
rect -8211 1255 -8043 1289
rect -7833 1255 -7665 1289
rect -7455 1255 -7287 1289
rect -7077 1255 -6909 1289
rect -6699 1255 -6531 1289
rect -6321 1255 -6153 1289
rect -5943 1255 -5775 1289
rect -5565 1255 -5397 1289
rect -5187 1255 -5019 1289
rect -4809 1255 -4641 1289
rect -4431 1255 -4263 1289
rect -4053 1255 -3885 1289
rect -3675 1255 -3507 1289
rect -3297 1255 -3129 1289
rect -2919 1255 -2751 1289
rect -2541 1255 -2373 1289
rect -2163 1255 -1995 1289
rect -1785 1255 -1617 1289
rect -1407 1255 -1239 1289
rect -1029 1255 -861 1289
rect -651 1255 -483 1289
rect -273 1255 -105 1289
rect 105 1255 273 1289
rect 483 1255 651 1289
rect 861 1255 1029 1289
rect 1239 1255 1407 1289
rect 1617 1255 1785 1289
rect 1995 1255 2163 1289
rect 2373 1255 2541 1289
rect 2751 1255 2919 1289
rect 3129 1255 3297 1289
rect 3507 1255 3675 1289
rect 3885 1255 4053 1289
rect 4263 1255 4431 1289
rect 4641 1255 4809 1289
rect 5019 1255 5187 1289
rect 5397 1255 5565 1289
rect 5775 1255 5943 1289
rect 6153 1255 6321 1289
rect 6531 1255 6699 1289
rect 6909 1255 7077 1289
rect 7287 1255 7455 1289
rect 7665 1255 7833 1289
rect 8043 1255 8211 1289
rect 8421 1255 8589 1289
rect 8799 1255 8967 1289
rect 9177 1255 9345 1289
rect -9345 1147 -9177 1181
rect -8967 1147 -8799 1181
rect -8589 1147 -8421 1181
rect -8211 1147 -8043 1181
rect -7833 1147 -7665 1181
rect -7455 1147 -7287 1181
rect -7077 1147 -6909 1181
rect -6699 1147 -6531 1181
rect -6321 1147 -6153 1181
rect -5943 1147 -5775 1181
rect -5565 1147 -5397 1181
rect -5187 1147 -5019 1181
rect -4809 1147 -4641 1181
rect -4431 1147 -4263 1181
rect -4053 1147 -3885 1181
rect -3675 1147 -3507 1181
rect -3297 1147 -3129 1181
rect -2919 1147 -2751 1181
rect -2541 1147 -2373 1181
rect -2163 1147 -1995 1181
rect -1785 1147 -1617 1181
rect -1407 1147 -1239 1181
rect -1029 1147 -861 1181
rect -651 1147 -483 1181
rect -273 1147 -105 1181
rect 105 1147 273 1181
rect 483 1147 651 1181
rect 861 1147 1029 1181
rect 1239 1147 1407 1181
rect 1617 1147 1785 1181
rect 1995 1147 2163 1181
rect 2373 1147 2541 1181
rect 2751 1147 2919 1181
rect 3129 1147 3297 1181
rect 3507 1147 3675 1181
rect 3885 1147 4053 1181
rect 4263 1147 4431 1181
rect 4641 1147 4809 1181
rect 5019 1147 5187 1181
rect 5397 1147 5565 1181
rect 5775 1147 5943 1181
rect 6153 1147 6321 1181
rect 6531 1147 6699 1181
rect 6909 1147 7077 1181
rect 7287 1147 7455 1181
rect 7665 1147 7833 1181
rect 8043 1147 8211 1181
rect 8421 1147 8589 1181
rect 8799 1147 8967 1181
rect 9177 1147 9345 1181
rect -9345 37 -9177 71
rect -8967 37 -8799 71
rect -8589 37 -8421 71
rect -8211 37 -8043 71
rect -7833 37 -7665 71
rect -7455 37 -7287 71
rect -7077 37 -6909 71
rect -6699 37 -6531 71
rect -6321 37 -6153 71
rect -5943 37 -5775 71
rect -5565 37 -5397 71
rect -5187 37 -5019 71
rect -4809 37 -4641 71
rect -4431 37 -4263 71
rect -4053 37 -3885 71
rect -3675 37 -3507 71
rect -3297 37 -3129 71
rect -2919 37 -2751 71
rect -2541 37 -2373 71
rect -2163 37 -1995 71
rect -1785 37 -1617 71
rect -1407 37 -1239 71
rect -1029 37 -861 71
rect -651 37 -483 71
rect -273 37 -105 71
rect 105 37 273 71
rect 483 37 651 71
rect 861 37 1029 71
rect 1239 37 1407 71
rect 1617 37 1785 71
rect 1995 37 2163 71
rect 2373 37 2541 71
rect 2751 37 2919 71
rect 3129 37 3297 71
rect 3507 37 3675 71
rect 3885 37 4053 71
rect 4263 37 4431 71
rect 4641 37 4809 71
rect 5019 37 5187 71
rect 5397 37 5565 71
rect 5775 37 5943 71
rect 6153 37 6321 71
rect 6531 37 6699 71
rect 6909 37 7077 71
rect 7287 37 7455 71
rect 7665 37 7833 71
rect 8043 37 8211 71
rect 8421 37 8589 71
rect 8799 37 8967 71
rect 9177 37 9345 71
rect -9345 -71 -9177 -37
rect -8967 -71 -8799 -37
rect -8589 -71 -8421 -37
rect -8211 -71 -8043 -37
rect -7833 -71 -7665 -37
rect -7455 -71 -7287 -37
rect -7077 -71 -6909 -37
rect -6699 -71 -6531 -37
rect -6321 -71 -6153 -37
rect -5943 -71 -5775 -37
rect -5565 -71 -5397 -37
rect -5187 -71 -5019 -37
rect -4809 -71 -4641 -37
rect -4431 -71 -4263 -37
rect -4053 -71 -3885 -37
rect -3675 -71 -3507 -37
rect -3297 -71 -3129 -37
rect -2919 -71 -2751 -37
rect -2541 -71 -2373 -37
rect -2163 -71 -1995 -37
rect -1785 -71 -1617 -37
rect -1407 -71 -1239 -37
rect -1029 -71 -861 -37
rect -651 -71 -483 -37
rect -273 -71 -105 -37
rect 105 -71 273 -37
rect 483 -71 651 -37
rect 861 -71 1029 -37
rect 1239 -71 1407 -37
rect 1617 -71 1785 -37
rect 1995 -71 2163 -37
rect 2373 -71 2541 -37
rect 2751 -71 2919 -37
rect 3129 -71 3297 -37
rect 3507 -71 3675 -37
rect 3885 -71 4053 -37
rect 4263 -71 4431 -37
rect 4641 -71 4809 -37
rect 5019 -71 5187 -37
rect 5397 -71 5565 -37
rect 5775 -71 5943 -37
rect 6153 -71 6321 -37
rect 6531 -71 6699 -37
rect 6909 -71 7077 -37
rect 7287 -71 7455 -37
rect 7665 -71 7833 -37
rect 8043 -71 8211 -37
rect 8421 -71 8589 -37
rect 8799 -71 8967 -37
rect 9177 -71 9345 -37
rect -9345 -1181 -9177 -1147
rect -8967 -1181 -8799 -1147
rect -8589 -1181 -8421 -1147
rect -8211 -1181 -8043 -1147
rect -7833 -1181 -7665 -1147
rect -7455 -1181 -7287 -1147
rect -7077 -1181 -6909 -1147
rect -6699 -1181 -6531 -1147
rect -6321 -1181 -6153 -1147
rect -5943 -1181 -5775 -1147
rect -5565 -1181 -5397 -1147
rect -5187 -1181 -5019 -1147
rect -4809 -1181 -4641 -1147
rect -4431 -1181 -4263 -1147
rect -4053 -1181 -3885 -1147
rect -3675 -1181 -3507 -1147
rect -3297 -1181 -3129 -1147
rect -2919 -1181 -2751 -1147
rect -2541 -1181 -2373 -1147
rect -2163 -1181 -1995 -1147
rect -1785 -1181 -1617 -1147
rect -1407 -1181 -1239 -1147
rect -1029 -1181 -861 -1147
rect -651 -1181 -483 -1147
rect -273 -1181 -105 -1147
rect 105 -1181 273 -1147
rect 483 -1181 651 -1147
rect 861 -1181 1029 -1147
rect 1239 -1181 1407 -1147
rect 1617 -1181 1785 -1147
rect 1995 -1181 2163 -1147
rect 2373 -1181 2541 -1147
rect 2751 -1181 2919 -1147
rect 3129 -1181 3297 -1147
rect 3507 -1181 3675 -1147
rect 3885 -1181 4053 -1147
rect 4263 -1181 4431 -1147
rect 4641 -1181 4809 -1147
rect 5019 -1181 5187 -1147
rect 5397 -1181 5565 -1147
rect 5775 -1181 5943 -1147
rect 6153 -1181 6321 -1147
rect 6531 -1181 6699 -1147
rect 6909 -1181 7077 -1147
rect 7287 -1181 7455 -1147
rect 7665 -1181 7833 -1147
rect 8043 -1181 8211 -1147
rect 8421 -1181 8589 -1147
rect 8799 -1181 8967 -1147
rect 9177 -1181 9345 -1147
rect -9345 -1289 -9177 -1255
rect -8967 -1289 -8799 -1255
rect -8589 -1289 -8421 -1255
rect -8211 -1289 -8043 -1255
rect -7833 -1289 -7665 -1255
rect -7455 -1289 -7287 -1255
rect -7077 -1289 -6909 -1255
rect -6699 -1289 -6531 -1255
rect -6321 -1289 -6153 -1255
rect -5943 -1289 -5775 -1255
rect -5565 -1289 -5397 -1255
rect -5187 -1289 -5019 -1255
rect -4809 -1289 -4641 -1255
rect -4431 -1289 -4263 -1255
rect -4053 -1289 -3885 -1255
rect -3675 -1289 -3507 -1255
rect -3297 -1289 -3129 -1255
rect -2919 -1289 -2751 -1255
rect -2541 -1289 -2373 -1255
rect -2163 -1289 -1995 -1255
rect -1785 -1289 -1617 -1255
rect -1407 -1289 -1239 -1255
rect -1029 -1289 -861 -1255
rect -651 -1289 -483 -1255
rect -273 -1289 -105 -1255
rect 105 -1289 273 -1255
rect 483 -1289 651 -1255
rect 861 -1289 1029 -1255
rect 1239 -1289 1407 -1255
rect 1617 -1289 1785 -1255
rect 1995 -1289 2163 -1255
rect 2373 -1289 2541 -1255
rect 2751 -1289 2919 -1255
rect 3129 -1289 3297 -1255
rect 3507 -1289 3675 -1255
rect 3885 -1289 4053 -1255
rect 4263 -1289 4431 -1255
rect 4641 -1289 4809 -1255
rect 5019 -1289 5187 -1255
rect 5397 -1289 5565 -1255
rect 5775 -1289 5943 -1255
rect 6153 -1289 6321 -1255
rect 6531 -1289 6699 -1255
rect 6909 -1289 7077 -1255
rect 7287 -1289 7455 -1255
rect 7665 -1289 7833 -1255
rect 8043 -1289 8211 -1255
rect 8421 -1289 8589 -1255
rect 8799 -1289 8967 -1255
rect 9177 -1289 9345 -1255
rect -9345 -2399 -9177 -2365
rect -8967 -2399 -8799 -2365
rect -8589 -2399 -8421 -2365
rect -8211 -2399 -8043 -2365
rect -7833 -2399 -7665 -2365
rect -7455 -2399 -7287 -2365
rect -7077 -2399 -6909 -2365
rect -6699 -2399 -6531 -2365
rect -6321 -2399 -6153 -2365
rect -5943 -2399 -5775 -2365
rect -5565 -2399 -5397 -2365
rect -5187 -2399 -5019 -2365
rect -4809 -2399 -4641 -2365
rect -4431 -2399 -4263 -2365
rect -4053 -2399 -3885 -2365
rect -3675 -2399 -3507 -2365
rect -3297 -2399 -3129 -2365
rect -2919 -2399 -2751 -2365
rect -2541 -2399 -2373 -2365
rect -2163 -2399 -1995 -2365
rect -1785 -2399 -1617 -2365
rect -1407 -2399 -1239 -2365
rect -1029 -2399 -861 -2365
rect -651 -2399 -483 -2365
rect -273 -2399 -105 -2365
rect 105 -2399 273 -2365
rect 483 -2399 651 -2365
rect 861 -2399 1029 -2365
rect 1239 -2399 1407 -2365
rect 1617 -2399 1785 -2365
rect 1995 -2399 2163 -2365
rect 2373 -2399 2541 -2365
rect 2751 -2399 2919 -2365
rect 3129 -2399 3297 -2365
rect 3507 -2399 3675 -2365
rect 3885 -2399 4053 -2365
rect 4263 -2399 4431 -2365
rect 4641 -2399 4809 -2365
rect 5019 -2399 5187 -2365
rect 5397 -2399 5565 -2365
rect 5775 -2399 5943 -2365
rect 6153 -2399 6321 -2365
rect 6531 -2399 6699 -2365
rect 6909 -2399 7077 -2365
rect 7287 -2399 7455 -2365
rect 7665 -2399 7833 -2365
rect 8043 -2399 8211 -2365
rect 8421 -2399 8589 -2365
rect 8799 -2399 8967 -2365
rect 9177 -2399 9345 -2365
<< locali >>
rect -9541 2503 -9445 2537
rect 9445 2503 9541 2537
rect -9541 2441 -9507 2503
rect 9507 2441 9541 2503
rect -9361 2365 -9345 2399
rect -9177 2365 -9161 2399
rect -8983 2365 -8967 2399
rect -8799 2365 -8783 2399
rect -8605 2365 -8589 2399
rect -8421 2365 -8405 2399
rect -8227 2365 -8211 2399
rect -8043 2365 -8027 2399
rect -7849 2365 -7833 2399
rect -7665 2365 -7649 2399
rect -7471 2365 -7455 2399
rect -7287 2365 -7271 2399
rect -7093 2365 -7077 2399
rect -6909 2365 -6893 2399
rect -6715 2365 -6699 2399
rect -6531 2365 -6515 2399
rect -6337 2365 -6321 2399
rect -6153 2365 -6137 2399
rect -5959 2365 -5943 2399
rect -5775 2365 -5759 2399
rect -5581 2365 -5565 2399
rect -5397 2365 -5381 2399
rect -5203 2365 -5187 2399
rect -5019 2365 -5003 2399
rect -4825 2365 -4809 2399
rect -4641 2365 -4625 2399
rect -4447 2365 -4431 2399
rect -4263 2365 -4247 2399
rect -4069 2365 -4053 2399
rect -3885 2365 -3869 2399
rect -3691 2365 -3675 2399
rect -3507 2365 -3491 2399
rect -3313 2365 -3297 2399
rect -3129 2365 -3113 2399
rect -2935 2365 -2919 2399
rect -2751 2365 -2735 2399
rect -2557 2365 -2541 2399
rect -2373 2365 -2357 2399
rect -2179 2365 -2163 2399
rect -1995 2365 -1979 2399
rect -1801 2365 -1785 2399
rect -1617 2365 -1601 2399
rect -1423 2365 -1407 2399
rect -1239 2365 -1223 2399
rect -1045 2365 -1029 2399
rect -861 2365 -845 2399
rect -667 2365 -651 2399
rect -483 2365 -467 2399
rect -289 2365 -273 2399
rect -105 2365 -89 2399
rect 89 2365 105 2399
rect 273 2365 289 2399
rect 467 2365 483 2399
rect 651 2365 667 2399
rect 845 2365 861 2399
rect 1029 2365 1045 2399
rect 1223 2365 1239 2399
rect 1407 2365 1423 2399
rect 1601 2365 1617 2399
rect 1785 2365 1801 2399
rect 1979 2365 1995 2399
rect 2163 2365 2179 2399
rect 2357 2365 2373 2399
rect 2541 2365 2557 2399
rect 2735 2365 2751 2399
rect 2919 2365 2935 2399
rect 3113 2365 3129 2399
rect 3297 2365 3313 2399
rect 3491 2365 3507 2399
rect 3675 2365 3691 2399
rect 3869 2365 3885 2399
rect 4053 2365 4069 2399
rect 4247 2365 4263 2399
rect 4431 2365 4447 2399
rect 4625 2365 4641 2399
rect 4809 2365 4825 2399
rect 5003 2365 5019 2399
rect 5187 2365 5203 2399
rect 5381 2365 5397 2399
rect 5565 2365 5581 2399
rect 5759 2365 5775 2399
rect 5943 2365 5959 2399
rect 6137 2365 6153 2399
rect 6321 2365 6337 2399
rect 6515 2365 6531 2399
rect 6699 2365 6715 2399
rect 6893 2365 6909 2399
rect 7077 2365 7093 2399
rect 7271 2365 7287 2399
rect 7455 2365 7471 2399
rect 7649 2365 7665 2399
rect 7833 2365 7849 2399
rect 8027 2365 8043 2399
rect 8211 2365 8227 2399
rect 8405 2365 8421 2399
rect 8589 2365 8605 2399
rect 8783 2365 8799 2399
rect 8967 2365 8983 2399
rect 9161 2365 9177 2399
rect 9345 2365 9361 2399
rect -9407 2315 -9373 2331
rect -9407 1323 -9373 1339
rect -9149 2315 -9115 2331
rect -9149 1323 -9115 1339
rect -9029 2315 -8995 2331
rect -9029 1323 -8995 1339
rect -8771 2315 -8737 2331
rect -8771 1323 -8737 1339
rect -8651 2315 -8617 2331
rect -8651 1323 -8617 1339
rect -8393 2315 -8359 2331
rect -8393 1323 -8359 1339
rect -8273 2315 -8239 2331
rect -8273 1323 -8239 1339
rect -8015 2315 -7981 2331
rect -8015 1323 -7981 1339
rect -7895 2315 -7861 2331
rect -7895 1323 -7861 1339
rect -7637 2315 -7603 2331
rect -7637 1323 -7603 1339
rect -7517 2315 -7483 2331
rect -7517 1323 -7483 1339
rect -7259 2315 -7225 2331
rect -7259 1323 -7225 1339
rect -7139 2315 -7105 2331
rect -7139 1323 -7105 1339
rect -6881 2315 -6847 2331
rect -6881 1323 -6847 1339
rect -6761 2315 -6727 2331
rect -6761 1323 -6727 1339
rect -6503 2315 -6469 2331
rect -6503 1323 -6469 1339
rect -6383 2315 -6349 2331
rect -6383 1323 -6349 1339
rect -6125 2315 -6091 2331
rect -6125 1323 -6091 1339
rect -6005 2315 -5971 2331
rect -6005 1323 -5971 1339
rect -5747 2315 -5713 2331
rect -5747 1323 -5713 1339
rect -5627 2315 -5593 2331
rect -5627 1323 -5593 1339
rect -5369 2315 -5335 2331
rect -5369 1323 -5335 1339
rect -5249 2315 -5215 2331
rect -5249 1323 -5215 1339
rect -4991 2315 -4957 2331
rect -4991 1323 -4957 1339
rect -4871 2315 -4837 2331
rect -4871 1323 -4837 1339
rect -4613 2315 -4579 2331
rect -4613 1323 -4579 1339
rect -4493 2315 -4459 2331
rect -4493 1323 -4459 1339
rect -4235 2315 -4201 2331
rect -4235 1323 -4201 1339
rect -4115 2315 -4081 2331
rect -4115 1323 -4081 1339
rect -3857 2315 -3823 2331
rect -3857 1323 -3823 1339
rect -3737 2315 -3703 2331
rect -3737 1323 -3703 1339
rect -3479 2315 -3445 2331
rect -3479 1323 -3445 1339
rect -3359 2315 -3325 2331
rect -3359 1323 -3325 1339
rect -3101 2315 -3067 2331
rect -3101 1323 -3067 1339
rect -2981 2315 -2947 2331
rect -2981 1323 -2947 1339
rect -2723 2315 -2689 2331
rect -2723 1323 -2689 1339
rect -2603 2315 -2569 2331
rect -2603 1323 -2569 1339
rect -2345 2315 -2311 2331
rect -2345 1323 -2311 1339
rect -2225 2315 -2191 2331
rect -2225 1323 -2191 1339
rect -1967 2315 -1933 2331
rect -1967 1323 -1933 1339
rect -1847 2315 -1813 2331
rect -1847 1323 -1813 1339
rect -1589 2315 -1555 2331
rect -1589 1323 -1555 1339
rect -1469 2315 -1435 2331
rect -1469 1323 -1435 1339
rect -1211 2315 -1177 2331
rect -1211 1323 -1177 1339
rect -1091 2315 -1057 2331
rect -1091 1323 -1057 1339
rect -833 2315 -799 2331
rect -833 1323 -799 1339
rect -713 2315 -679 2331
rect -713 1323 -679 1339
rect -455 2315 -421 2331
rect -455 1323 -421 1339
rect -335 2315 -301 2331
rect -335 1323 -301 1339
rect -77 2315 -43 2331
rect -77 1323 -43 1339
rect 43 2315 77 2331
rect 43 1323 77 1339
rect 301 2315 335 2331
rect 301 1323 335 1339
rect 421 2315 455 2331
rect 421 1323 455 1339
rect 679 2315 713 2331
rect 679 1323 713 1339
rect 799 2315 833 2331
rect 799 1323 833 1339
rect 1057 2315 1091 2331
rect 1057 1323 1091 1339
rect 1177 2315 1211 2331
rect 1177 1323 1211 1339
rect 1435 2315 1469 2331
rect 1435 1323 1469 1339
rect 1555 2315 1589 2331
rect 1555 1323 1589 1339
rect 1813 2315 1847 2331
rect 1813 1323 1847 1339
rect 1933 2315 1967 2331
rect 1933 1323 1967 1339
rect 2191 2315 2225 2331
rect 2191 1323 2225 1339
rect 2311 2315 2345 2331
rect 2311 1323 2345 1339
rect 2569 2315 2603 2331
rect 2569 1323 2603 1339
rect 2689 2315 2723 2331
rect 2689 1323 2723 1339
rect 2947 2315 2981 2331
rect 2947 1323 2981 1339
rect 3067 2315 3101 2331
rect 3067 1323 3101 1339
rect 3325 2315 3359 2331
rect 3325 1323 3359 1339
rect 3445 2315 3479 2331
rect 3445 1323 3479 1339
rect 3703 2315 3737 2331
rect 3703 1323 3737 1339
rect 3823 2315 3857 2331
rect 3823 1323 3857 1339
rect 4081 2315 4115 2331
rect 4081 1323 4115 1339
rect 4201 2315 4235 2331
rect 4201 1323 4235 1339
rect 4459 2315 4493 2331
rect 4459 1323 4493 1339
rect 4579 2315 4613 2331
rect 4579 1323 4613 1339
rect 4837 2315 4871 2331
rect 4837 1323 4871 1339
rect 4957 2315 4991 2331
rect 4957 1323 4991 1339
rect 5215 2315 5249 2331
rect 5215 1323 5249 1339
rect 5335 2315 5369 2331
rect 5335 1323 5369 1339
rect 5593 2315 5627 2331
rect 5593 1323 5627 1339
rect 5713 2315 5747 2331
rect 5713 1323 5747 1339
rect 5971 2315 6005 2331
rect 5971 1323 6005 1339
rect 6091 2315 6125 2331
rect 6091 1323 6125 1339
rect 6349 2315 6383 2331
rect 6349 1323 6383 1339
rect 6469 2315 6503 2331
rect 6469 1323 6503 1339
rect 6727 2315 6761 2331
rect 6727 1323 6761 1339
rect 6847 2315 6881 2331
rect 6847 1323 6881 1339
rect 7105 2315 7139 2331
rect 7105 1323 7139 1339
rect 7225 2315 7259 2331
rect 7225 1323 7259 1339
rect 7483 2315 7517 2331
rect 7483 1323 7517 1339
rect 7603 2315 7637 2331
rect 7603 1323 7637 1339
rect 7861 2315 7895 2331
rect 7861 1323 7895 1339
rect 7981 2315 8015 2331
rect 7981 1323 8015 1339
rect 8239 2315 8273 2331
rect 8239 1323 8273 1339
rect 8359 2315 8393 2331
rect 8359 1323 8393 1339
rect 8617 2315 8651 2331
rect 8617 1323 8651 1339
rect 8737 2315 8771 2331
rect 8737 1323 8771 1339
rect 8995 2315 9029 2331
rect 8995 1323 9029 1339
rect 9115 2315 9149 2331
rect 9115 1323 9149 1339
rect 9373 2315 9407 2331
rect 9373 1323 9407 1339
rect -9361 1255 -9345 1289
rect -9177 1255 -9161 1289
rect -8983 1255 -8967 1289
rect -8799 1255 -8783 1289
rect -8605 1255 -8589 1289
rect -8421 1255 -8405 1289
rect -8227 1255 -8211 1289
rect -8043 1255 -8027 1289
rect -7849 1255 -7833 1289
rect -7665 1255 -7649 1289
rect -7471 1255 -7455 1289
rect -7287 1255 -7271 1289
rect -7093 1255 -7077 1289
rect -6909 1255 -6893 1289
rect -6715 1255 -6699 1289
rect -6531 1255 -6515 1289
rect -6337 1255 -6321 1289
rect -6153 1255 -6137 1289
rect -5959 1255 -5943 1289
rect -5775 1255 -5759 1289
rect -5581 1255 -5565 1289
rect -5397 1255 -5381 1289
rect -5203 1255 -5187 1289
rect -5019 1255 -5003 1289
rect -4825 1255 -4809 1289
rect -4641 1255 -4625 1289
rect -4447 1255 -4431 1289
rect -4263 1255 -4247 1289
rect -4069 1255 -4053 1289
rect -3885 1255 -3869 1289
rect -3691 1255 -3675 1289
rect -3507 1255 -3491 1289
rect -3313 1255 -3297 1289
rect -3129 1255 -3113 1289
rect -2935 1255 -2919 1289
rect -2751 1255 -2735 1289
rect -2557 1255 -2541 1289
rect -2373 1255 -2357 1289
rect -2179 1255 -2163 1289
rect -1995 1255 -1979 1289
rect -1801 1255 -1785 1289
rect -1617 1255 -1601 1289
rect -1423 1255 -1407 1289
rect -1239 1255 -1223 1289
rect -1045 1255 -1029 1289
rect -861 1255 -845 1289
rect -667 1255 -651 1289
rect -483 1255 -467 1289
rect -289 1255 -273 1289
rect -105 1255 -89 1289
rect 89 1255 105 1289
rect 273 1255 289 1289
rect 467 1255 483 1289
rect 651 1255 667 1289
rect 845 1255 861 1289
rect 1029 1255 1045 1289
rect 1223 1255 1239 1289
rect 1407 1255 1423 1289
rect 1601 1255 1617 1289
rect 1785 1255 1801 1289
rect 1979 1255 1995 1289
rect 2163 1255 2179 1289
rect 2357 1255 2373 1289
rect 2541 1255 2557 1289
rect 2735 1255 2751 1289
rect 2919 1255 2935 1289
rect 3113 1255 3129 1289
rect 3297 1255 3313 1289
rect 3491 1255 3507 1289
rect 3675 1255 3691 1289
rect 3869 1255 3885 1289
rect 4053 1255 4069 1289
rect 4247 1255 4263 1289
rect 4431 1255 4447 1289
rect 4625 1255 4641 1289
rect 4809 1255 4825 1289
rect 5003 1255 5019 1289
rect 5187 1255 5203 1289
rect 5381 1255 5397 1289
rect 5565 1255 5581 1289
rect 5759 1255 5775 1289
rect 5943 1255 5959 1289
rect 6137 1255 6153 1289
rect 6321 1255 6337 1289
rect 6515 1255 6531 1289
rect 6699 1255 6715 1289
rect 6893 1255 6909 1289
rect 7077 1255 7093 1289
rect 7271 1255 7287 1289
rect 7455 1255 7471 1289
rect 7649 1255 7665 1289
rect 7833 1255 7849 1289
rect 8027 1255 8043 1289
rect 8211 1255 8227 1289
rect 8405 1255 8421 1289
rect 8589 1255 8605 1289
rect 8783 1255 8799 1289
rect 8967 1255 8983 1289
rect 9161 1255 9177 1289
rect 9345 1255 9361 1289
rect -9361 1147 -9345 1181
rect -9177 1147 -9161 1181
rect -8983 1147 -8967 1181
rect -8799 1147 -8783 1181
rect -8605 1147 -8589 1181
rect -8421 1147 -8405 1181
rect -8227 1147 -8211 1181
rect -8043 1147 -8027 1181
rect -7849 1147 -7833 1181
rect -7665 1147 -7649 1181
rect -7471 1147 -7455 1181
rect -7287 1147 -7271 1181
rect -7093 1147 -7077 1181
rect -6909 1147 -6893 1181
rect -6715 1147 -6699 1181
rect -6531 1147 -6515 1181
rect -6337 1147 -6321 1181
rect -6153 1147 -6137 1181
rect -5959 1147 -5943 1181
rect -5775 1147 -5759 1181
rect -5581 1147 -5565 1181
rect -5397 1147 -5381 1181
rect -5203 1147 -5187 1181
rect -5019 1147 -5003 1181
rect -4825 1147 -4809 1181
rect -4641 1147 -4625 1181
rect -4447 1147 -4431 1181
rect -4263 1147 -4247 1181
rect -4069 1147 -4053 1181
rect -3885 1147 -3869 1181
rect -3691 1147 -3675 1181
rect -3507 1147 -3491 1181
rect -3313 1147 -3297 1181
rect -3129 1147 -3113 1181
rect -2935 1147 -2919 1181
rect -2751 1147 -2735 1181
rect -2557 1147 -2541 1181
rect -2373 1147 -2357 1181
rect -2179 1147 -2163 1181
rect -1995 1147 -1979 1181
rect -1801 1147 -1785 1181
rect -1617 1147 -1601 1181
rect -1423 1147 -1407 1181
rect -1239 1147 -1223 1181
rect -1045 1147 -1029 1181
rect -861 1147 -845 1181
rect -667 1147 -651 1181
rect -483 1147 -467 1181
rect -289 1147 -273 1181
rect -105 1147 -89 1181
rect 89 1147 105 1181
rect 273 1147 289 1181
rect 467 1147 483 1181
rect 651 1147 667 1181
rect 845 1147 861 1181
rect 1029 1147 1045 1181
rect 1223 1147 1239 1181
rect 1407 1147 1423 1181
rect 1601 1147 1617 1181
rect 1785 1147 1801 1181
rect 1979 1147 1995 1181
rect 2163 1147 2179 1181
rect 2357 1147 2373 1181
rect 2541 1147 2557 1181
rect 2735 1147 2751 1181
rect 2919 1147 2935 1181
rect 3113 1147 3129 1181
rect 3297 1147 3313 1181
rect 3491 1147 3507 1181
rect 3675 1147 3691 1181
rect 3869 1147 3885 1181
rect 4053 1147 4069 1181
rect 4247 1147 4263 1181
rect 4431 1147 4447 1181
rect 4625 1147 4641 1181
rect 4809 1147 4825 1181
rect 5003 1147 5019 1181
rect 5187 1147 5203 1181
rect 5381 1147 5397 1181
rect 5565 1147 5581 1181
rect 5759 1147 5775 1181
rect 5943 1147 5959 1181
rect 6137 1147 6153 1181
rect 6321 1147 6337 1181
rect 6515 1147 6531 1181
rect 6699 1147 6715 1181
rect 6893 1147 6909 1181
rect 7077 1147 7093 1181
rect 7271 1147 7287 1181
rect 7455 1147 7471 1181
rect 7649 1147 7665 1181
rect 7833 1147 7849 1181
rect 8027 1147 8043 1181
rect 8211 1147 8227 1181
rect 8405 1147 8421 1181
rect 8589 1147 8605 1181
rect 8783 1147 8799 1181
rect 8967 1147 8983 1181
rect 9161 1147 9177 1181
rect 9345 1147 9361 1181
rect -9407 1097 -9373 1113
rect -9407 105 -9373 121
rect -9149 1097 -9115 1113
rect -9149 105 -9115 121
rect -9029 1097 -8995 1113
rect -9029 105 -8995 121
rect -8771 1097 -8737 1113
rect -8771 105 -8737 121
rect -8651 1097 -8617 1113
rect -8651 105 -8617 121
rect -8393 1097 -8359 1113
rect -8393 105 -8359 121
rect -8273 1097 -8239 1113
rect -8273 105 -8239 121
rect -8015 1097 -7981 1113
rect -8015 105 -7981 121
rect -7895 1097 -7861 1113
rect -7895 105 -7861 121
rect -7637 1097 -7603 1113
rect -7637 105 -7603 121
rect -7517 1097 -7483 1113
rect -7517 105 -7483 121
rect -7259 1097 -7225 1113
rect -7259 105 -7225 121
rect -7139 1097 -7105 1113
rect -7139 105 -7105 121
rect -6881 1097 -6847 1113
rect -6881 105 -6847 121
rect -6761 1097 -6727 1113
rect -6761 105 -6727 121
rect -6503 1097 -6469 1113
rect -6503 105 -6469 121
rect -6383 1097 -6349 1113
rect -6383 105 -6349 121
rect -6125 1097 -6091 1113
rect -6125 105 -6091 121
rect -6005 1097 -5971 1113
rect -6005 105 -5971 121
rect -5747 1097 -5713 1113
rect -5747 105 -5713 121
rect -5627 1097 -5593 1113
rect -5627 105 -5593 121
rect -5369 1097 -5335 1113
rect -5369 105 -5335 121
rect -5249 1097 -5215 1113
rect -5249 105 -5215 121
rect -4991 1097 -4957 1113
rect -4991 105 -4957 121
rect -4871 1097 -4837 1113
rect -4871 105 -4837 121
rect -4613 1097 -4579 1113
rect -4613 105 -4579 121
rect -4493 1097 -4459 1113
rect -4493 105 -4459 121
rect -4235 1097 -4201 1113
rect -4235 105 -4201 121
rect -4115 1097 -4081 1113
rect -4115 105 -4081 121
rect -3857 1097 -3823 1113
rect -3857 105 -3823 121
rect -3737 1097 -3703 1113
rect -3737 105 -3703 121
rect -3479 1097 -3445 1113
rect -3479 105 -3445 121
rect -3359 1097 -3325 1113
rect -3359 105 -3325 121
rect -3101 1097 -3067 1113
rect -3101 105 -3067 121
rect -2981 1097 -2947 1113
rect -2981 105 -2947 121
rect -2723 1097 -2689 1113
rect -2723 105 -2689 121
rect -2603 1097 -2569 1113
rect -2603 105 -2569 121
rect -2345 1097 -2311 1113
rect -2345 105 -2311 121
rect -2225 1097 -2191 1113
rect -2225 105 -2191 121
rect -1967 1097 -1933 1113
rect -1967 105 -1933 121
rect -1847 1097 -1813 1113
rect -1847 105 -1813 121
rect -1589 1097 -1555 1113
rect -1589 105 -1555 121
rect -1469 1097 -1435 1113
rect -1469 105 -1435 121
rect -1211 1097 -1177 1113
rect -1211 105 -1177 121
rect -1091 1097 -1057 1113
rect -1091 105 -1057 121
rect -833 1097 -799 1113
rect -833 105 -799 121
rect -713 1097 -679 1113
rect -713 105 -679 121
rect -455 1097 -421 1113
rect -455 105 -421 121
rect -335 1097 -301 1113
rect -335 105 -301 121
rect -77 1097 -43 1113
rect -77 105 -43 121
rect 43 1097 77 1113
rect 43 105 77 121
rect 301 1097 335 1113
rect 301 105 335 121
rect 421 1097 455 1113
rect 421 105 455 121
rect 679 1097 713 1113
rect 679 105 713 121
rect 799 1097 833 1113
rect 799 105 833 121
rect 1057 1097 1091 1113
rect 1057 105 1091 121
rect 1177 1097 1211 1113
rect 1177 105 1211 121
rect 1435 1097 1469 1113
rect 1435 105 1469 121
rect 1555 1097 1589 1113
rect 1555 105 1589 121
rect 1813 1097 1847 1113
rect 1813 105 1847 121
rect 1933 1097 1967 1113
rect 1933 105 1967 121
rect 2191 1097 2225 1113
rect 2191 105 2225 121
rect 2311 1097 2345 1113
rect 2311 105 2345 121
rect 2569 1097 2603 1113
rect 2569 105 2603 121
rect 2689 1097 2723 1113
rect 2689 105 2723 121
rect 2947 1097 2981 1113
rect 2947 105 2981 121
rect 3067 1097 3101 1113
rect 3067 105 3101 121
rect 3325 1097 3359 1113
rect 3325 105 3359 121
rect 3445 1097 3479 1113
rect 3445 105 3479 121
rect 3703 1097 3737 1113
rect 3703 105 3737 121
rect 3823 1097 3857 1113
rect 3823 105 3857 121
rect 4081 1097 4115 1113
rect 4081 105 4115 121
rect 4201 1097 4235 1113
rect 4201 105 4235 121
rect 4459 1097 4493 1113
rect 4459 105 4493 121
rect 4579 1097 4613 1113
rect 4579 105 4613 121
rect 4837 1097 4871 1113
rect 4837 105 4871 121
rect 4957 1097 4991 1113
rect 4957 105 4991 121
rect 5215 1097 5249 1113
rect 5215 105 5249 121
rect 5335 1097 5369 1113
rect 5335 105 5369 121
rect 5593 1097 5627 1113
rect 5593 105 5627 121
rect 5713 1097 5747 1113
rect 5713 105 5747 121
rect 5971 1097 6005 1113
rect 5971 105 6005 121
rect 6091 1097 6125 1113
rect 6091 105 6125 121
rect 6349 1097 6383 1113
rect 6349 105 6383 121
rect 6469 1097 6503 1113
rect 6469 105 6503 121
rect 6727 1097 6761 1113
rect 6727 105 6761 121
rect 6847 1097 6881 1113
rect 6847 105 6881 121
rect 7105 1097 7139 1113
rect 7105 105 7139 121
rect 7225 1097 7259 1113
rect 7225 105 7259 121
rect 7483 1097 7517 1113
rect 7483 105 7517 121
rect 7603 1097 7637 1113
rect 7603 105 7637 121
rect 7861 1097 7895 1113
rect 7861 105 7895 121
rect 7981 1097 8015 1113
rect 7981 105 8015 121
rect 8239 1097 8273 1113
rect 8239 105 8273 121
rect 8359 1097 8393 1113
rect 8359 105 8393 121
rect 8617 1097 8651 1113
rect 8617 105 8651 121
rect 8737 1097 8771 1113
rect 8737 105 8771 121
rect 8995 1097 9029 1113
rect 8995 105 9029 121
rect 9115 1097 9149 1113
rect 9115 105 9149 121
rect 9373 1097 9407 1113
rect 9373 105 9407 121
rect -9361 37 -9345 71
rect -9177 37 -9161 71
rect -8983 37 -8967 71
rect -8799 37 -8783 71
rect -8605 37 -8589 71
rect -8421 37 -8405 71
rect -8227 37 -8211 71
rect -8043 37 -8027 71
rect -7849 37 -7833 71
rect -7665 37 -7649 71
rect -7471 37 -7455 71
rect -7287 37 -7271 71
rect -7093 37 -7077 71
rect -6909 37 -6893 71
rect -6715 37 -6699 71
rect -6531 37 -6515 71
rect -6337 37 -6321 71
rect -6153 37 -6137 71
rect -5959 37 -5943 71
rect -5775 37 -5759 71
rect -5581 37 -5565 71
rect -5397 37 -5381 71
rect -5203 37 -5187 71
rect -5019 37 -5003 71
rect -4825 37 -4809 71
rect -4641 37 -4625 71
rect -4447 37 -4431 71
rect -4263 37 -4247 71
rect -4069 37 -4053 71
rect -3885 37 -3869 71
rect -3691 37 -3675 71
rect -3507 37 -3491 71
rect -3313 37 -3297 71
rect -3129 37 -3113 71
rect -2935 37 -2919 71
rect -2751 37 -2735 71
rect -2557 37 -2541 71
rect -2373 37 -2357 71
rect -2179 37 -2163 71
rect -1995 37 -1979 71
rect -1801 37 -1785 71
rect -1617 37 -1601 71
rect -1423 37 -1407 71
rect -1239 37 -1223 71
rect -1045 37 -1029 71
rect -861 37 -845 71
rect -667 37 -651 71
rect -483 37 -467 71
rect -289 37 -273 71
rect -105 37 -89 71
rect 89 37 105 71
rect 273 37 289 71
rect 467 37 483 71
rect 651 37 667 71
rect 845 37 861 71
rect 1029 37 1045 71
rect 1223 37 1239 71
rect 1407 37 1423 71
rect 1601 37 1617 71
rect 1785 37 1801 71
rect 1979 37 1995 71
rect 2163 37 2179 71
rect 2357 37 2373 71
rect 2541 37 2557 71
rect 2735 37 2751 71
rect 2919 37 2935 71
rect 3113 37 3129 71
rect 3297 37 3313 71
rect 3491 37 3507 71
rect 3675 37 3691 71
rect 3869 37 3885 71
rect 4053 37 4069 71
rect 4247 37 4263 71
rect 4431 37 4447 71
rect 4625 37 4641 71
rect 4809 37 4825 71
rect 5003 37 5019 71
rect 5187 37 5203 71
rect 5381 37 5397 71
rect 5565 37 5581 71
rect 5759 37 5775 71
rect 5943 37 5959 71
rect 6137 37 6153 71
rect 6321 37 6337 71
rect 6515 37 6531 71
rect 6699 37 6715 71
rect 6893 37 6909 71
rect 7077 37 7093 71
rect 7271 37 7287 71
rect 7455 37 7471 71
rect 7649 37 7665 71
rect 7833 37 7849 71
rect 8027 37 8043 71
rect 8211 37 8227 71
rect 8405 37 8421 71
rect 8589 37 8605 71
rect 8783 37 8799 71
rect 8967 37 8983 71
rect 9161 37 9177 71
rect 9345 37 9361 71
rect -9361 -71 -9345 -37
rect -9177 -71 -9161 -37
rect -8983 -71 -8967 -37
rect -8799 -71 -8783 -37
rect -8605 -71 -8589 -37
rect -8421 -71 -8405 -37
rect -8227 -71 -8211 -37
rect -8043 -71 -8027 -37
rect -7849 -71 -7833 -37
rect -7665 -71 -7649 -37
rect -7471 -71 -7455 -37
rect -7287 -71 -7271 -37
rect -7093 -71 -7077 -37
rect -6909 -71 -6893 -37
rect -6715 -71 -6699 -37
rect -6531 -71 -6515 -37
rect -6337 -71 -6321 -37
rect -6153 -71 -6137 -37
rect -5959 -71 -5943 -37
rect -5775 -71 -5759 -37
rect -5581 -71 -5565 -37
rect -5397 -71 -5381 -37
rect -5203 -71 -5187 -37
rect -5019 -71 -5003 -37
rect -4825 -71 -4809 -37
rect -4641 -71 -4625 -37
rect -4447 -71 -4431 -37
rect -4263 -71 -4247 -37
rect -4069 -71 -4053 -37
rect -3885 -71 -3869 -37
rect -3691 -71 -3675 -37
rect -3507 -71 -3491 -37
rect -3313 -71 -3297 -37
rect -3129 -71 -3113 -37
rect -2935 -71 -2919 -37
rect -2751 -71 -2735 -37
rect -2557 -71 -2541 -37
rect -2373 -71 -2357 -37
rect -2179 -71 -2163 -37
rect -1995 -71 -1979 -37
rect -1801 -71 -1785 -37
rect -1617 -71 -1601 -37
rect -1423 -71 -1407 -37
rect -1239 -71 -1223 -37
rect -1045 -71 -1029 -37
rect -861 -71 -845 -37
rect -667 -71 -651 -37
rect -483 -71 -467 -37
rect -289 -71 -273 -37
rect -105 -71 -89 -37
rect 89 -71 105 -37
rect 273 -71 289 -37
rect 467 -71 483 -37
rect 651 -71 667 -37
rect 845 -71 861 -37
rect 1029 -71 1045 -37
rect 1223 -71 1239 -37
rect 1407 -71 1423 -37
rect 1601 -71 1617 -37
rect 1785 -71 1801 -37
rect 1979 -71 1995 -37
rect 2163 -71 2179 -37
rect 2357 -71 2373 -37
rect 2541 -71 2557 -37
rect 2735 -71 2751 -37
rect 2919 -71 2935 -37
rect 3113 -71 3129 -37
rect 3297 -71 3313 -37
rect 3491 -71 3507 -37
rect 3675 -71 3691 -37
rect 3869 -71 3885 -37
rect 4053 -71 4069 -37
rect 4247 -71 4263 -37
rect 4431 -71 4447 -37
rect 4625 -71 4641 -37
rect 4809 -71 4825 -37
rect 5003 -71 5019 -37
rect 5187 -71 5203 -37
rect 5381 -71 5397 -37
rect 5565 -71 5581 -37
rect 5759 -71 5775 -37
rect 5943 -71 5959 -37
rect 6137 -71 6153 -37
rect 6321 -71 6337 -37
rect 6515 -71 6531 -37
rect 6699 -71 6715 -37
rect 6893 -71 6909 -37
rect 7077 -71 7093 -37
rect 7271 -71 7287 -37
rect 7455 -71 7471 -37
rect 7649 -71 7665 -37
rect 7833 -71 7849 -37
rect 8027 -71 8043 -37
rect 8211 -71 8227 -37
rect 8405 -71 8421 -37
rect 8589 -71 8605 -37
rect 8783 -71 8799 -37
rect 8967 -71 8983 -37
rect 9161 -71 9177 -37
rect 9345 -71 9361 -37
rect -9407 -121 -9373 -105
rect -9407 -1113 -9373 -1097
rect -9149 -121 -9115 -105
rect -9149 -1113 -9115 -1097
rect -9029 -121 -8995 -105
rect -9029 -1113 -8995 -1097
rect -8771 -121 -8737 -105
rect -8771 -1113 -8737 -1097
rect -8651 -121 -8617 -105
rect -8651 -1113 -8617 -1097
rect -8393 -121 -8359 -105
rect -8393 -1113 -8359 -1097
rect -8273 -121 -8239 -105
rect -8273 -1113 -8239 -1097
rect -8015 -121 -7981 -105
rect -8015 -1113 -7981 -1097
rect -7895 -121 -7861 -105
rect -7895 -1113 -7861 -1097
rect -7637 -121 -7603 -105
rect -7637 -1113 -7603 -1097
rect -7517 -121 -7483 -105
rect -7517 -1113 -7483 -1097
rect -7259 -121 -7225 -105
rect -7259 -1113 -7225 -1097
rect -7139 -121 -7105 -105
rect -7139 -1113 -7105 -1097
rect -6881 -121 -6847 -105
rect -6881 -1113 -6847 -1097
rect -6761 -121 -6727 -105
rect -6761 -1113 -6727 -1097
rect -6503 -121 -6469 -105
rect -6503 -1113 -6469 -1097
rect -6383 -121 -6349 -105
rect -6383 -1113 -6349 -1097
rect -6125 -121 -6091 -105
rect -6125 -1113 -6091 -1097
rect -6005 -121 -5971 -105
rect -6005 -1113 -5971 -1097
rect -5747 -121 -5713 -105
rect -5747 -1113 -5713 -1097
rect -5627 -121 -5593 -105
rect -5627 -1113 -5593 -1097
rect -5369 -121 -5335 -105
rect -5369 -1113 -5335 -1097
rect -5249 -121 -5215 -105
rect -5249 -1113 -5215 -1097
rect -4991 -121 -4957 -105
rect -4991 -1113 -4957 -1097
rect -4871 -121 -4837 -105
rect -4871 -1113 -4837 -1097
rect -4613 -121 -4579 -105
rect -4613 -1113 -4579 -1097
rect -4493 -121 -4459 -105
rect -4493 -1113 -4459 -1097
rect -4235 -121 -4201 -105
rect -4235 -1113 -4201 -1097
rect -4115 -121 -4081 -105
rect -4115 -1113 -4081 -1097
rect -3857 -121 -3823 -105
rect -3857 -1113 -3823 -1097
rect -3737 -121 -3703 -105
rect -3737 -1113 -3703 -1097
rect -3479 -121 -3445 -105
rect -3479 -1113 -3445 -1097
rect -3359 -121 -3325 -105
rect -3359 -1113 -3325 -1097
rect -3101 -121 -3067 -105
rect -3101 -1113 -3067 -1097
rect -2981 -121 -2947 -105
rect -2981 -1113 -2947 -1097
rect -2723 -121 -2689 -105
rect -2723 -1113 -2689 -1097
rect -2603 -121 -2569 -105
rect -2603 -1113 -2569 -1097
rect -2345 -121 -2311 -105
rect -2345 -1113 -2311 -1097
rect -2225 -121 -2191 -105
rect -2225 -1113 -2191 -1097
rect -1967 -121 -1933 -105
rect -1967 -1113 -1933 -1097
rect -1847 -121 -1813 -105
rect -1847 -1113 -1813 -1097
rect -1589 -121 -1555 -105
rect -1589 -1113 -1555 -1097
rect -1469 -121 -1435 -105
rect -1469 -1113 -1435 -1097
rect -1211 -121 -1177 -105
rect -1211 -1113 -1177 -1097
rect -1091 -121 -1057 -105
rect -1091 -1113 -1057 -1097
rect -833 -121 -799 -105
rect -833 -1113 -799 -1097
rect -713 -121 -679 -105
rect -713 -1113 -679 -1097
rect -455 -121 -421 -105
rect -455 -1113 -421 -1097
rect -335 -121 -301 -105
rect -335 -1113 -301 -1097
rect -77 -121 -43 -105
rect -77 -1113 -43 -1097
rect 43 -121 77 -105
rect 43 -1113 77 -1097
rect 301 -121 335 -105
rect 301 -1113 335 -1097
rect 421 -121 455 -105
rect 421 -1113 455 -1097
rect 679 -121 713 -105
rect 679 -1113 713 -1097
rect 799 -121 833 -105
rect 799 -1113 833 -1097
rect 1057 -121 1091 -105
rect 1057 -1113 1091 -1097
rect 1177 -121 1211 -105
rect 1177 -1113 1211 -1097
rect 1435 -121 1469 -105
rect 1435 -1113 1469 -1097
rect 1555 -121 1589 -105
rect 1555 -1113 1589 -1097
rect 1813 -121 1847 -105
rect 1813 -1113 1847 -1097
rect 1933 -121 1967 -105
rect 1933 -1113 1967 -1097
rect 2191 -121 2225 -105
rect 2191 -1113 2225 -1097
rect 2311 -121 2345 -105
rect 2311 -1113 2345 -1097
rect 2569 -121 2603 -105
rect 2569 -1113 2603 -1097
rect 2689 -121 2723 -105
rect 2689 -1113 2723 -1097
rect 2947 -121 2981 -105
rect 2947 -1113 2981 -1097
rect 3067 -121 3101 -105
rect 3067 -1113 3101 -1097
rect 3325 -121 3359 -105
rect 3325 -1113 3359 -1097
rect 3445 -121 3479 -105
rect 3445 -1113 3479 -1097
rect 3703 -121 3737 -105
rect 3703 -1113 3737 -1097
rect 3823 -121 3857 -105
rect 3823 -1113 3857 -1097
rect 4081 -121 4115 -105
rect 4081 -1113 4115 -1097
rect 4201 -121 4235 -105
rect 4201 -1113 4235 -1097
rect 4459 -121 4493 -105
rect 4459 -1113 4493 -1097
rect 4579 -121 4613 -105
rect 4579 -1113 4613 -1097
rect 4837 -121 4871 -105
rect 4837 -1113 4871 -1097
rect 4957 -121 4991 -105
rect 4957 -1113 4991 -1097
rect 5215 -121 5249 -105
rect 5215 -1113 5249 -1097
rect 5335 -121 5369 -105
rect 5335 -1113 5369 -1097
rect 5593 -121 5627 -105
rect 5593 -1113 5627 -1097
rect 5713 -121 5747 -105
rect 5713 -1113 5747 -1097
rect 5971 -121 6005 -105
rect 5971 -1113 6005 -1097
rect 6091 -121 6125 -105
rect 6091 -1113 6125 -1097
rect 6349 -121 6383 -105
rect 6349 -1113 6383 -1097
rect 6469 -121 6503 -105
rect 6469 -1113 6503 -1097
rect 6727 -121 6761 -105
rect 6727 -1113 6761 -1097
rect 6847 -121 6881 -105
rect 6847 -1113 6881 -1097
rect 7105 -121 7139 -105
rect 7105 -1113 7139 -1097
rect 7225 -121 7259 -105
rect 7225 -1113 7259 -1097
rect 7483 -121 7517 -105
rect 7483 -1113 7517 -1097
rect 7603 -121 7637 -105
rect 7603 -1113 7637 -1097
rect 7861 -121 7895 -105
rect 7861 -1113 7895 -1097
rect 7981 -121 8015 -105
rect 7981 -1113 8015 -1097
rect 8239 -121 8273 -105
rect 8239 -1113 8273 -1097
rect 8359 -121 8393 -105
rect 8359 -1113 8393 -1097
rect 8617 -121 8651 -105
rect 8617 -1113 8651 -1097
rect 8737 -121 8771 -105
rect 8737 -1113 8771 -1097
rect 8995 -121 9029 -105
rect 8995 -1113 9029 -1097
rect 9115 -121 9149 -105
rect 9115 -1113 9149 -1097
rect 9373 -121 9407 -105
rect 9373 -1113 9407 -1097
rect -9361 -1181 -9345 -1147
rect -9177 -1181 -9161 -1147
rect -8983 -1181 -8967 -1147
rect -8799 -1181 -8783 -1147
rect -8605 -1181 -8589 -1147
rect -8421 -1181 -8405 -1147
rect -8227 -1181 -8211 -1147
rect -8043 -1181 -8027 -1147
rect -7849 -1181 -7833 -1147
rect -7665 -1181 -7649 -1147
rect -7471 -1181 -7455 -1147
rect -7287 -1181 -7271 -1147
rect -7093 -1181 -7077 -1147
rect -6909 -1181 -6893 -1147
rect -6715 -1181 -6699 -1147
rect -6531 -1181 -6515 -1147
rect -6337 -1181 -6321 -1147
rect -6153 -1181 -6137 -1147
rect -5959 -1181 -5943 -1147
rect -5775 -1181 -5759 -1147
rect -5581 -1181 -5565 -1147
rect -5397 -1181 -5381 -1147
rect -5203 -1181 -5187 -1147
rect -5019 -1181 -5003 -1147
rect -4825 -1181 -4809 -1147
rect -4641 -1181 -4625 -1147
rect -4447 -1181 -4431 -1147
rect -4263 -1181 -4247 -1147
rect -4069 -1181 -4053 -1147
rect -3885 -1181 -3869 -1147
rect -3691 -1181 -3675 -1147
rect -3507 -1181 -3491 -1147
rect -3313 -1181 -3297 -1147
rect -3129 -1181 -3113 -1147
rect -2935 -1181 -2919 -1147
rect -2751 -1181 -2735 -1147
rect -2557 -1181 -2541 -1147
rect -2373 -1181 -2357 -1147
rect -2179 -1181 -2163 -1147
rect -1995 -1181 -1979 -1147
rect -1801 -1181 -1785 -1147
rect -1617 -1181 -1601 -1147
rect -1423 -1181 -1407 -1147
rect -1239 -1181 -1223 -1147
rect -1045 -1181 -1029 -1147
rect -861 -1181 -845 -1147
rect -667 -1181 -651 -1147
rect -483 -1181 -467 -1147
rect -289 -1181 -273 -1147
rect -105 -1181 -89 -1147
rect 89 -1181 105 -1147
rect 273 -1181 289 -1147
rect 467 -1181 483 -1147
rect 651 -1181 667 -1147
rect 845 -1181 861 -1147
rect 1029 -1181 1045 -1147
rect 1223 -1181 1239 -1147
rect 1407 -1181 1423 -1147
rect 1601 -1181 1617 -1147
rect 1785 -1181 1801 -1147
rect 1979 -1181 1995 -1147
rect 2163 -1181 2179 -1147
rect 2357 -1181 2373 -1147
rect 2541 -1181 2557 -1147
rect 2735 -1181 2751 -1147
rect 2919 -1181 2935 -1147
rect 3113 -1181 3129 -1147
rect 3297 -1181 3313 -1147
rect 3491 -1181 3507 -1147
rect 3675 -1181 3691 -1147
rect 3869 -1181 3885 -1147
rect 4053 -1181 4069 -1147
rect 4247 -1181 4263 -1147
rect 4431 -1181 4447 -1147
rect 4625 -1181 4641 -1147
rect 4809 -1181 4825 -1147
rect 5003 -1181 5019 -1147
rect 5187 -1181 5203 -1147
rect 5381 -1181 5397 -1147
rect 5565 -1181 5581 -1147
rect 5759 -1181 5775 -1147
rect 5943 -1181 5959 -1147
rect 6137 -1181 6153 -1147
rect 6321 -1181 6337 -1147
rect 6515 -1181 6531 -1147
rect 6699 -1181 6715 -1147
rect 6893 -1181 6909 -1147
rect 7077 -1181 7093 -1147
rect 7271 -1181 7287 -1147
rect 7455 -1181 7471 -1147
rect 7649 -1181 7665 -1147
rect 7833 -1181 7849 -1147
rect 8027 -1181 8043 -1147
rect 8211 -1181 8227 -1147
rect 8405 -1181 8421 -1147
rect 8589 -1181 8605 -1147
rect 8783 -1181 8799 -1147
rect 8967 -1181 8983 -1147
rect 9161 -1181 9177 -1147
rect 9345 -1181 9361 -1147
rect -9361 -1289 -9345 -1255
rect -9177 -1289 -9161 -1255
rect -8983 -1289 -8967 -1255
rect -8799 -1289 -8783 -1255
rect -8605 -1289 -8589 -1255
rect -8421 -1289 -8405 -1255
rect -8227 -1289 -8211 -1255
rect -8043 -1289 -8027 -1255
rect -7849 -1289 -7833 -1255
rect -7665 -1289 -7649 -1255
rect -7471 -1289 -7455 -1255
rect -7287 -1289 -7271 -1255
rect -7093 -1289 -7077 -1255
rect -6909 -1289 -6893 -1255
rect -6715 -1289 -6699 -1255
rect -6531 -1289 -6515 -1255
rect -6337 -1289 -6321 -1255
rect -6153 -1289 -6137 -1255
rect -5959 -1289 -5943 -1255
rect -5775 -1289 -5759 -1255
rect -5581 -1289 -5565 -1255
rect -5397 -1289 -5381 -1255
rect -5203 -1289 -5187 -1255
rect -5019 -1289 -5003 -1255
rect -4825 -1289 -4809 -1255
rect -4641 -1289 -4625 -1255
rect -4447 -1289 -4431 -1255
rect -4263 -1289 -4247 -1255
rect -4069 -1289 -4053 -1255
rect -3885 -1289 -3869 -1255
rect -3691 -1289 -3675 -1255
rect -3507 -1289 -3491 -1255
rect -3313 -1289 -3297 -1255
rect -3129 -1289 -3113 -1255
rect -2935 -1289 -2919 -1255
rect -2751 -1289 -2735 -1255
rect -2557 -1289 -2541 -1255
rect -2373 -1289 -2357 -1255
rect -2179 -1289 -2163 -1255
rect -1995 -1289 -1979 -1255
rect -1801 -1289 -1785 -1255
rect -1617 -1289 -1601 -1255
rect -1423 -1289 -1407 -1255
rect -1239 -1289 -1223 -1255
rect -1045 -1289 -1029 -1255
rect -861 -1289 -845 -1255
rect -667 -1289 -651 -1255
rect -483 -1289 -467 -1255
rect -289 -1289 -273 -1255
rect -105 -1289 -89 -1255
rect 89 -1289 105 -1255
rect 273 -1289 289 -1255
rect 467 -1289 483 -1255
rect 651 -1289 667 -1255
rect 845 -1289 861 -1255
rect 1029 -1289 1045 -1255
rect 1223 -1289 1239 -1255
rect 1407 -1289 1423 -1255
rect 1601 -1289 1617 -1255
rect 1785 -1289 1801 -1255
rect 1979 -1289 1995 -1255
rect 2163 -1289 2179 -1255
rect 2357 -1289 2373 -1255
rect 2541 -1289 2557 -1255
rect 2735 -1289 2751 -1255
rect 2919 -1289 2935 -1255
rect 3113 -1289 3129 -1255
rect 3297 -1289 3313 -1255
rect 3491 -1289 3507 -1255
rect 3675 -1289 3691 -1255
rect 3869 -1289 3885 -1255
rect 4053 -1289 4069 -1255
rect 4247 -1289 4263 -1255
rect 4431 -1289 4447 -1255
rect 4625 -1289 4641 -1255
rect 4809 -1289 4825 -1255
rect 5003 -1289 5019 -1255
rect 5187 -1289 5203 -1255
rect 5381 -1289 5397 -1255
rect 5565 -1289 5581 -1255
rect 5759 -1289 5775 -1255
rect 5943 -1289 5959 -1255
rect 6137 -1289 6153 -1255
rect 6321 -1289 6337 -1255
rect 6515 -1289 6531 -1255
rect 6699 -1289 6715 -1255
rect 6893 -1289 6909 -1255
rect 7077 -1289 7093 -1255
rect 7271 -1289 7287 -1255
rect 7455 -1289 7471 -1255
rect 7649 -1289 7665 -1255
rect 7833 -1289 7849 -1255
rect 8027 -1289 8043 -1255
rect 8211 -1289 8227 -1255
rect 8405 -1289 8421 -1255
rect 8589 -1289 8605 -1255
rect 8783 -1289 8799 -1255
rect 8967 -1289 8983 -1255
rect 9161 -1289 9177 -1255
rect 9345 -1289 9361 -1255
rect -9407 -1339 -9373 -1323
rect -9407 -2331 -9373 -2315
rect -9149 -1339 -9115 -1323
rect -9149 -2331 -9115 -2315
rect -9029 -1339 -8995 -1323
rect -9029 -2331 -8995 -2315
rect -8771 -1339 -8737 -1323
rect -8771 -2331 -8737 -2315
rect -8651 -1339 -8617 -1323
rect -8651 -2331 -8617 -2315
rect -8393 -1339 -8359 -1323
rect -8393 -2331 -8359 -2315
rect -8273 -1339 -8239 -1323
rect -8273 -2331 -8239 -2315
rect -8015 -1339 -7981 -1323
rect -8015 -2331 -7981 -2315
rect -7895 -1339 -7861 -1323
rect -7895 -2331 -7861 -2315
rect -7637 -1339 -7603 -1323
rect -7637 -2331 -7603 -2315
rect -7517 -1339 -7483 -1323
rect -7517 -2331 -7483 -2315
rect -7259 -1339 -7225 -1323
rect -7259 -2331 -7225 -2315
rect -7139 -1339 -7105 -1323
rect -7139 -2331 -7105 -2315
rect -6881 -1339 -6847 -1323
rect -6881 -2331 -6847 -2315
rect -6761 -1339 -6727 -1323
rect -6761 -2331 -6727 -2315
rect -6503 -1339 -6469 -1323
rect -6503 -2331 -6469 -2315
rect -6383 -1339 -6349 -1323
rect -6383 -2331 -6349 -2315
rect -6125 -1339 -6091 -1323
rect -6125 -2331 -6091 -2315
rect -6005 -1339 -5971 -1323
rect -6005 -2331 -5971 -2315
rect -5747 -1339 -5713 -1323
rect -5747 -2331 -5713 -2315
rect -5627 -1339 -5593 -1323
rect -5627 -2331 -5593 -2315
rect -5369 -1339 -5335 -1323
rect -5369 -2331 -5335 -2315
rect -5249 -1339 -5215 -1323
rect -5249 -2331 -5215 -2315
rect -4991 -1339 -4957 -1323
rect -4991 -2331 -4957 -2315
rect -4871 -1339 -4837 -1323
rect -4871 -2331 -4837 -2315
rect -4613 -1339 -4579 -1323
rect -4613 -2331 -4579 -2315
rect -4493 -1339 -4459 -1323
rect -4493 -2331 -4459 -2315
rect -4235 -1339 -4201 -1323
rect -4235 -2331 -4201 -2315
rect -4115 -1339 -4081 -1323
rect -4115 -2331 -4081 -2315
rect -3857 -1339 -3823 -1323
rect -3857 -2331 -3823 -2315
rect -3737 -1339 -3703 -1323
rect -3737 -2331 -3703 -2315
rect -3479 -1339 -3445 -1323
rect -3479 -2331 -3445 -2315
rect -3359 -1339 -3325 -1323
rect -3359 -2331 -3325 -2315
rect -3101 -1339 -3067 -1323
rect -3101 -2331 -3067 -2315
rect -2981 -1339 -2947 -1323
rect -2981 -2331 -2947 -2315
rect -2723 -1339 -2689 -1323
rect -2723 -2331 -2689 -2315
rect -2603 -1339 -2569 -1323
rect -2603 -2331 -2569 -2315
rect -2345 -1339 -2311 -1323
rect -2345 -2331 -2311 -2315
rect -2225 -1339 -2191 -1323
rect -2225 -2331 -2191 -2315
rect -1967 -1339 -1933 -1323
rect -1967 -2331 -1933 -2315
rect -1847 -1339 -1813 -1323
rect -1847 -2331 -1813 -2315
rect -1589 -1339 -1555 -1323
rect -1589 -2331 -1555 -2315
rect -1469 -1339 -1435 -1323
rect -1469 -2331 -1435 -2315
rect -1211 -1339 -1177 -1323
rect -1211 -2331 -1177 -2315
rect -1091 -1339 -1057 -1323
rect -1091 -2331 -1057 -2315
rect -833 -1339 -799 -1323
rect -833 -2331 -799 -2315
rect -713 -1339 -679 -1323
rect -713 -2331 -679 -2315
rect -455 -1339 -421 -1323
rect -455 -2331 -421 -2315
rect -335 -1339 -301 -1323
rect -335 -2331 -301 -2315
rect -77 -1339 -43 -1323
rect -77 -2331 -43 -2315
rect 43 -1339 77 -1323
rect 43 -2331 77 -2315
rect 301 -1339 335 -1323
rect 301 -2331 335 -2315
rect 421 -1339 455 -1323
rect 421 -2331 455 -2315
rect 679 -1339 713 -1323
rect 679 -2331 713 -2315
rect 799 -1339 833 -1323
rect 799 -2331 833 -2315
rect 1057 -1339 1091 -1323
rect 1057 -2331 1091 -2315
rect 1177 -1339 1211 -1323
rect 1177 -2331 1211 -2315
rect 1435 -1339 1469 -1323
rect 1435 -2331 1469 -2315
rect 1555 -1339 1589 -1323
rect 1555 -2331 1589 -2315
rect 1813 -1339 1847 -1323
rect 1813 -2331 1847 -2315
rect 1933 -1339 1967 -1323
rect 1933 -2331 1967 -2315
rect 2191 -1339 2225 -1323
rect 2191 -2331 2225 -2315
rect 2311 -1339 2345 -1323
rect 2311 -2331 2345 -2315
rect 2569 -1339 2603 -1323
rect 2569 -2331 2603 -2315
rect 2689 -1339 2723 -1323
rect 2689 -2331 2723 -2315
rect 2947 -1339 2981 -1323
rect 2947 -2331 2981 -2315
rect 3067 -1339 3101 -1323
rect 3067 -2331 3101 -2315
rect 3325 -1339 3359 -1323
rect 3325 -2331 3359 -2315
rect 3445 -1339 3479 -1323
rect 3445 -2331 3479 -2315
rect 3703 -1339 3737 -1323
rect 3703 -2331 3737 -2315
rect 3823 -1339 3857 -1323
rect 3823 -2331 3857 -2315
rect 4081 -1339 4115 -1323
rect 4081 -2331 4115 -2315
rect 4201 -1339 4235 -1323
rect 4201 -2331 4235 -2315
rect 4459 -1339 4493 -1323
rect 4459 -2331 4493 -2315
rect 4579 -1339 4613 -1323
rect 4579 -2331 4613 -2315
rect 4837 -1339 4871 -1323
rect 4837 -2331 4871 -2315
rect 4957 -1339 4991 -1323
rect 4957 -2331 4991 -2315
rect 5215 -1339 5249 -1323
rect 5215 -2331 5249 -2315
rect 5335 -1339 5369 -1323
rect 5335 -2331 5369 -2315
rect 5593 -1339 5627 -1323
rect 5593 -2331 5627 -2315
rect 5713 -1339 5747 -1323
rect 5713 -2331 5747 -2315
rect 5971 -1339 6005 -1323
rect 5971 -2331 6005 -2315
rect 6091 -1339 6125 -1323
rect 6091 -2331 6125 -2315
rect 6349 -1339 6383 -1323
rect 6349 -2331 6383 -2315
rect 6469 -1339 6503 -1323
rect 6469 -2331 6503 -2315
rect 6727 -1339 6761 -1323
rect 6727 -2331 6761 -2315
rect 6847 -1339 6881 -1323
rect 6847 -2331 6881 -2315
rect 7105 -1339 7139 -1323
rect 7105 -2331 7139 -2315
rect 7225 -1339 7259 -1323
rect 7225 -2331 7259 -2315
rect 7483 -1339 7517 -1323
rect 7483 -2331 7517 -2315
rect 7603 -1339 7637 -1323
rect 7603 -2331 7637 -2315
rect 7861 -1339 7895 -1323
rect 7861 -2331 7895 -2315
rect 7981 -1339 8015 -1323
rect 7981 -2331 8015 -2315
rect 8239 -1339 8273 -1323
rect 8239 -2331 8273 -2315
rect 8359 -1339 8393 -1323
rect 8359 -2331 8393 -2315
rect 8617 -1339 8651 -1323
rect 8617 -2331 8651 -2315
rect 8737 -1339 8771 -1323
rect 8737 -2331 8771 -2315
rect 8995 -1339 9029 -1323
rect 8995 -2331 9029 -2315
rect 9115 -1339 9149 -1323
rect 9115 -2331 9149 -2315
rect 9373 -1339 9407 -1323
rect 9373 -2331 9407 -2315
rect -9361 -2399 -9345 -2365
rect -9177 -2399 -9161 -2365
rect -8983 -2399 -8967 -2365
rect -8799 -2399 -8783 -2365
rect -8605 -2399 -8589 -2365
rect -8421 -2399 -8405 -2365
rect -8227 -2399 -8211 -2365
rect -8043 -2399 -8027 -2365
rect -7849 -2399 -7833 -2365
rect -7665 -2399 -7649 -2365
rect -7471 -2399 -7455 -2365
rect -7287 -2399 -7271 -2365
rect -7093 -2399 -7077 -2365
rect -6909 -2399 -6893 -2365
rect -6715 -2399 -6699 -2365
rect -6531 -2399 -6515 -2365
rect -6337 -2399 -6321 -2365
rect -6153 -2399 -6137 -2365
rect -5959 -2399 -5943 -2365
rect -5775 -2399 -5759 -2365
rect -5581 -2399 -5565 -2365
rect -5397 -2399 -5381 -2365
rect -5203 -2399 -5187 -2365
rect -5019 -2399 -5003 -2365
rect -4825 -2399 -4809 -2365
rect -4641 -2399 -4625 -2365
rect -4447 -2399 -4431 -2365
rect -4263 -2399 -4247 -2365
rect -4069 -2399 -4053 -2365
rect -3885 -2399 -3869 -2365
rect -3691 -2399 -3675 -2365
rect -3507 -2399 -3491 -2365
rect -3313 -2399 -3297 -2365
rect -3129 -2399 -3113 -2365
rect -2935 -2399 -2919 -2365
rect -2751 -2399 -2735 -2365
rect -2557 -2399 -2541 -2365
rect -2373 -2399 -2357 -2365
rect -2179 -2399 -2163 -2365
rect -1995 -2399 -1979 -2365
rect -1801 -2399 -1785 -2365
rect -1617 -2399 -1601 -2365
rect -1423 -2399 -1407 -2365
rect -1239 -2399 -1223 -2365
rect -1045 -2399 -1029 -2365
rect -861 -2399 -845 -2365
rect -667 -2399 -651 -2365
rect -483 -2399 -467 -2365
rect -289 -2399 -273 -2365
rect -105 -2399 -89 -2365
rect 89 -2399 105 -2365
rect 273 -2399 289 -2365
rect 467 -2399 483 -2365
rect 651 -2399 667 -2365
rect 845 -2399 861 -2365
rect 1029 -2399 1045 -2365
rect 1223 -2399 1239 -2365
rect 1407 -2399 1423 -2365
rect 1601 -2399 1617 -2365
rect 1785 -2399 1801 -2365
rect 1979 -2399 1995 -2365
rect 2163 -2399 2179 -2365
rect 2357 -2399 2373 -2365
rect 2541 -2399 2557 -2365
rect 2735 -2399 2751 -2365
rect 2919 -2399 2935 -2365
rect 3113 -2399 3129 -2365
rect 3297 -2399 3313 -2365
rect 3491 -2399 3507 -2365
rect 3675 -2399 3691 -2365
rect 3869 -2399 3885 -2365
rect 4053 -2399 4069 -2365
rect 4247 -2399 4263 -2365
rect 4431 -2399 4447 -2365
rect 4625 -2399 4641 -2365
rect 4809 -2399 4825 -2365
rect 5003 -2399 5019 -2365
rect 5187 -2399 5203 -2365
rect 5381 -2399 5397 -2365
rect 5565 -2399 5581 -2365
rect 5759 -2399 5775 -2365
rect 5943 -2399 5959 -2365
rect 6137 -2399 6153 -2365
rect 6321 -2399 6337 -2365
rect 6515 -2399 6531 -2365
rect 6699 -2399 6715 -2365
rect 6893 -2399 6909 -2365
rect 7077 -2399 7093 -2365
rect 7271 -2399 7287 -2365
rect 7455 -2399 7471 -2365
rect 7649 -2399 7665 -2365
rect 7833 -2399 7849 -2365
rect 8027 -2399 8043 -2365
rect 8211 -2399 8227 -2365
rect 8405 -2399 8421 -2365
rect 8589 -2399 8605 -2365
rect 8783 -2399 8799 -2365
rect 8967 -2399 8983 -2365
rect 9161 -2399 9177 -2365
rect 9345 -2399 9361 -2365
rect -9541 -2503 -9507 -2441
rect 9507 -2503 9541 -2441
rect -9541 -2537 -9445 -2503
rect 9445 -2537 9541 -2503
<< viali >>
rect -9345 2365 -9177 2399
rect -8967 2365 -8799 2399
rect -8589 2365 -8421 2399
rect -8211 2365 -8043 2399
rect -7833 2365 -7665 2399
rect -7455 2365 -7287 2399
rect -7077 2365 -6909 2399
rect -6699 2365 -6531 2399
rect -6321 2365 -6153 2399
rect -5943 2365 -5775 2399
rect -5565 2365 -5397 2399
rect -5187 2365 -5019 2399
rect -4809 2365 -4641 2399
rect -4431 2365 -4263 2399
rect -4053 2365 -3885 2399
rect -3675 2365 -3507 2399
rect -3297 2365 -3129 2399
rect -2919 2365 -2751 2399
rect -2541 2365 -2373 2399
rect -2163 2365 -1995 2399
rect -1785 2365 -1617 2399
rect -1407 2365 -1239 2399
rect -1029 2365 -861 2399
rect -651 2365 -483 2399
rect -273 2365 -105 2399
rect 105 2365 273 2399
rect 483 2365 651 2399
rect 861 2365 1029 2399
rect 1239 2365 1407 2399
rect 1617 2365 1785 2399
rect 1995 2365 2163 2399
rect 2373 2365 2541 2399
rect 2751 2365 2919 2399
rect 3129 2365 3297 2399
rect 3507 2365 3675 2399
rect 3885 2365 4053 2399
rect 4263 2365 4431 2399
rect 4641 2365 4809 2399
rect 5019 2365 5187 2399
rect 5397 2365 5565 2399
rect 5775 2365 5943 2399
rect 6153 2365 6321 2399
rect 6531 2365 6699 2399
rect 6909 2365 7077 2399
rect 7287 2365 7455 2399
rect 7665 2365 7833 2399
rect 8043 2365 8211 2399
rect 8421 2365 8589 2399
rect 8799 2365 8967 2399
rect 9177 2365 9345 2399
rect -9407 1339 -9373 2315
rect -9149 1339 -9115 2315
rect -9029 1339 -8995 2315
rect -8771 1339 -8737 2315
rect -8651 1339 -8617 2315
rect -8393 1339 -8359 2315
rect -8273 1339 -8239 2315
rect -8015 1339 -7981 2315
rect -7895 1339 -7861 2315
rect -7637 1339 -7603 2315
rect -7517 1339 -7483 2315
rect -7259 1339 -7225 2315
rect -7139 1339 -7105 2315
rect -6881 1339 -6847 2315
rect -6761 1339 -6727 2315
rect -6503 1339 -6469 2315
rect -6383 1339 -6349 2315
rect -6125 1339 -6091 2315
rect -6005 1339 -5971 2315
rect -5747 1339 -5713 2315
rect -5627 1339 -5593 2315
rect -5369 1339 -5335 2315
rect -5249 1339 -5215 2315
rect -4991 1339 -4957 2315
rect -4871 1339 -4837 2315
rect -4613 1339 -4579 2315
rect -4493 1339 -4459 2315
rect -4235 1339 -4201 2315
rect -4115 1339 -4081 2315
rect -3857 1339 -3823 2315
rect -3737 1339 -3703 2315
rect -3479 1339 -3445 2315
rect -3359 1339 -3325 2315
rect -3101 1339 -3067 2315
rect -2981 1339 -2947 2315
rect -2723 1339 -2689 2315
rect -2603 1339 -2569 2315
rect -2345 1339 -2311 2315
rect -2225 1339 -2191 2315
rect -1967 1339 -1933 2315
rect -1847 1339 -1813 2315
rect -1589 1339 -1555 2315
rect -1469 1339 -1435 2315
rect -1211 1339 -1177 2315
rect -1091 1339 -1057 2315
rect -833 1339 -799 2315
rect -713 1339 -679 2315
rect -455 1339 -421 2315
rect -335 1339 -301 2315
rect -77 1339 -43 2315
rect 43 1339 77 2315
rect 301 1339 335 2315
rect 421 1339 455 2315
rect 679 1339 713 2315
rect 799 1339 833 2315
rect 1057 1339 1091 2315
rect 1177 1339 1211 2315
rect 1435 1339 1469 2315
rect 1555 1339 1589 2315
rect 1813 1339 1847 2315
rect 1933 1339 1967 2315
rect 2191 1339 2225 2315
rect 2311 1339 2345 2315
rect 2569 1339 2603 2315
rect 2689 1339 2723 2315
rect 2947 1339 2981 2315
rect 3067 1339 3101 2315
rect 3325 1339 3359 2315
rect 3445 1339 3479 2315
rect 3703 1339 3737 2315
rect 3823 1339 3857 2315
rect 4081 1339 4115 2315
rect 4201 1339 4235 2315
rect 4459 1339 4493 2315
rect 4579 1339 4613 2315
rect 4837 1339 4871 2315
rect 4957 1339 4991 2315
rect 5215 1339 5249 2315
rect 5335 1339 5369 2315
rect 5593 1339 5627 2315
rect 5713 1339 5747 2315
rect 5971 1339 6005 2315
rect 6091 1339 6125 2315
rect 6349 1339 6383 2315
rect 6469 1339 6503 2315
rect 6727 1339 6761 2315
rect 6847 1339 6881 2315
rect 7105 1339 7139 2315
rect 7225 1339 7259 2315
rect 7483 1339 7517 2315
rect 7603 1339 7637 2315
rect 7861 1339 7895 2315
rect 7981 1339 8015 2315
rect 8239 1339 8273 2315
rect 8359 1339 8393 2315
rect 8617 1339 8651 2315
rect 8737 1339 8771 2315
rect 8995 1339 9029 2315
rect 9115 1339 9149 2315
rect 9373 1339 9407 2315
rect -9345 1255 -9177 1289
rect -8967 1255 -8799 1289
rect -8589 1255 -8421 1289
rect -8211 1255 -8043 1289
rect -7833 1255 -7665 1289
rect -7455 1255 -7287 1289
rect -7077 1255 -6909 1289
rect -6699 1255 -6531 1289
rect -6321 1255 -6153 1289
rect -5943 1255 -5775 1289
rect -5565 1255 -5397 1289
rect -5187 1255 -5019 1289
rect -4809 1255 -4641 1289
rect -4431 1255 -4263 1289
rect -4053 1255 -3885 1289
rect -3675 1255 -3507 1289
rect -3297 1255 -3129 1289
rect -2919 1255 -2751 1289
rect -2541 1255 -2373 1289
rect -2163 1255 -1995 1289
rect -1785 1255 -1617 1289
rect -1407 1255 -1239 1289
rect -1029 1255 -861 1289
rect -651 1255 -483 1289
rect -273 1255 -105 1289
rect 105 1255 273 1289
rect 483 1255 651 1289
rect 861 1255 1029 1289
rect 1239 1255 1407 1289
rect 1617 1255 1785 1289
rect 1995 1255 2163 1289
rect 2373 1255 2541 1289
rect 2751 1255 2919 1289
rect 3129 1255 3297 1289
rect 3507 1255 3675 1289
rect 3885 1255 4053 1289
rect 4263 1255 4431 1289
rect 4641 1255 4809 1289
rect 5019 1255 5187 1289
rect 5397 1255 5565 1289
rect 5775 1255 5943 1289
rect 6153 1255 6321 1289
rect 6531 1255 6699 1289
rect 6909 1255 7077 1289
rect 7287 1255 7455 1289
rect 7665 1255 7833 1289
rect 8043 1255 8211 1289
rect 8421 1255 8589 1289
rect 8799 1255 8967 1289
rect 9177 1255 9345 1289
rect -9345 1147 -9177 1181
rect -8967 1147 -8799 1181
rect -8589 1147 -8421 1181
rect -8211 1147 -8043 1181
rect -7833 1147 -7665 1181
rect -7455 1147 -7287 1181
rect -7077 1147 -6909 1181
rect -6699 1147 -6531 1181
rect -6321 1147 -6153 1181
rect -5943 1147 -5775 1181
rect -5565 1147 -5397 1181
rect -5187 1147 -5019 1181
rect -4809 1147 -4641 1181
rect -4431 1147 -4263 1181
rect -4053 1147 -3885 1181
rect -3675 1147 -3507 1181
rect -3297 1147 -3129 1181
rect -2919 1147 -2751 1181
rect -2541 1147 -2373 1181
rect -2163 1147 -1995 1181
rect -1785 1147 -1617 1181
rect -1407 1147 -1239 1181
rect -1029 1147 -861 1181
rect -651 1147 -483 1181
rect -273 1147 -105 1181
rect 105 1147 273 1181
rect 483 1147 651 1181
rect 861 1147 1029 1181
rect 1239 1147 1407 1181
rect 1617 1147 1785 1181
rect 1995 1147 2163 1181
rect 2373 1147 2541 1181
rect 2751 1147 2919 1181
rect 3129 1147 3297 1181
rect 3507 1147 3675 1181
rect 3885 1147 4053 1181
rect 4263 1147 4431 1181
rect 4641 1147 4809 1181
rect 5019 1147 5187 1181
rect 5397 1147 5565 1181
rect 5775 1147 5943 1181
rect 6153 1147 6321 1181
rect 6531 1147 6699 1181
rect 6909 1147 7077 1181
rect 7287 1147 7455 1181
rect 7665 1147 7833 1181
rect 8043 1147 8211 1181
rect 8421 1147 8589 1181
rect 8799 1147 8967 1181
rect 9177 1147 9345 1181
rect -9407 121 -9373 1097
rect -9149 121 -9115 1097
rect -9029 121 -8995 1097
rect -8771 121 -8737 1097
rect -8651 121 -8617 1097
rect -8393 121 -8359 1097
rect -8273 121 -8239 1097
rect -8015 121 -7981 1097
rect -7895 121 -7861 1097
rect -7637 121 -7603 1097
rect -7517 121 -7483 1097
rect -7259 121 -7225 1097
rect -7139 121 -7105 1097
rect -6881 121 -6847 1097
rect -6761 121 -6727 1097
rect -6503 121 -6469 1097
rect -6383 121 -6349 1097
rect -6125 121 -6091 1097
rect -6005 121 -5971 1097
rect -5747 121 -5713 1097
rect -5627 121 -5593 1097
rect -5369 121 -5335 1097
rect -5249 121 -5215 1097
rect -4991 121 -4957 1097
rect -4871 121 -4837 1097
rect -4613 121 -4579 1097
rect -4493 121 -4459 1097
rect -4235 121 -4201 1097
rect -4115 121 -4081 1097
rect -3857 121 -3823 1097
rect -3737 121 -3703 1097
rect -3479 121 -3445 1097
rect -3359 121 -3325 1097
rect -3101 121 -3067 1097
rect -2981 121 -2947 1097
rect -2723 121 -2689 1097
rect -2603 121 -2569 1097
rect -2345 121 -2311 1097
rect -2225 121 -2191 1097
rect -1967 121 -1933 1097
rect -1847 121 -1813 1097
rect -1589 121 -1555 1097
rect -1469 121 -1435 1097
rect -1211 121 -1177 1097
rect -1091 121 -1057 1097
rect -833 121 -799 1097
rect -713 121 -679 1097
rect -455 121 -421 1097
rect -335 121 -301 1097
rect -77 121 -43 1097
rect 43 121 77 1097
rect 301 121 335 1097
rect 421 121 455 1097
rect 679 121 713 1097
rect 799 121 833 1097
rect 1057 121 1091 1097
rect 1177 121 1211 1097
rect 1435 121 1469 1097
rect 1555 121 1589 1097
rect 1813 121 1847 1097
rect 1933 121 1967 1097
rect 2191 121 2225 1097
rect 2311 121 2345 1097
rect 2569 121 2603 1097
rect 2689 121 2723 1097
rect 2947 121 2981 1097
rect 3067 121 3101 1097
rect 3325 121 3359 1097
rect 3445 121 3479 1097
rect 3703 121 3737 1097
rect 3823 121 3857 1097
rect 4081 121 4115 1097
rect 4201 121 4235 1097
rect 4459 121 4493 1097
rect 4579 121 4613 1097
rect 4837 121 4871 1097
rect 4957 121 4991 1097
rect 5215 121 5249 1097
rect 5335 121 5369 1097
rect 5593 121 5627 1097
rect 5713 121 5747 1097
rect 5971 121 6005 1097
rect 6091 121 6125 1097
rect 6349 121 6383 1097
rect 6469 121 6503 1097
rect 6727 121 6761 1097
rect 6847 121 6881 1097
rect 7105 121 7139 1097
rect 7225 121 7259 1097
rect 7483 121 7517 1097
rect 7603 121 7637 1097
rect 7861 121 7895 1097
rect 7981 121 8015 1097
rect 8239 121 8273 1097
rect 8359 121 8393 1097
rect 8617 121 8651 1097
rect 8737 121 8771 1097
rect 8995 121 9029 1097
rect 9115 121 9149 1097
rect 9373 121 9407 1097
rect -9345 37 -9177 71
rect -8967 37 -8799 71
rect -8589 37 -8421 71
rect -8211 37 -8043 71
rect -7833 37 -7665 71
rect -7455 37 -7287 71
rect -7077 37 -6909 71
rect -6699 37 -6531 71
rect -6321 37 -6153 71
rect -5943 37 -5775 71
rect -5565 37 -5397 71
rect -5187 37 -5019 71
rect -4809 37 -4641 71
rect -4431 37 -4263 71
rect -4053 37 -3885 71
rect -3675 37 -3507 71
rect -3297 37 -3129 71
rect -2919 37 -2751 71
rect -2541 37 -2373 71
rect -2163 37 -1995 71
rect -1785 37 -1617 71
rect -1407 37 -1239 71
rect -1029 37 -861 71
rect -651 37 -483 71
rect -273 37 -105 71
rect 105 37 273 71
rect 483 37 651 71
rect 861 37 1029 71
rect 1239 37 1407 71
rect 1617 37 1785 71
rect 1995 37 2163 71
rect 2373 37 2541 71
rect 2751 37 2919 71
rect 3129 37 3297 71
rect 3507 37 3675 71
rect 3885 37 4053 71
rect 4263 37 4431 71
rect 4641 37 4809 71
rect 5019 37 5187 71
rect 5397 37 5565 71
rect 5775 37 5943 71
rect 6153 37 6321 71
rect 6531 37 6699 71
rect 6909 37 7077 71
rect 7287 37 7455 71
rect 7665 37 7833 71
rect 8043 37 8211 71
rect 8421 37 8589 71
rect 8799 37 8967 71
rect 9177 37 9345 71
rect -9345 -71 -9177 -37
rect -8967 -71 -8799 -37
rect -8589 -71 -8421 -37
rect -8211 -71 -8043 -37
rect -7833 -71 -7665 -37
rect -7455 -71 -7287 -37
rect -7077 -71 -6909 -37
rect -6699 -71 -6531 -37
rect -6321 -71 -6153 -37
rect -5943 -71 -5775 -37
rect -5565 -71 -5397 -37
rect -5187 -71 -5019 -37
rect -4809 -71 -4641 -37
rect -4431 -71 -4263 -37
rect -4053 -71 -3885 -37
rect -3675 -71 -3507 -37
rect -3297 -71 -3129 -37
rect -2919 -71 -2751 -37
rect -2541 -71 -2373 -37
rect -2163 -71 -1995 -37
rect -1785 -71 -1617 -37
rect -1407 -71 -1239 -37
rect -1029 -71 -861 -37
rect -651 -71 -483 -37
rect -273 -71 -105 -37
rect 105 -71 273 -37
rect 483 -71 651 -37
rect 861 -71 1029 -37
rect 1239 -71 1407 -37
rect 1617 -71 1785 -37
rect 1995 -71 2163 -37
rect 2373 -71 2541 -37
rect 2751 -71 2919 -37
rect 3129 -71 3297 -37
rect 3507 -71 3675 -37
rect 3885 -71 4053 -37
rect 4263 -71 4431 -37
rect 4641 -71 4809 -37
rect 5019 -71 5187 -37
rect 5397 -71 5565 -37
rect 5775 -71 5943 -37
rect 6153 -71 6321 -37
rect 6531 -71 6699 -37
rect 6909 -71 7077 -37
rect 7287 -71 7455 -37
rect 7665 -71 7833 -37
rect 8043 -71 8211 -37
rect 8421 -71 8589 -37
rect 8799 -71 8967 -37
rect 9177 -71 9345 -37
rect -9407 -1097 -9373 -121
rect -9149 -1097 -9115 -121
rect -9029 -1097 -8995 -121
rect -8771 -1097 -8737 -121
rect -8651 -1097 -8617 -121
rect -8393 -1097 -8359 -121
rect -8273 -1097 -8239 -121
rect -8015 -1097 -7981 -121
rect -7895 -1097 -7861 -121
rect -7637 -1097 -7603 -121
rect -7517 -1097 -7483 -121
rect -7259 -1097 -7225 -121
rect -7139 -1097 -7105 -121
rect -6881 -1097 -6847 -121
rect -6761 -1097 -6727 -121
rect -6503 -1097 -6469 -121
rect -6383 -1097 -6349 -121
rect -6125 -1097 -6091 -121
rect -6005 -1097 -5971 -121
rect -5747 -1097 -5713 -121
rect -5627 -1097 -5593 -121
rect -5369 -1097 -5335 -121
rect -5249 -1097 -5215 -121
rect -4991 -1097 -4957 -121
rect -4871 -1097 -4837 -121
rect -4613 -1097 -4579 -121
rect -4493 -1097 -4459 -121
rect -4235 -1097 -4201 -121
rect -4115 -1097 -4081 -121
rect -3857 -1097 -3823 -121
rect -3737 -1097 -3703 -121
rect -3479 -1097 -3445 -121
rect -3359 -1097 -3325 -121
rect -3101 -1097 -3067 -121
rect -2981 -1097 -2947 -121
rect -2723 -1097 -2689 -121
rect -2603 -1097 -2569 -121
rect -2345 -1097 -2311 -121
rect -2225 -1097 -2191 -121
rect -1967 -1097 -1933 -121
rect -1847 -1097 -1813 -121
rect -1589 -1097 -1555 -121
rect -1469 -1097 -1435 -121
rect -1211 -1097 -1177 -121
rect -1091 -1097 -1057 -121
rect -833 -1097 -799 -121
rect -713 -1097 -679 -121
rect -455 -1097 -421 -121
rect -335 -1097 -301 -121
rect -77 -1097 -43 -121
rect 43 -1097 77 -121
rect 301 -1097 335 -121
rect 421 -1097 455 -121
rect 679 -1097 713 -121
rect 799 -1097 833 -121
rect 1057 -1097 1091 -121
rect 1177 -1097 1211 -121
rect 1435 -1097 1469 -121
rect 1555 -1097 1589 -121
rect 1813 -1097 1847 -121
rect 1933 -1097 1967 -121
rect 2191 -1097 2225 -121
rect 2311 -1097 2345 -121
rect 2569 -1097 2603 -121
rect 2689 -1097 2723 -121
rect 2947 -1097 2981 -121
rect 3067 -1097 3101 -121
rect 3325 -1097 3359 -121
rect 3445 -1097 3479 -121
rect 3703 -1097 3737 -121
rect 3823 -1097 3857 -121
rect 4081 -1097 4115 -121
rect 4201 -1097 4235 -121
rect 4459 -1097 4493 -121
rect 4579 -1097 4613 -121
rect 4837 -1097 4871 -121
rect 4957 -1097 4991 -121
rect 5215 -1097 5249 -121
rect 5335 -1097 5369 -121
rect 5593 -1097 5627 -121
rect 5713 -1097 5747 -121
rect 5971 -1097 6005 -121
rect 6091 -1097 6125 -121
rect 6349 -1097 6383 -121
rect 6469 -1097 6503 -121
rect 6727 -1097 6761 -121
rect 6847 -1097 6881 -121
rect 7105 -1097 7139 -121
rect 7225 -1097 7259 -121
rect 7483 -1097 7517 -121
rect 7603 -1097 7637 -121
rect 7861 -1097 7895 -121
rect 7981 -1097 8015 -121
rect 8239 -1097 8273 -121
rect 8359 -1097 8393 -121
rect 8617 -1097 8651 -121
rect 8737 -1097 8771 -121
rect 8995 -1097 9029 -121
rect 9115 -1097 9149 -121
rect 9373 -1097 9407 -121
rect -9345 -1181 -9177 -1147
rect -8967 -1181 -8799 -1147
rect -8589 -1181 -8421 -1147
rect -8211 -1181 -8043 -1147
rect -7833 -1181 -7665 -1147
rect -7455 -1181 -7287 -1147
rect -7077 -1181 -6909 -1147
rect -6699 -1181 -6531 -1147
rect -6321 -1181 -6153 -1147
rect -5943 -1181 -5775 -1147
rect -5565 -1181 -5397 -1147
rect -5187 -1181 -5019 -1147
rect -4809 -1181 -4641 -1147
rect -4431 -1181 -4263 -1147
rect -4053 -1181 -3885 -1147
rect -3675 -1181 -3507 -1147
rect -3297 -1181 -3129 -1147
rect -2919 -1181 -2751 -1147
rect -2541 -1181 -2373 -1147
rect -2163 -1181 -1995 -1147
rect -1785 -1181 -1617 -1147
rect -1407 -1181 -1239 -1147
rect -1029 -1181 -861 -1147
rect -651 -1181 -483 -1147
rect -273 -1181 -105 -1147
rect 105 -1181 273 -1147
rect 483 -1181 651 -1147
rect 861 -1181 1029 -1147
rect 1239 -1181 1407 -1147
rect 1617 -1181 1785 -1147
rect 1995 -1181 2163 -1147
rect 2373 -1181 2541 -1147
rect 2751 -1181 2919 -1147
rect 3129 -1181 3297 -1147
rect 3507 -1181 3675 -1147
rect 3885 -1181 4053 -1147
rect 4263 -1181 4431 -1147
rect 4641 -1181 4809 -1147
rect 5019 -1181 5187 -1147
rect 5397 -1181 5565 -1147
rect 5775 -1181 5943 -1147
rect 6153 -1181 6321 -1147
rect 6531 -1181 6699 -1147
rect 6909 -1181 7077 -1147
rect 7287 -1181 7455 -1147
rect 7665 -1181 7833 -1147
rect 8043 -1181 8211 -1147
rect 8421 -1181 8589 -1147
rect 8799 -1181 8967 -1147
rect 9177 -1181 9345 -1147
rect -9345 -1289 -9177 -1255
rect -8967 -1289 -8799 -1255
rect -8589 -1289 -8421 -1255
rect -8211 -1289 -8043 -1255
rect -7833 -1289 -7665 -1255
rect -7455 -1289 -7287 -1255
rect -7077 -1289 -6909 -1255
rect -6699 -1289 -6531 -1255
rect -6321 -1289 -6153 -1255
rect -5943 -1289 -5775 -1255
rect -5565 -1289 -5397 -1255
rect -5187 -1289 -5019 -1255
rect -4809 -1289 -4641 -1255
rect -4431 -1289 -4263 -1255
rect -4053 -1289 -3885 -1255
rect -3675 -1289 -3507 -1255
rect -3297 -1289 -3129 -1255
rect -2919 -1289 -2751 -1255
rect -2541 -1289 -2373 -1255
rect -2163 -1289 -1995 -1255
rect -1785 -1289 -1617 -1255
rect -1407 -1289 -1239 -1255
rect -1029 -1289 -861 -1255
rect -651 -1289 -483 -1255
rect -273 -1289 -105 -1255
rect 105 -1289 273 -1255
rect 483 -1289 651 -1255
rect 861 -1289 1029 -1255
rect 1239 -1289 1407 -1255
rect 1617 -1289 1785 -1255
rect 1995 -1289 2163 -1255
rect 2373 -1289 2541 -1255
rect 2751 -1289 2919 -1255
rect 3129 -1289 3297 -1255
rect 3507 -1289 3675 -1255
rect 3885 -1289 4053 -1255
rect 4263 -1289 4431 -1255
rect 4641 -1289 4809 -1255
rect 5019 -1289 5187 -1255
rect 5397 -1289 5565 -1255
rect 5775 -1289 5943 -1255
rect 6153 -1289 6321 -1255
rect 6531 -1289 6699 -1255
rect 6909 -1289 7077 -1255
rect 7287 -1289 7455 -1255
rect 7665 -1289 7833 -1255
rect 8043 -1289 8211 -1255
rect 8421 -1289 8589 -1255
rect 8799 -1289 8967 -1255
rect 9177 -1289 9345 -1255
rect -9407 -2315 -9373 -1339
rect -9149 -2315 -9115 -1339
rect -9029 -2315 -8995 -1339
rect -8771 -2315 -8737 -1339
rect -8651 -2315 -8617 -1339
rect -8393 -2315 -8359 -1339
rect -8273 -2315 -8239 -1339
rect -8015 -2315 -7981 -1339
rect -7895 -2315 -7861 -1339
rect -7637 -2315 -7603 -1339
rect -7517 -2315 -7483 -1339
rect -7259 -2315 -7225 -1339
rect -7139 -2315 -7105 -1339
rect -6881 -2315 -6847 -1339
rect -6761 -2315 -6727 -1339
rect -6503 -2315 -6469 -1339
rect -6383 -2315 -6349 -1339
rect -6125 -2315 -6091 -1339
rect -6005 -2315 -5971 -1339
rect -5747 -2315 -5713 -1339
rect -5627 -2315 -5593 -1339
rect -5369 -2315 -5335 -1339
rect -5249 -2315 -5215 -1339
rect -4991 -2315 -4957 -1339
rect -4871 -2315 -4837 -1339
rect -4613 -2315 -4579 -1339
rect -4493 -2315 -4459 -1339
rect -4235 -2315 -4201 -1339
rect -4115 -2315 -4081 -1339
rect -3857 -2315 -3823 -1339
rect -3737 -2315 -3703 -1339
rect -3479 -2315 -3445 -1339
rect -3359 -2315 -3325 -1339
rect -3101 -2315 -3067 -1339
rect -2981 -2315 -2947 -1339
rect -2723 -2315 -2689 -1339
rect -2603 -2315 -2569 -1339
rect -2345 -2315 -2311 -1339
rect -2225 -2315 -2191 -1339
rect -1967 -2315 -1933 -1339
rect -1847 -2315 -1813 -1339
rect -1589 -2315 -1555 -1339
rect -1469 -2315 -1435 -1339
rect -1211 -2315 -1177 -1339
rect -1091 -2315 -1057 -1339
rect -833 -2315 -799 -1339
rect -713 -2315 -679 -1339
rect -455 -2315 -421 -1339
rect -335 -2315 -301 -1339
rect -77 -2315 -43 -1339
rect 43 -2315 77 -1339
rect 301 -2315 335 -1339
rect 421 -2315 455 -1339
rect 679 -2315 713 -1339
rect 799 -2315 833 -1339
rect 1057 -2315 1091 -1339
rect 1177 -2315 1211 -1339
rect 1435 -2315 1469 -1339
rect 1555 -2315 1589 -1339
rect 1813 -2315 1847 -1339
rect 1933 -2315 1967 -1339
rect 2191 -2315 2225 -1339
rect 2311 -2315 2345 -1339
rect 2569 -2315 2603 -1339
rect 2689 -2315 2723 -1339
rect 2947 -2315 2981 -1339
rect 3067 -2315 3101 -1339
rect 3325 -2315 3359 -1339
rect 3445 -2315 3479 -1339
rect 3703 -2315 3737 -1339
rect 3823 -2315 3857 -1339
rect 4081 -2315 4115 -1339
rect 4201 -2315 4235 -1339
rect 4459 -2315 4493 -1339
rect 4579 -2315 4613 -1339
rect 4837 -2315 4871 -1339
rect 4957 -2315 4991 -1339
rect 5215 -2315 5249 -1339
rect 5335 -2315 5369 -1339
rect 5593 -2315 5627 -1339
rect 5713 -2315 5747 -1339
rect 5971 -2315 6005 -1339
rect 6091 -2315 6125 -1339
rect 6349 -2315 6383 -1339
rect 6469 -2315 6503 -1339
rect 6727 -2315 6761 -1339
rect 6847 -2315 6881 -1339
rect 7105 -2315 7139 -1339
rect 7225 -2315 7259 -1339
rect 7483 -2315 7517 -1339
rect 7603 -2315 7637 -1339
rect 7861 -2315 7895 -1339
rect 7981 -2315 8015 -1339
rect 8239 -2315 8273 -1339
rect 8359 -2315 8393 -1339
rect 8617 -2315 8651 -1339
rect 8737 -2315 8771 -1339
rect 8995 -2315 9029 -1339
rect 9115 -2315 9149 -1339
rect 9373 -2315 9407 -1339
rect -9345 -2399 -9177 -2365
rect -8967 -2399 -8799 -2365
rect -8589 -2399 -8421 -2365
rect -8211 -2399 -8043 -2365
rect -7833 -2399 -7665 -2365
rect -7455 -2399 -7287 -2365
rect -7077 -2399 -6909 -2365
rect -6699 -2399 -6531 -2365
rect -6321 -2399 -6153 -2365
rect -5943 -2399 -5775 -2365
rect -5565 -2399 -5397 -2365
rect -5187 -2399 -5019 -2365
rect -4809 -2399 -4641 -2365
rect -4431 -2399 -4263 -2365
rect -4053 -2399 -3885 -2365
rect -3675 -2399 -3507 -2365
rect -3297 -2399 -3129 -2365
rect -2919 -2399 -2751 -2365
rect -2541 -2399 -2373 -2365
rect -2163 -2399 -1995 -2365
rect -1785 -2399 -1617 -2365
rect -1407 -2399 -1239 -2365
rect -1029 -2399 -861 -2365
rect -651 -2399 -483 -2365
rect -273 -2399 -105 -2365
rect 105 -2399 273 -2365
rect 483 -2399 651 -2365
rect 861 -2399 1029 -2365
rect 1239 -2399 1407 -2365
rect 1617 -2399 1785 -2365
rect 1995 -2399 2163 -2365
rect 2373 -2399 2541 -2365
rect 2751 -2399 2919 -2365
rect 3129 -2399 3297 -2365
rect 3507 -2399 3675 -2365
rect 3885 -2399 4053 -2365
rect 4263 -2399 4431 -2365
rect 4641 -2399 4809 -2365
rect 5019 -2399 5187 -2365
rect 5397 -2399 5565 -2365
rect 5775 -2399 5943 -2365
rect 6153 -2399 6321 -2365
rect 6531 -2399 6699 -2365
rect 6909 -2399 7077 -2365
rect 7287 -2399 7455 -2365
rect 7665 -2399 7833 -2365
rect 8043 -2399 8211 -2365
rect 8421 -2399 8589 -2365
rect 8799 -2399 8967 -2365
rect 9177 -2399 9345 -2365
<< metal1 >>
rect -9357 2399 -9165 2405
rect -9357 2365 -9345 2399
rect -9177 2365 -9165 2399
rect -9357 2359 -9165 2365
rect -8979 2399 -8787 2405
rect -8979 2365 -8967 2399
rect -8799 2365 -8787 2399
rect -8979 2359 -8787 2365
rect -8601 2399 -8409 2405
rect -8601 2365 -8589 2399
rect -8421 2365 -8409 2399
rect -8601 2359 -8409 2365
rect -8223 2399 -8031 2405
rect -8223 2365 -8211 2399
rect -8043 2365 -8031 2399
rect -8223 2359 -8031 2365
rect -7845 2399 -7653 2405
rect -7845 2365 -7833 2399
rect -7665 2365 -7653 2399
rect -7845 2359 -7653 2365
rect -7467 2399 -7275 2405
rect -7467 2365 -7455 2399
rect -7287 2365 -7275 2399
rect -7467 2359 -7275 2365
rect -7089 2399 -6897 2405
rect -7089 2365 -7077 2399
rect -6909 2365 -6897 2399
rect -7089 2359 -6897 2365
rect -6711 2399 -6519 2405
rect -6711 2365 -6699 2399
rect -6531 2365 -6519 2399
rect -6711 2359 -6519 2365
rect -6333 2399 -6141 2405
rect -6333 2365 -6321 2399
rect -6153 2365 -6141 2399
rect -6333 2359 -6141 2365
rect -5955 2399 -5763 2405
rect -5955 2365 -5943 2399
rect -5775 2365 -5763 2399
rect -5955 2359 -5763 2365
rect -5577 2399 -5385 2405
rect -5577 2365 -5565 2399
rect -5397 2365 -5385 2399
rect -5577 2359 -5385 2365
rect -5199 2399 -5007 2405
rect -5199 2365 -5187 2399
rect -5019 2365 -5007 2399
rect -5199 2359 -5007 2365
rect -4821 2399 -4629 2405
rect -4821 2365 -4809 2399
rect -4641 2365 -4629 2399
rect -4821 2359 -4629 2365
rect -4443 2399 -4251 2405
rect -4443 2365 -4431 2399
rect -4263 2365 -4251 2399
rect -4443 2359 -4251 2365
rect -4065 2399 -3873 2405
rect -4065 2365 -4053 2399
rect -3885 2365 -3873 2399
rect -4065 2359 -3873 2365
rect -3687 2399 -3495 2405
rect -3687 2365 -3675 2399
rect -3507 2365 -3495 2399
rect -3687 2359 -3495 2365
rect -3309 2399 -3117 2405
rect -3309 2365 -3297 2399
rect -3129 2365 -3117 2399
rect -3309 2359 -3117 2365
rect -2931 2399 -2739 2405
rect -2931 2365 -2919 2399
rect -2751 2365 -2739 2399
rect -2931 2359 -2739 2365
rect -2553 2399 -2361 2405
rect -2553 2365 -2541 2399
rect -2373 2365 -2361 2399
rect -2553 2359 -2361 2365
rect -2175 2399 -1983 2405
rect -2175 2365 -2163 2399
rect -1995 2365 -1983 2399
rect -2175 2359 -1983 2365
rect -1797 2399 -1605 2405
rect -1797 2365 -1785 2399
rect -1617 2365 -1605 2399
rect -1797 2359 -1605 2365
rect -1419 2399 -1227 2405
rect -1419 2365 -1407 2399
rect -1239 2365 -1227 2399
rect -1419 2359 -1227 2365
rect -1041 2399 -849 2405
rect -1041 2365 -1029 2399
rect -861 2365 -849 2399
rect -1041 2359 -849 2365
rect -663 2399 -471 2405
rect -663 2365 -651 2399
rect -483 2365 -471 2399
rect -663 2359 -471 2365
rect -285 2399 -93 2405
rect -285 2365 -273 2399
rect -105 2365 -93 2399
rect -285 2359 -93 2365
rect 93 2399 285 2405
rect 93 2365 105 2399
rect 273 2365 285 2399
rect 93 2359 285 2365
rect 471 2399 663 2405
rect 471 2365 483 2399
rect 651 2365 663 2399
rect 471 2359 663 2365
rect 849 2399 1041 2405
rect 849 2365 861 2399
rect 1029 2365 1041 2399
rect 849 2359 1041 2365
rect 1227 2399 1419 2405
rect 1227 2365 1239 2399
rect 1407 2365 1419 2399
rect 1227 2359 1419 2365
rect 1605 2399 1797 2405
rect 1605 2365 1617 2399
rect 1785 2365 1797 2399
rect 1605 2359 1797 2365
rect 1983 2399 2175 2405
rect 1983 2365 1995 2399
rect 2163 2365 2175 2399
rect 1983 2359 2175 2365
rect 2361 2399 2553 2405
rect 2361 2365 2373 2399
rect 2541 2365 2553 2399
rect 2361 2359 2553 2365
rect 2739 2399 2931 2405
rect 2739 2365 2751 2399
rect 2919 2365 2931 2399
rect 2739 2359 2931 2365
rect 3117 2399 3309 2405
rect 3117 2365 3129 2399
rect 3297 2365 3309 2399
rect 3117 2359 3309 2365
rect 3495 2399 3687 2405
rect 3495 2365 3507 2399
rect 3675 2365 3687 2399
rect 3495 2359 3687 2365
rect 3873 2399 4065 2405
rect 3873 2365 3885 2399
rect 4053 2365 4065 2399
rect 3873 2359 4065 2365
rect 4251 2399 4443 2405
rect 4251 2365 4263 2399
rect 4431 2365 4443 2399
rect 4251 2359 4443 2365
rect 4629 2399 4821 2405
rect 4629 2365 4641 2399
rect 4809 2365 4821 2399
rect 4629 2359 4821 2365
rect 5007 2399 5199 2405
rect 5007 2365 5019 2399
rect 5187 2365 5199 2399
rect 5007 2359 5199 2365
rect 5385 2399 5577 2405
rect 5385 2365 5397 2399
rect 5565 2365 5577 2399
rect 5385 2359 5577 2365
rect 5763 2399 5955 2405
rect 5763 2365 5775 2399
rect 5943 2365 5955 2399
rect 5763 2359 5955 2365
rect 6141 2399 6333 2405
rect 6141 2365 6153 2399
rect 6321 2365 6333 2399
rect 6141 2359 6333 2365
rect 6519 2399 6711 2405
rect 6519 2365 6531 2399
rect 6699 2365 6711 2399
rect 6519 2359 6711 2365
rect 6897 2399 7089 2405
rect 6897 2365 6909 2399
rect 7077 2365 7089 2399
rect 6897 2359 7089 2365
rect 7275 2399 7467 2405
rect 7275 2365 7287 2399
rect 7455 2365 7467 2399
rect 7275 2359 7467 2365
rect 7653 2399 7845 2405
rect 7653 2365 7665 2399
rect 7833 2365 7845 2399
rect 7653 2359 7845 2365
rect 8031 2399 8223 2405
rect 8031 2365 8043 2399
rect 8211 2365 8223 2399
rect 8031 2359 8223 2365
rect 8409 2399 8601 2405
rect 8409 2365 8421 2399
rect 8589 2365 8601 2399
rect 8409 2359 8601 2365
rect 8787 2399 8979 2405
rect 8787 2365 8799 2399
rect 8967 2365 8979 2399
rect 8787 2359 8979 2365
rect 9165 2399 9357 2405
rect 9165 2365 9177 2399
rect 9345 2365 9357 2399
rect 9165 2359 9357 2365
rect -9413 2315 -9367 2327
rect -9413 1339 -9407 2315
rect -9373 1339 -9367 2315
rect -9413 1327 -9367 1339
rect -9155 2315 -9109 2327
rect -9155 1339 -9149 2315
rect -9115 1339 -9109 2315
rect -9155 1327 -9109 1339
rect -9035 2315 -8989 2327
rect -9035 1339 -9029 2315
rect -8995 1339 -8989 2315
rect -9035 1327 -8989 1339
rect -8777 2315 -8731 2327
rect -8777 1339 -8771 2315
rect -8737 1339 -8731 2315
rect -8777 1327 -8731 1339
rect -8657 2315 -8611 2327
rect -8657 1339 -8651 2315
rect -8617 1339 -8611 2315
rect -8657 1327 -8611 1339
rect -8399 2315 -8353 2327
rect -8399 1339 -8393 2315
rect -8359 1339 -8353 2315
rect -8399 1327 -8353 1339
rect -8279 2315 -8233 2327
rect -8279 1339 -8273 2315
rect -8239 1339 -8233 2315
rect -8279 1327 -8233 1339
rect -8021 2315 -7975 2327
rect -8021 1339 -8015 2315
rect -7981 1339 -7975 2315
rect -8021 1327 -7975 1339
rect -7901 2315 -7855 2327
rect -7901 1339 -7895 2315
rect -7861 1339 -7855 2315
rect -7901 1327 -7855 1339
rect -7643 2315 -7597 2327
rect -7643 1339 -7637 2315
rect -7603 1339 -7597 2315
rect -7643 1327 -7597 1339
rect -7523 2315 -7477 2327
rect -7523 1339 -7517 2315
rect -7483 1339 -7477 2315
rect -7523 1327 -7477 1339
rect -7265 2315 -7219 2327
rect -7265 1339 -7259 2315
rect -7225 1339 -7219 2315
rect -7265 1327 -7219 1339
rect -7145 2315 -7099 2327
rect -7145 1339 -7139 2315
rect -7105 1339 -7099 2315
rect -7145 1327 -7099 1339
rect -6887 2315 -6841 2327
rect -6887 1339 -6881 2315
rect -6847 1339 -6841 2315
rect -6887 1327 -6841 1339
rect -6767 2315 -6721 2327
rect -6767 1339 -6761 2315
rect -6727 1339 -6721 2315
rect -6767 1327 -6721 1339
rect -6509 2315 -6463 2327
rect -6509 1339 -6503 2315
rect -6469 1339 -6463 2315
rect -6509 1327 -6463 1339
rect -6389 2315 -6343 2327
rect -6389 1339 -6383 2315
rect -6349 1339 -6343 2315
rect -6389 1327 -6343 1339
rect -6131 2315 -6085 2327
rect -6131 1339 -6125 2315
rect -6091 1339 -6085 2315
rect -6131 1327 -6085 1339
rect -6011 2315 -5965 2327
rect -6011 1339 -6005 2315
rect -5971 1339 -5965 2315
rect -6011 1327 -5965 1339
rect -5753 2315 -5707 2327
rect -5753 1339 -5747 2315
rect -5713 1339 -5707 2315
rect -5753 1327 -5707 1339
rect -5633 2315 -5587 2327
rect -5633 1339 -5627 2315
rect -5593 1339 -5587 2315
rect -5633 1327 -5587 1339
rect -5375 2315 -5329 2327
rect -5375 1339 -5369 2315
rect -5335 1339 -5329 2315
rect -5375 1327 -5329 1339
rect -5255 2315 -5209 2327
rect -5255 1339 -5249 2315
rect -5215 1339 -5209 2315
rect -5255 1327 -5209 1339
rect -4997 2315 -4951 2327
rect -4997 1339 -4991 2315
rect -4957 1339 -4951 2315
rect -4997 1327 -4951 1339
rect -4877 2315 -4831 2327
rect -4877 1339 -4871 2315
rect -4837 1339 -4831 2315
rect -4877 1327 -4831 1339
rect -4619 2315 -4573 2327
rect -4619 1339 -4613 2315
rect -4579 1339 -4573 2315
rect -4619 1327 -4573 1339
rect -4499 2315 -4453 2327
rect -4499 1339 -4493 2315
rect -4459 1339 -4453 2315
rect -4499 1327 -4453 1339
rect -4241 2315 -4195 2327
rect -4241 1339 -4235 2315
rect -4201 1339 -4195 2315
rect -4241 1327 -4195 1339
rect -4121 2315 -4075 2327
rect -4121 1339 -4115 2315
rect -4081 1339 -4075 2315
rect -4121 1327 -4075 1339
rect -3863 2315 -3817 2327
rect -3863 1339 -3857 2315
rect -3823 1339 -3817 2315
rect -3863 1327 -3817 1339
rect -3743 2315 -3697 2327
rect -3743 1339 -3737 2315
rect -3703 1339 -3697 2315
rect -3743 1327 -3697 1339
rect -3485 2315 -3439 2327
rect -3485 1339 -3479 2315
rect -3445 1339 -3439 2315
rect -3485 1327 -3439 1339
rect -3365 2315 -3319 2327
rect -3365 1339 -3359 2315
rect -3325 1339 -3319 2315
rect -3365 1327 -3319 1339
rect -3107 2315 -3061 2327
rect -3107 1339 -3101 2315
rect -3067 1339 -3061 2315
rect -3107 1327 -3061 1339
rect -2987 2315 -2941 2327
rect -2987 1339 -2981 2315
rect -2947 1339 -2941 2315
rect -2987 1327 -2941 1339
rect -2729 2315 -2683 2327
rect -2729 1339 -2723 2315
rect -2689 1339 -2683 2315
rect -2729 1327 -2683 1339
rect -2609 2315 -2563 2327
rect -2609 1339 -2603 2315
rect -2569 1339 -2563 2315
rect -2609 1327 -2563 1339
rect -2351 2315 -2305 2327
rect -2351 1339 -2345 2315
rect -2311 1339 -2305 2315
rect -2351 1327 -2305 1339
rect -2231 2315 -2185 2327
rect -2231 1339 -2225 2315
rect -2191 1339 -2185 2315
rect -2231 1327 -2185 1339
rect -1973 2315 -1927 2327
rect -1973 1339 -1967 2315
rect -1933 1339 -1927 2315
rect -1973 1327 -1927 1339
rect -1853 2315 -1807 2327
rect -1853 1339 -1847 2315
rect -1813 1339 -1807 2315
rect -1853 1327 -1807 1339
rect -1595 2315 -1549 2327
rect -1595 1339 -1589 2315
rect -1555 1339 -1549 2315
rect -1595 1327 -1549 1339
rect -1475 2315 -1429 2327
rect -1475 1339 -1469 2315
rect -1435 1339 -1429 2315
rect -1475 1327 -1429 1339
rect -1217 2315 -1171 2327
rect -1217 1339 -1211 2315
rect -1177 1339 -1171 2315
rect -1217 1327 -1171 1339
rect -1097 2315 -1051 2327
rect -1097 1339 -1091 2315
rect -1057 1339 -1051 2315
rect -1097 1327 -1051 1339
rect -839 2315 -793 2327
rect -839 1339 -833 2315
rect -799 1339 -793 2315
rect -839 1327 -793 1339
rect -719 2315 -673 2327
rect -719 1339 -713 2315
rect -679 1339 -673 2315
rect -719 1327 -673 1339
rect -461 2315 -415 2327
rect -461 1339 -455 2315
rect -421 1339 -415 2315
rect -461 1327 -415 1339
rect -341 2315 -295 2327
rect -341 1339 -335 2315
rect -301 1339 -295 2315
rect -341 1327 -295 1339
rect -83 2315 -37 2327
rect -83 1339 -77 2315
rect -43 1339 -37 2315
rect -83 1327 -37 1339
rect 37 2315 83 2327
rect 37 1339 43 2315
rect 77 1339 83 2315
rect 37 1327 83 1339
rect 295 2315 341 2327
rect 295 1339 301 2315
rect 335 1339 341 2315
rect 295 1327 341 1339
rect 415 2315 461 2327
rect 415 1339 421 2315
rect 455 1339 461 2315
rect 415 1327 461 1339
rect 673 2315 719 2327
rect 673 1339 679 2315
rect 713 1339 719 2315
rect 673 1327 719 1339
rect 793 2315 839 2327
rect 793 1339 799 2315
rect 833 1339 839 2315
rect 793 1327 839 1339
rect 1051 2315 1097 2327
rect 1051 1339 1057 2315
rect 1091 1339 1097 2315
rect 1051 1327 1097 1339
rect 1171 2315 1217 2327
rect 1171 1339 1177 2315
rect 1211 1339 1217 2315
rect 1171 1327 1217 1339
rect 1429 2315 1475 2327
rect 1429 1339 1435 2315
rect 1469 1339 1475 2315
rect 1429 1327 1475 1339
rect 1549 2315 1595 2327
rect 1549 1339 1555 2315
rect 1589 1339 1595 2315
rect 1549 1327 1595 1339
rect 1807 2315 1853 2327
rect 1807 1339 1813 2315
rect 1847 1339 1853 2315
rect 1807 1327 1853 1339
rect 1927 2315 1973 2327
rect 1927 1339 1933 2315
rect 1967 1339 1973 2315
rect 1927 1327 1973 1339
rect 2185 2315 2231 2327
rect 2185 1339 2191 2315
rect 2225 1339 2231 2315
rect 2185 1327 2231 1339
rect 2305 2315 2351 2327
rect 2305 1339 2311 2315
rect 2345 1339 2351 2315
rect 2305 1327 2351 1339
rect 2563 2315 2609 2327
rect 2563 1339 2569 2315
rect 2603 1339 2609 2315
rect 2563 1327 2609 1339
rect 2683 2315 2729 2327
rect 2683 1339 2689 2315
rect 2723 1339 2729 2315
rect 2683 1327 2729 1339
rect 2941 2315 2987 2327
rect 2941 1339 2947 2315
rect 2981 1339 2987 2315
rect 2941 1327 2987 1339
rect 3061 2315 3107 2327
rect 3061 1339 3067 2315
rect 3101 1339 3107 2315
rect 3061 1327 3107 1339
rect 3319 2315 3365 2327
rect 3319 1339 3325 2315
rect 3359 1339 3365 2315
rect 3319 1327 3365 1339
rect 3439 2315 3485 2327
rect 3439 1339 3445 2315
rect 3479 1339 3485 2315
rect 3439 1327 3485 1339
rect 3697 2315 3743 2327
rect 3697 1339 3703 2315
rect 3737 1339 3743 2315
rect 3697 1327 3743 1339
rect 3817 2315 3863 2327
rect 3817 1339 3823 2315
rect 3857 1339 3863 2315
rect 3817 1327 3863 1339
rect 4075 2315 4121 2327
rect 4075 1339 4081 2315
rect 4115 1339 4121 2315
rect 4075 1327 4121 1339
rect 4195 2315 4241 2327
rect 4195 1339 4201 2315
rect 4235 1339 4241 2315
rect 4195 1327 4241 1339
rect 4453 2315 4499 2327
rect 4453 1339 4459 2315
rect 4493 1339 4499 2315
rect 4453 1327 4499 1339
rect 4573 2315 4619 2327
rect 4573 1339 4579 2315
rect 4613 1339 4619 2315
rect 4573 1327 4619 1339
rect 4831 2315 4877 2327
rect 4831 1339 4837 2315
rect 4871 1339 4877 2315
rect 4831 1327 4877 1339
rect 4951 2315 4997 2327
rect 4951 1339 4957 2315
rect 4991 1339 4997 2315
rect 4951 1327 4997 1339
rect 5209 2315 5255 2327
rect 5209 1339 5215 2315
rect 5249 1339 5255 2315
rect 5209 1327 5255 1339
rect 5329 2315 5375 2327
rect 5329 1339 5335 2315
rect 5369 1339 5375 2315
rect 5329 1327 5375 1339
rect 5587 2315 5633 2327
rect 5587 1339 5593 2315
rect 5627 1339 5633 2315
rect 5587 1327 5633 1339
rect 5707 2315 5753 2327
rect 5707 1339 5713 2315
rect 5747 1339 5753 2315
rect 5707 1327 5753 1339
rect 5965 2315 6011 2327
rect 5965 1339 5971 2315
rect 6005 1339 6011 2315
rect 5965 1327 6011 1339
rect 6085 2315 6131 2327
rect 6085 1339 6091 2315
rect 6125 1339 6131 2315
rect 6085 1327 6131 1339
rect 6343 2315 6389 2327
rect 6343 1339 6349 2315
rect 6383 1339 6389 2315
rect 6343 1327 6389 1339
rect 6463 2315 6509 2327
rect 6463 1339 6469 2315
rect 6503 1339 6509 2315
rect 6463 1327 6509 1339
rect 6721 2315 6767 2327
rect 6721 1339 6727 2315
rect 6761 1339 6767 2315
rect 6721 1327 6767 1339
rect 6841 2315 6887 2327
rect 6841 1339 6847 2315
rect 6881 1339 6887 2315
rect 6841 1327 6887 1339
rect 7099 2315 7145 2327
rect 7099 1339 7105 2315
rect 7139 1339 7145 2315
rect 7099 1327 7145 1339
rect 7219 2315 7265 2327
rect 7219 1339 7225 2315
rect 7259 1339 7265 2315
rect 7219 1327 7265 1339
rect 7477 2315 7523 2327
rect 7477 1339 7483 2315
rect 7517 1339 7523 2315
rect 7477 1327 7523 1339
rect 7597 2315 7643 2327
rect 7597 1339 7603 2315
rect 7637 1339 7643 2315
rect 7597 1327 7643 1339
rect 7855 2315 7901 2327
rect 7855 1339 7861 2315
rect 7895 1339 7901 2315
rect 7855 1327 7901 1339
rect 7975 2315 8021 2327
rect 7975 1339 7981 2315
rect 8015 1339 8021 2315
rect 7975 1327 8021 1339
rect 8233 2315 8279 2327
rect 8233 1339 8239 2315
rect 8273 1339 8279 2315
rect 8233 1327 8279 1339
rect 8353 2315 8399 2327
rect 8353 1339 8359 2315
rect 8393 1339 8399 2315
rect 8353 1327 8399 1339
rect 8611 2315 8657 2327
rect 8611 1339 8617 2315
rect 8651 1339 8657 2315
rect 8611 1327 8657 1339
rect 8731 2315 8777 2327
rect 8731 1339 8737 2315
rect 8771 1339 8777 2315
rect 8731 1327 8777 1339
rect 8989 2315 9035 2327
rect 8989 1339 8995 2315
rect 9029 1339 9035 2315
rect 8989 1327 9035 1339
rect 9109 2315 9155 2327
rect 9109 1339 9115 2315
rect 9149 1339 9155 2315
rect 9109 1327 9155 1339
rect 9367 2315 9413 2327
rect 9367 1339 9373 2315
rect 9407 1339 9413 2315
rect 9367 1327 9413 1339
rect -9357 1289 -9165 1295
rect -9357 1255 -9345 1289
rect -9177 1255 -9165 1289
rect -9357 1249 -9165 1255
rect -8979 1289 -8787 1295
rect -8979 1255 -8967 1289
rect -8799 1255 -8787 1289
rect -8979 1249 -8787 1255
rect -8601 1289 -8409 1295
rect -8601 1255 -8589 1289
rect -8421 1255 -8409 1289
rect -8601 1249 -8409 1255
rect -8223 1289 -8031 1295
rect -8223 1255 -8211 1289
rect -8043 1255 -8031 1289
rect -8223 1249 -8031 1255
rect -7845 1289 -7653 1295
rect -7845 1255 -7833 1289
rect -7665 1255 -7653 1289
rect -7845 1249 -7653 1255
rect -7467 1289 -7275 1295
rect -7467 1255 -7455 1289
rect -7287 1255 -7275 1289
rect -7467 1249 -7275 1255
rect -7089 1289 -6897 1295
rect -7089 1255 -7077 1289
rect -6909 1255 -6897 1289
rect -7089 1249 -6897 1255
rect -6711 1289 -6519 1295
rect -6711 1255 -6699 1289
rect -6531 1255 -6519 1289
rect -6711 1249 -6519 1255
rect -6333 1289 -6141 1295
rect -6333 1255 -6321 1289
rect -6153 1255 -6141 1289
rect -6333 1249 -6141 1255
rect -5955 1289 -5763 1295
rect -5955 1255 -5943 1289
rect -5775 1255 -5763 1289
rect -5955 1249 -5763 1255
rect -5577 1289 -5385 1295
rect -5577 1255 -5565 1289
rect -5397 1255 -5385 1289
rect -5577 1249 -5385 1255
rect -5199 1289 -5007 1295
rect -5199 1255 -5187 1289
rect -5019 1255 -5007 1289
rect -5199 1249 -5007 1255
rect -4821 1289 -4629 1295
rect -4821 1255 -4809 1289
rect -4641 1255 -4629 1289
rect -4821 1249 -4629 1255
rect -4443 1289 -4251 1295
rect -4443 1255 -4431 1289
rect -4263 1255 -4251 1289
rect -4443 1249 -4251 1255
rect -4065 1289 -3873 1295
rect -4065 1255 -4053 1289
rect -3885 1255 -3873 1289
rect -4065 1249 -3873 1255
rect -3687 1289 -3495 1295
rect -3687 1255 -3675 1289
rect -3507 1255 -3495 1289
rect -3687 1249 -3495 1255
rect -3309 1289 -3117 1295
rect -3309 1255 -3297 1289
rect -3129 1255 -3117 1289
rect -3309 1249 -3117 1255
rect -2931 1289 -2739 1295
rect -2931 1255 -2919 1289
rect -2751 1255 -2739 1289
rect -2931 1249 -2739 1255
rect -2553 1289 -2361 1295
rect -2553 1255 -2541 1289
rect -2373 1255 -2361 1289
rect -2553 1249 -2361 1255
rect -2175 1289 -1983 1295
rect -2175 1255 -2163 1289
rect -1995 1255 -1983 1289
rect -2175 1249 -1983 1255
rect -1797 1289 -1605 1295
rect -1797 1255 -1785 1289
rect -1617 1255 -1605 1289
rect -1797 1249 -1605 1255
rect -1419 1289 -1227 1295
rect -1419 1255 -1407 1289
rect -1239 1255 -1227 1289
rect -1419 1249 -1227 1255
rect -1041 1289 -849 1295
rect -1041 1255 -1029 1289
rect -861 1255 -849 1289
rect -1041 1249 -849 1255
rect -663 1289 -471 1295
rect -663 1255 -651 1289
rect -483 1255 -471 1289
rect -663 1249 -471 1255
rect -285 1289 -93 1295
rect -285 1255 -273 1289
rect -105 1255 -93 1289
rect -285 1249 -93 1255
rect 93 1289 285 1295
rect 93 1255 105 1289
rect 273 1255 285 1289
rect 93 1249 285 1255
rect 471 1289 663 1295
rect 471 1255 483 1289
rect 651 1255 663 1289
rect 471 1249 663 1255
rect 849 1289 1041 1295
rect 849 1255 861 1289
rect 1029 1255 1041 1289
rect 849 1249 1041 1255
rect 1227 1289 1419 1295
rect 1227 1255 1239 1289
rect 1407 1255 1419 1289
rect 1227 1249 1419 1255
rect 1605 1289 1797 1295
rect 1605 1255 1617 1289
rect 1785 1255 1797 1289
rect 1605 1249 1797 1255
rect 1983 1289 2175 1295
rect 1983 1255 1995 1289
rect 2163 1255 2175 1289
rect 1983 1249 2175 1255
rect 2361 1289 2553 1295
rect 2361 1255 2373 1289
rect 2541 1255 2553 1289
rect 2361 1249 2553 1255
rect 2739 1289 2931 1295
rect 2739 1255 2751 1289
rect 2919 1255 2931 1289
rect 2739 1249 2931 1255
rect 3117 1289 3309 1295
rect 3117 1255 3129 1289
rect 3297 1255 3309 1289
rect 3117 1249 3309 1255
rect 3495 1289 3687 1295
rect 3495 1255 3507 1289
rect 3675 1255 3687 1289
rect 3495 1249 3687 1255
rect 3873 1289 4065 1295
rect 3873 1255 3885 1289
rect 4053 1255 4065 1289
rect 3873 1249 4065 1255
rect 4251 1289 4443 1295
rect 4251 1255 4263 1289
rect 4431 1255 4443 1289
rect 4251 1249 4443 1255
rect 4629 1289 4821 1295
rect 4629 1255 4641 1289
rect 4809 1255 4821 1289
rect 4629 1249 4821 1255
rect 5007 1289 5199 1295
rect 5007 1255 5019 1289
rect 5187 1255 5199 1289
rect 5007 1249 5199 1255
rect 5385 1289 5577 1295
rect 5385 1255 5397 1289
rect 5565 1255 5577 1289
rect 5385 1249 5577 1255
rect 5763 1289 5955 1295
rect 5763 1255 5775 1289
rect 5943 1255 5955 1289
rect 5763 1249 5955 1255
rect 6141 1289 6333 1295
rect 6141 1255 6153 1289
rect 6321 1255 6333 1289
rect 6141 1249 6333 1255
rect 6519 1289 6711 1295
rect 6519 1255 6531 1289
rect 6699 1255 6711 1289
rect 6519 1249 6711 1255
rect 6897 1289 7089 1295
rect 6897 1255 6909 1289
rect 7077 1255 7089 1289
rect 6897 1249 7089 1255
rect 7275 1289 7467 1295
rect 7275 1255 7287 1289
rect 7455 1255 7467 1289
rect 7275 1249 7467 1255
rect 7653 1289 7845 1295
rect 7653 1255 7665 1289
rect 7833 1255 7845 1289
rect 7653 1249 7845 1255
rect 8031 1289 8223 1295
rect 8031 1255 8043 1289
rect 8211 1255 8223 1289
rect 8031 1249 8223 1255
rect 8409 1289 8601 1295
rect 8409 1255 8421 1289
rect 8589 1255 8601 1289
rect 8409 1249 8601 1255
rect 8787 1289 8979 1295
rect 8787 1255 8799 1289
rect 8967 1255 8979 1289
rect 8787 1249 8979 1255
rect 9165 1289 9357 1295
rect 9165 1255 9177 1289
rect 9345 1255 9357 1289
rect 9165 1249 9357 1255
rect -9357 1181 -9165 1187
rect -9357 1147 -9345 1181
rect -9177 1147 -9165 1181
rect -9357 1141 -9165 1147
rect -8979 1181 -8787 1187
rect -8979 1147 -8967 1181
rect -8799 1147 -8787 1181
rect -8979 1141 -8787 1147
rect -8601 1181 -8409 1187
rect -8601 1147 -8589 1181
rect -8421 1147 -8409 1181
rect -8601 1141 -8409 1147
rect -8223 1181 -8031 1187
rect -8223 1147 -8211 1181
rect -8043 1147 -8031 1181
rect -8223 1141 -8031 1147
rect -7845 1181 -7653 1187
rect -7845 1147 -7833 1181
rect -7665 1147 -7653 1181
rect -7845 1141 -7653 1147
rect -7467 1181 -7275 1187
rect -7467 1147 -7455 1181
rect -7287 1147 -7275 1181
rect -7467 1141 -7275 1147
rect -7089 1181 -6897 1187
rect -7089 1147 -7077 1181
rect -6909 1147 -6897 1181
rect -7089 1141 -6897 1147
rect -6711 1181 -6519 1187
rect -6711 1147 -6699 1181
rect -6531 1147 -6519 1181
rect -6711 1141 -6519 1147
rect -6333 1181 -6141 1187
rect -6333 1147 -6321 1181
rect -6153 1147 -6141 1181
rect -6333 1141 -6141 1147
rect -5955 1181 -5763 1187
rect -5955 1147 -5943 1181
rect -5775 1147 -5763 1181
rect -5955 1141 -5763 1147
rect -5577 1181 -5385 1187
rect -5577 1147 -5565 1181
rect -5397 1147 -5385 1181
rect -5577 1141 -5385 1147
rect -5199 1181 -5007 1187
rect -5199 1147 -5187 1181
rect -5019 1147 -5007 1181
rect -5199 1141 -5007 1147
rect -4821 1181 -4629 1187
rect -4821 1147 -4809 1181
rect -4641 1147 -4629 1181
rect -4821 1141 -4629 1147
rect -4443 1181 -4251 1187
rect -4443 1147 -4431 1181
rect -4263 1147 -4251 1181
rect -4443 1141 -4251 1147
rect -4065 1181 -3873 1187
rect -4065 1147 -4053 1181
rect -3885 1147 -3873 1181
rect -4065 1141 -3873 1147
rect -3687 1181 -3495 1187
rect -3687 1147 -3675 1181
rect -3507 1147 -3495 1181
rect -3687 1141 -3495 1147
rect -3309 1181 -3117 1187
rect -3309 1147 -3297 1181
rect -3129 1147 -3117 1181
rect -3309 1141 -3117 1147
rect -2931 1181 -2739 1187
rect -2931 1147 -2919 1181
rect -2751 1147 -2739 1181
rect -2931 1141 -2739 1147
rect -2553 1181 -2361 1187
rect -2553 1147 -2541 1181
rect -2373 1147 -2361 1181
rect -2553 1141 -2361 1147
rect -2175 1181 -1983 1187
rect -2175 1147 -2163 1181
rect -1995 1147 -1983 1181
rect -2175 1141 -1983 1147
rect -1797 1181 -1605 1187
rect -1797 1147 -1785 1181
rect -1617 1147 -1605 1181
rect -1797 1141 -1605 1147
rect -1419 1181 -1227 1187
rect -1419 1147 -1407 1181
rect -1239 1147 -1227 1181
rect -1419 1141 -1227 1147
rect -1041 1181 -849 1187
rect -1041 1147 -1029 1181
rect -861 1147 -849 1181
rect -1041 1141 -849 1147
rect -663 1181 -471 1187
rect -663 1147 -651 1181
rect -483 1147 -471 1181
rect -663 1141 -471 1147
rect -285 1181 -93 1187
rect -285 1147 -273 1181
rect -105 1147 -93 1181
rect -285 1141 -93 1147
rect 93 1181 285 1187
rect 93 1147 105 1181
rect 273 1147 285 1181
rect 93 1141 285 1147
rect 471 1181 663 1187
rect 471 1147 483 1181
rect 651 1147 663 1181
rect 471 1141 663 1147
rect 849 1181 1041 1187
rect 849 1147 861 1181
rect 1029 1147 1041 1181
rect 849 1141 1041 1147
rect 1227 1181 1419 1187
rect 1227 1147 1239 1181
rect 1407 1147 1419 1181
rect 1227 1141 1419 1147
rect 1605 1181 1797 1187
rect 1605 1147 1617 1181
rect 1785 1147 1797 1181
rect 1605 1141 1797 1147
rect 1983 1181 2175 1187
rect 1983 1147 1995 1181
rect 2163 1147 2175 1181
rect 1983 1141 2175 1147
rect 2361 1181 2553 1187
rect 2361 1147 2373 1181
rect 2541 1147 2553 1181
rect 2361 1141 2553 1147
rect 2739 1181 2931 1187
rect 2739 1147 2751 1181
rect 2919 1147 2931 1181
rect 2739 1141 2931 1147
rect 3117 1181 3309 1187
rect 3117 1147 3129 1181
rect 3297 1147 3309 1181
rect 3117 1141 3309 1147
rect 3495 1181 3687 1187
rect 3495 1147 3507 1181
rect 3675 1147 3687 1181
rect 3495 1141 3687 1147
rect 3873 1181 4065 1187
rect 3873 1147 3885 1181
rect 4053 1147 4065 1181
rect 3873 1141 4065 1147
rect 4251 1181 4443 1187
rect 4251 1147 4263 1181
rect 4431 1147 4443 1181
rect 4251 1141 4443 1147
rect 4629 1181 4821 1187
rect 4629 1147 4641 1181
rect 4809 1147 4821 1181
rect 4629 1141 4821 1147
rect 5007 1181 5199 1187
rect 5007 1147 5019 1181
rect 5187 1147 5199 1181
rect 5007 1141 5199 1147
rect 5385 1181 5577 1187
rect 5385 1147 5397 1181
rect 5565 1147 5577 1181
rect 5385 1141 5577 1147
rect 5763 1181 5955 1187
rect 5763 1147 5775 1181
rect 5943 1147 5955 1181
rect 5763 1141 5955 1147
rect 6141 1181 6333 1187
rect 6141 1147 6153 1181
rect 6321 1147 6333 1181
rect 6141 1141 6333 1147
rect 6519 1181 6711 1187
rect 6519 1147 6531 1181
rect 6699 1147 6711 1181
rect 6519 1141 6711 1147
rect 6897 1181 7089 1187
rect 6897 1147 6909 1181
rect 7077 1147 7089 1181
rect 6897 1141 7089 1147
rect 7275 1181 7467 1187
rect 7275 1147 7287 1181
rect 7455 1147 7467 1181
rect 7275 1141 7467 1147
rect 7653 1181 7845 1187
rect 7653 1147 7665 1181
rect 7833 1147 7845 1181
rect 7653 1141 7845 1147
rect 8031 1181 8223 1187
rect 8031 1147 8043 1181
rect 8211 1147 8223 1181
rect 8031 1141 8223 1147
rect 8409 1181 8601 1187
rect 8409 1147 8421 1181
rect 8589 1147 8601 1181
rect 8409 1141 8601 1147
rect 8787 1181 8979 1187
rect 8787 1147 8799 1181
rect 8967 1147 8979 1181
rect 8787 1141 8979 1147
rect 9165 1181 9357 1187
rect 9165 1147 9177 1181
rect 9345 1147 9357 1181
rect 9165 1141 9357 1147
rect -9413 1097 -9367 1109
rect -9413 121 -9407 1097
rect -9373 121 -9367 1097
rect -9413 109 -9367 121
rect -9155 1097 -9109 1109
rect -9155 121 -9149 1097
rect -9115 121 -9109 1097
rect -9155 109 -9109 121
rect -9035 1097 -8989 1109
rect -9035 121 -9029 1097
rect -8995 121 -8989 1097
rect -9035 109 -8989 121
rect -8777 1097 -8731 1109
rect -8777 121 -8771 1097
rect -8737 121 -8731 1097
rect -8777 109 -8731 121
rect -8657 1097 -8611 1109
rect -8657 121 -8651 1097
rect -8617 121 -8611 1097
rect -8657 109 -8611 121
rect -8399 1097 -8353 1109
rect -8399 121 -8393 1097
rect -8359 121 -8353 1097
rect -8399 109 -8353 121
rect -8279 1097 -8233 1109
rect -8279 121 -8273 1097
rect -8239 121 -8233 1097
rect -8279 109 -8233 121
rect -8021 1097 -7975 1109
rect -8021 121 -8015 1097
rect -7981 121 -7975 1097
rect -8021 109 -7975 121
rect -7901 1097 -7855 1109
rect -7901 121 -7895 1097
rect -7861 121 -7855 1097
rect -7901 109 -7855 121
rect -7643 1097 -7597 1109
rect -7643 121 -7637 1097
rect -7603 121 -7597 1097
rect -7643 109 -7597 121
rect -7523 1097 -7477 1109
rect -7523 121 -7517 1097
rect -7483 121 -7477 1097
rect -7523 109 -7477 121
rect -7265 1097 -7219 1109
rect -7265 121 -7259 1097
rect -7225 121 -7219 1097
rect -7265 109 -7219 121
rect -7145 1097 -7099 1109
rect -7145 121 -7139 1097
rect -7105 121 -7099 1097
rect -7145 109 -7099 121
rect -6887 1097 -6841 1109
rect -6887 121 -6881 1097
rect -6847 121 -6841 1097
rect -6887 109 -6841 121
rect -6767 1097 -6721 1109
rect -6767 121 -6761 1097
rect -6727 121 -6721 1097
rect -6767 109 -6721 121
rect -6509 1097 -6463 1109
rect -6509 121 -6503 1097
rect -6469 121 -6463 1097
rect -6509 109 -6463 121
rect -6389 1097 -6343 1109
rect -6389 121 -6383 1097
rect -6349 121 -6343 1097
rect -6389 109 -6343 121
rect -6131 1097 -6085 1109
rect -6131 121 -6125 1097
rect -6091 121 -6085 1097
rect -6131 109 -6085 121
rect -6011 1097 -5965 1109
rect -6011 121 -6005 1097
rect -5971 121 -5965 1097
rect -6011 109 -5965 121
rect -5753 1097 -5707 1109
rect -5753 121 -5747 1097
rect -5713 121 -5707 1097
rect -5753 109 -5707 121
rect -5633 1097 -5587 1109
rect -5633 121 -5627 1097
rect -5593 121 -5587 1097
rect -5633 109 -5587 121
rect -5375 1097 -5329 1109
rect -5375 121 -5369 1097
rect -5335 121 -5329 1097
rect -5375 109 -5329 121
rect -5255 1097 -5209 1109
rect -5255 121 -5249 1097
rect -5215 121 -5209 1097
rect -5255 109 -5209 121
rect -4997 1097 -4951 1109
rect -4997 121 -4991 1097
rect -4957 121 -4951 1097
rect -4997 109 -4951 121
rect -4877 1097 -4831 1109
rect -4877 121 -4871 1097
rect -4837 121 -4831 1097
rect -4877 109 -4831 121
rect -4619 1097 -4573 1109
rect -4619 121 -4613 1097
rect -4579 121 -4573 1097
rect -4619 109 -4573 121
rect -4499 1097 -4453 1109
rect -4499 121 -4493 1097
rect -4459 121 -4453 1097
rect -4499 109 -4453 121
rect -4241 1097 -4195 1109
rect -4241 121 -4235 1097
rect -4201 121 -4195 1097
rect -4241 109 -4195 121
rect -4121 1097 -4075 1109
rect -4121 121 -4115 1097
rect -4081 121 -4075 1097
rect -4121 109 -4075 121
rect -3863 1097 -3817 1109
rect -3863 121 -3857 1097
rect -3823 121 -3817 1097
rect -3863 109 -3817 121
rect -3743 1097 -3697 1109
rect -3743 121 -3737 1097
rect -3703 121 -3697 1097
rect -3743 109 -3697 121
rect -3485 1097 -3439 1109
rect -3485 121 -3479 1097
rect -3445 121 -3439 1097
rect -3485 109 -3439 121
rect -3365 1097 -3319 1109
rect -3365 121 -3359 1097
rect -3325 121 -3319 1097
rect -3365 109 -3319 121
rect -3107 1097 -3061 1109
rect -3107 121 -3101 1097
rect -3067 121 -3061 1097
rect -3107 109 -3061 121
rect -2987 1097 -2941 1109
rect -2987 121 -2981 1097
rect -2947 121 -2941 1097
rect -2987 109 -2941 121
rect -2729 1097 -2683 1109
rect -2729 121 -2723 1097
rect -2689 121 -2683 1097
rect -2729 109 -2683 121
rect -2609 1097 -2563 1109
rect -2609 121 -2603 1097
rect -2569 121 -2563 1097
rect -2609 109 -2563 121
rect -2351 1097 -2305 1109
rect -2351 121 -2345 1097
rect -2311 121 -2305 1097
rect -2351 109 -2305 121
rect -2231 1097 -2185 1109
rect -2231 121 -2225 1097
rect -2191 121 -2185 1097
rect -2231 109 -2185 121
rect -1973 1097 -1927 1109
rect -1973 121 -1967 1097
rect -1933 121 -1927 1097
rect -1973 109 -1927 121
rect -1853 1097 -1807 1109
rect -1853 121 -1847 1097
rect -1813 121 -1807 1097
rect -1853 109 -1807 121
rect -1595 1097 -1549 1109
rect -1595 121 -1589 1097
rect -1555 121 -1549 1097
rect -1595 109 -1549 121
rect -1475 1097 -1429 1109
rect -1475 121 -1469 1097
rect -1435 121 -1429 1097
rect -1475 109 -1429 121
rect -1217 1097 -1171 1109
rect -1217 121 -1211 1097
rect -1177 121 -1171 1097
rect -1217 109 -1171 121
rect -1097 1097 -1051 1109
rect -1097 121 -1091 1097
rect -1057 121 -1051 1097
rect -1097 109 -1051 121
rect -839 1097 -793 1109
rect -839 121 -833 1097
rect -799 121 -793 1097
rect -839 109 -793 121
rect -719 1097 -673 1109
rect -719 121 -713 1097
rect -679 121 -673 1097
rect -719 109 -673 121
rect -461 1097 -415 1109
rect -461 121 -455 1097
rect -421 121 -415 1097
rect -461 109 -415 121
rect -341 1097 -295 1109
rect -341 121 -335 1097
rect -301 121 -295 1097
rect -341 109 -295 121
rect -83 1097 -37 1109
rect -83 121 -77 1097
rect -43 121 -37 1097
rect -83 109 -37 121
rect 37 1097 83 1109
rect 37 121 43 1097
rect 77 121 83 1097
rect 37 109 83 121
rect 295 1097 341 1109
rect 295 121 301 1097
rect 335 121 341 1097
rect 295 109 341 121
rect 415 1097 461 1109
rect 415 121 421 1097
rect 455 121 461 1097
rect 415 109 461 121
rect 673 1097 719 1109
rect 673 121 679 1097
rect 713 121 719 1097
rect 673 109 719 121
rect 793 1097 839 1109
rect 793 121 799 1097
rect 833 121 839 1097
rect 793 109 839 121
rect 1051 1097 1097 1109
rect 1051 121 1057 1097
rect 1091 121 1097 1097
rect 1051 109 1097 121
rect 1171 1097 1217 1109
rect 1171 121 1177 1097
rect 1211 121 1217 1097
rect 1171 109 1217 121
rect 1429 1097 1475 1109
rect 1429 121 1435 1097
rect 1469 121 1475 1097
rect 1429 109 1475 121
rect 1549 1097 1595 1109
rect 1549 121 1555 1097
rect 1589 121 1595 1097
rect 1549 109 1595 121
rect 1807 1097 1853 1109
rect 1807 121 1813 1097
rect 1847 121 1853 1097
rect 1807 109 1853 121
rect 1927 1097 1973 1109
rect 1927 121 1933 1097
rect 1967 121 1973 1097
rect 1927 109 1973 121
rect 2185 1097 2231 1109
rect 2185 121 2191 1097
rect 2225 121 2231 1097
rect 2185 109 2231 121
rect 2305 1097 2351 1109
rect 2305 121 2311 1097
rect 2345 121 2351 1097
rect 2305 109 2351 121
rect 2563 1097 2609 1109
rect 2563 121 2569 1097
rect 2603 121 2609 1097
rect 2563 109 2609 121
rect 2683 1097 2729 1109
rect 2683 121 2689 1097
rect 2723 121 2729 1097
rect 2683 109 2729 121
rect 2941 1097 2987 1109
rect 2941 121 2947 1097
rect 2981 121 2987 1097
rect 2941 109 2987 121
rect 3061 1097 3107 1109
rect 3061 121 3067 1097
rect 3101 121 3107 1097
rect 3061 109 3107 121
rect 3319 1097 3365 1109
rect 3319 121 3325 1097
rect 3359 121 3365 1097
rect 3319 109 3365 121
rect 3439 1097 3485 1109
rect 3439 121 3445 1097
rect 3479 121 3485 1097
rect 3439 109 3485 121
rect 3697 1097 3743 1109
rect 3697 121 3703 1097
rect 3737 121 3743 1097
rect 3697 109 3743 121
rect 3817 1097 3863 1109
rect 3817 121 3823 1097
rect 3857 121 3863 1097
rect 3817 109 3863 121
rect 4075 1097 4121 1109
rect 4075 121 4081 1097
rect 4115 121 4121 1097
rect 4075 109 4121 121
rect 4195 1097 4241 1109
rect 4195 121 4201 1097
rect 4235 121 4241 1097
rect 4195 109 4241 121
rect 4453 1097 4499 1109
rect 4453 121 4459 1097
rect 4493 121 4499 1097
rect 4453 109 4499 121
rect 4573 1097 4619 1109
rect 4573 121 4579 1097
rect 4613 121 4619 1097
rect 4573 109 4619 121
rect 4831 1097 4877 1109
rect 4831 121 4837 1097
rect 4871 121 4877 1097
rect 4831 109 4877 121
rect 4951 1097 4997 1109
rect 4951 121 4957 1097
rect 4991 121 4997 1097
rect 4951 109 4997 121
rect 5209 1097 5255 1109
rect 5209 121 5215 1097
rect 5249 121 5255 1097
rect 5209 109 5255 121
rect 5329 1097 5375 1109
rect 5329 121 5335 1097
rect 5369 121 5375 1097
rect 5329 109 5375 121
rect 5587 1097 5633 1109
rect 5587 121 5593 1097
rect 5627 121 5633 1097
rect 5587 109 5633 121
rect 5707 1097 5753 1109
rect 5707 121 5713 1097
rect 5747 121 5753 1097
rect 5707 109 5753 121
rect 5965 1097 6011 1109
rect 5965 121 5971 1097
rect 6005 121 6011 1097
rect 5965 109 6011 121
rect 6085 1097 6131 1109
rect 6085 121 6091 1097
rect 6125 121 6131 1097
rect 6085 109 6131 121
rect 6343 1097 6389 1109
rect 6343 121 6349 1097
rect 6383 121 6389 1097
rect 6343 109 6389 121
rect 6463 1097 6509 1109
rect 6463 121 6469 1097
rect 6503 121 6509 1097
rect 6463 109 6509 121
rect 6721 1097 6767 1109
rect 6721 121 6727 1097
rect 6761 121 6767 1097
rect 6721 109 6767 121
rect 6841 1097 6887 1109
rect 6841 121 6847 1097
rect 6881 121 6887 1097
rect 6841 109 6887 121
rect 7099 1097 7145 1109
rect 7099 121 7105 1097
rect 7139 121 7145 1097
rect 7099 109 7145 121
rect 7219 1097 7265 1109
rect 7219 121 7225 1097
rect 7259 121 7265 1097
rect 7219 109 7265 121
rect 7477 1097 7523 1109
rect 7477 121 7483 1097
rect 7517 121 7523 1097
rect 7477 109 7523 121
rect 7597 1097 7643 1109
rect 7597 121 7603 1097
rect 7637 121 7643 1097
rect 7597 109 7643 121
rect 7855 1097 7901 1109
rect 7855 121 7861 1097
rect 7895 121 7901 1097
rect 7855 109 7901 121
rect 7975 1097 8021 1109
rect 7975 121 7981 1097
rect 8015 121 8021 1097
rect 7975 109 8021 121
rect 8233 1097 8279 1109
rect 8233 121 8239 1097
rect 8273 121 8279 1097
rect 8233 109 8279 121
rect 8353 1097 8399 1109
rect 8353 121 8359 1097
rect 8393 121 8399 1097
rect 8353 109 8399 121
rect 8611 1097 8657 1109
rect 8611 121 8617 1097
rect 8651 121 8657 1097
rect 8611 109 8657 121
rect 8731 1097 8777 1109
rect 8731 121 8737 1097
rect 8771 121 8777 1097
rect 8731 109 8777 121
rect 8989 1097 9035 1109
rect 8989 121 8995 1097
rect 9029 121 9035 1097
rect 8989 109 9035 121
rect 9109 1097 9155 1109
rect 9109 121 9115 1097
rect 9149 121 9155 1097
rect 9109 109 9155 121
rect 9367 1097 9413 1109
rect 9367 121 9373 1097
rect 9407 121 9413 1097
rect 9367 109 9413 121
rect -9357 71 -9165 77
rect -9357 37 -9345 71
rect -9177 37 -9165 71
rect -9357 31 -9165 37
rect -8979 71 -8787 77
rect -8979 37 -8967 71
rect -8799 37 -8787 71
rect -8979 31 -8787 37
rect -8601 71 -8409 77
rect -8601 37 -8589 71
rect -8421 37 -8409 71
rect -8601 31 -8409 37
rect -8223 71 -8031 77
rect -8223 37 -8211 71
rect -8043 37 -8031 71
rect -8223 31 -8031 37
rect -7845 71 -7653 77
rect -7845 37 -7833 71
rect -7665 37 -7653 71
rect -7845 31 -7653 37
rect -7467 71 -7275 77
rect -7467 37 -7455 71
rect -7287 37 -7275 71
rect -7467 31 -7275 37
rect -7089 71 -6897 77
rect -7089 37 -7077 71
rect -6909 37 -6897 71
rect -7089 31 -6897 37
rect -6711 71 -6519 77
rect -6711 37 -6699 71
rect -6531 37 -6519 71
rect -6711 31 -6519 37
rect -6333 71 -6141 77
rect -6333 37 -6321 71
rect -6153 37 -6141 71
rect -6333 31 -6141 37
rect -5955 71 -5763 77
rect -5955 37 -5943 71
rect -5775 37 -5763 71
rect -5955 31 -5763 37
rect -5577 71 -5385 77
rect -5577 37 -5565 71
rect -5397 37 -5385 71
rect -5577 31 -5385 37
rect -5199 71 -5007 77
rect -5199 37 -5187 71
rect -5019 37 -5007 71
rect -5199 31 -5007 37
rect -4821 71 -4629 77
rect -4821 37 -4809 71
rect -4641 37 -4629 71
rect -4821 31 -4629 37
rect -4443 71 -4251 77
rect -4443 37 -4431 71
rect -4263 37 -4251 71
rect -4443 31 -4251 37
rect -4065 71 -3873 77
rect -4065 37 -4053 71
rect -3885 37 -3873 71
rect -4065 31 -3873 37
rect -3687 71 -3495 77
rect -3687 37 -3675 71
rect -3507 37 -3495 71
rect -3687 31 -3495 37
rect -3309 71 -3117 77
rect -3309 37 -3297 71
rect -3129 37 -3117 71
rect -3309 31 -3117 37
rect -2931 71 -2739 77
rect -2931 37 -2919 71
rect -2751 37 -2739 71
rect -2931 31 -2739 37
rect -2553 71 -2361 77
rect -2553 37 -2541 71
rect -2373 37 -2361 71
rect -2553 31 -2361 37
rect -2175 71 -1983 77
rect -2175 37 -2163 71
rect -1995 37 -1983 71
rect -2175 31 -1983 37
rect -1797 71 -1605 77
rect -1797 37 -1785 71
rect -1617 37 -1605 71
rect -1797 31 -1605 37
rect -1419 71 -1227 77
rect -1419 37 -1407 71
rect -1239 37 -1227 71
rect -1419 31 -1227 37
rect -1041 71 -849 77
rect -1041 37 -1029 71
rect -861 37 -849 71
rect -1041 31 -849 37
rect -663 71 -471 77
rect -663 37 -651 71
rect -483 37 -471 71
rect -663 31 -471 37
rect -285 71 -93 77
rect -285 37 -273 71
rect -105 37 -93 71
rect -285 31 -93 37
rect 93 71 285 77
rect 93 37 105 71
rect 273 37 285 71
rect 93 31 285 37
rect 471 71 663 77
rect 471 37 483 71
rect 651 37 663 71
rect 471 31 663 37
rect 849 71 1041 77
rect 849 37 861 71
rect 1029 37 1041 71
rect 849 31 1041 37
rect 1227 71 1419 77
rect 1227 37 1239 71
rect 1407 37 1419 71
rect 1227 31 1419 37
rect 1605 71 1797 77
rect 1605 37 1617 71
rect 1785 37 1797 71
rect 1605 31 1797 37
rect 1983 71 2175 77
rect 1983 37 1995 71
rect 2163 37 2175 71
rect 1983 31 2175 37
rect 2361 71 2553 77
rect 2361 37 2373 71
rect 2541 37 2553 71
rect 2361 31 2553 37
rect 2739 71 2931 77
rect 2739 37 2751 71
rect 2919 37 2931 71
rect 2739 31 2931 37
rect 3117 71 3309 77
rect 3117 37 3129 71
rect 3297 37 3309 71
rect 3117 31 3309 37
rect 3495 71 3687 77
rect 3495 37 3507 71
rect 3675 37 3687 71
rect 3495 31 3687 37
rect 3873 71 4065 77
rect 3873 37 3885 71
rect 4053 37 4065 71
rect 3873 31 4065 37
rect 4251 71 4443 77
rect 4251 37 4263 71
rect 4431 37 4443 71
rect 4251 31 4443 37
rect 4629 71 4821 77
rect 4629 37 4641 71
rect 4809 37 4821 71
rect 4629 31 4821 37
rect 5007 71 5199 77
rect 5007 37 5019 71
rect 5187 37 5199 71
rect 5007 31 5199 37
rect 5385 71 5577 77
rect 5385 37 5397 71
rect 5565 37 5577 71
rect 5385 31 5577 37
rect 5763 71 5955 77
rect 5763 37 5775 71
rect 5943 37 5955 71
rect 5763 31 5955 37
rect 6141 71 6333 77
rect 6141 37 6153 71
rect 6321 37 6333 71
rect 6141 31 6333 37
rect 6519 71 6711 77
rect 6519 37 6531 71
rect 6699 37 6711 71
rect 6519 31 6711 37
rect 6897 71 7089 77
rect 6897 37 6909 71
rect 7077 37 7089 71
rect 6897 31 7089 37
rect 7275 71 7467 77
rect 7275 37 7287 71
rect 7455 37 7467 71
rect 7275 31 7467 37
rect 7653 71 7845 77
rect 7653 37 7665 71
rect 7833 37 7845 71
rect 7653 31 7845 37
rect 8031 71 8223 77
rect 8031 37 8043 71
rect 8211 37 8223 71
rect 8031 31 8223 37
rect 8409 71 8601 77
rect 8409 37 8421 71
rect 8589 37 8601 71
rect 8409 31 8601 37
rect 8787 71 8979 77
rect 8787 37 8799 71
rect 8967 37 8979 71
rect 8787 31 8979 37
rect 9165 71 9357 77
rect 9165 37 9177 71
rect 9345 37 9357 71
rect 9165 31 9357 37
rect -9357 -37 -9165 -31
rect -9357 -71 -9345 -37
rect -9177 -71 -9165 -37
rect -9357 -77 -9165 -71
rect -8979 -37 -8787 -31
rect -8979 -71 -8967 -37
rect -8799 -71 -8787 -37
rect -8979 -77 -8787 -71
rect -8601 -37 -8409 -31
rect -8601 -71 -8589 -37
rect -8421 -71 -8409 -37
rect -8601 -77 -8409 -71
rect -8223 -37 -8031 -31
rect -8223 -71 -8211 -37
rect -8043 -71 -8031 -37
rect -8223 -77 -8031 -71
rect -7845 -37 -7653 -31
rect -7845 -71 -7833 -37
rect -7665 -71 -7653 -37
rect -7845 -77 -7653 -71
rect -7467 -37 -7275 -31
rect -7467 -71 -7455 -37
rect -7287 -71 -7275 -37
rect -7467 -77 -7275 -71
rect -7089 -37 -6897 -31
rect -7089 -71 -7077 -37
rect -6909 -71 -6897 -37
rect -7089 -77 -6897 -71
rect -6711 -37 -6519 -31
rect -6711 -71 -6699 -37
rect -6531 -71 -6519 -37
rect -6711 -77 -6519 -71
rect -6333 -37 -6141 -31
rect -6333 -71 -6321 -37
rect -6153 -71 -6141 -37
rect -6333 -77 -6141 -71
rect -5955 -37 -5763 -31
rect -5955 -71 -5943 -37
rect -5775 -71 -5763 -37
rect -5955 -77 -5763 -71
rect -5577 -37 -5385 -31
rect -5577 -71 -5565 -37
rect -5397 -71 -5385 -37
rect -5577 -77 -5385 -71
rect -5199 -37 -5007 -31
rect -5199 -71 -5187 -37
rect -5019 -71 -5007 -37
rect -5199 -77 -5007 -71
rect -4821 -37 -4629 -31
rect -4821 -71 -4809 -37
rect -4641 -71 -4629 -37
rect -4821 -77 -4629 -71
rect -4443 -37 -4251 -31
rect -4443 -71 -4431 -37
rect -4263 -71 -4251 -37
rect -4443 -77 -4251 -71
rect -4065 -37 -3873 -31
rect -4065 -71 -4053 -37
rect -3885 -71 -3873 -37
rect -4065 -77 -3873 -71
rect -3687 -37 -3495 -31
rect -3687 -71 -3675 -37
rect -3507 -71 -3495 -37
rect -3687 -77 -3495 -71
rect -3309 -37 -3117 -31
rect -3309 -71 -3297 -37
rect -3129 -71 -3117 -37
rect -3309 -77 -3117 -71
rect -2931 -37 -2739 -31
rect -2931 -71 -2919 -37
rect -2751 -71 -2739 -37
rect -2931 -77 -2739 -71
rect -2553 -37 -2361 -31
rect -2553 -71 -2541 -37
rect -2373 -71 -2361 -37
rect -2553 -77 -2361 -71
rect -2175 -37 -1983 -31
rect -2175 -71 -2163 -37
rect -1995 -71 -1983 -37
rect -2175 -77 -1983 -71
rect -1797 -37 -1605 -31
rect -1797 -71 -1785 -37
rect -1617 -71 -1605 -37
rect -1797 -77 -1605 -71
rect -1419 -37 -1227 -31
rect -1419 -71 -1407 -37
rect -1239 -71 -1227 -37
rect -1419 -77 -1227 -71
rect -1041 -37 -849 -31
rect -1041 -71 -1029 -37
rect -861 -71 -849 -37
rect -1041 -77 -849 -71
rect -663 -37 -471 -31
rect -663 -71 -651 -37
rect -483 -71 -471 -37
rect -663 -77 -471 -71
rect -285 -37 -93 -31
rect -285 -71 -273 -37
rect -105 -71 -93 -37
rect -285 -77 -93 -71
rect 93 -37 285 -31
rect 93 -71 105 -37
rect 273 -71 285 -37
rect 93 -77 285 -71
rect 471 -37 663 -31
rect 471 -71 483 -37
rect 651 -71 663 -37
rect 471 -77 663 -71
rect 849 -37 1041 -31
rect 849 -71 861 -37
rect 1029 -71 1041 -37
rect 849 -77 1041 -71
rect 1227 -37 1419 -31
rect 1227 -71 1239 -37
rect 1407 -71 1419 -37
rect 1227 -77 1419 -71
rect 1605 -37 1797 -31
rect 1605 -71 1617 -37
rect 1785 -71 1797 -37
rect 1605 -77 1797 -71
rect 1983 -37 2175 -31
rect 1983 -71 1995 -37
rect 2163 -71 2175 -37
rect 1983 -77 2175 -71
rect 2361 -37 2553 -31
rect 2361 -71 2373 -37
rect 2541 -71 2553 -37
rect 2361 -77 2553 -71
rect 2739 -37 2931 -31
rect 2739 -71 2751 -37
rect 2919 -71 2931 -37
rect 2739 -77 2931 -71
rect 3117 -37 3309 -31
rect 3117 -71 3129 -37
rect 3297 -71 3309 -37
rect 3117 -77 3309 -71
rect 3495 -37 3687 -31
rect 3495 -71 3507 -37
rect 3675 -71 3687 -37
rect 3495 -77 3687 -71
rect 3873 -37 4065 -31
rect 3873 -71 3885 -37
rect 4053 -71 4065 -37
rect 3873 -77 4065 -71
rect 4251 -37 4443 -31
rect 4251 -71 4263 -37
rect 4431 -71 4443 -37
rect 4251 -77 4443 -71
rect 4629 -37 4821 -31
rect 4629 -71 4641 -37
rect 4809 -71 4821 -37
rect 4629 -77 4821 -71
rect 5007 -37 5199 -31
rect 5007 -71 5019 -37
rect 5187 -71 5199 -37
rect 5007 -77 5199 -71
rect 5385 -37 5577 -31
rect 5385 -71 5397 -37
rect 5565 -71 5577 -37
rect 5385 -77 5577 -71
rect 5763 -37 5955 -31
rect 5763 -71 5775 -37
rect 5943 -71 5955 -37
rect 5763 -77 5955 -71
rect 6141 -37 6333 -31
rect 6141 -71 6153 -37
rect 6321 -71 6333 -37
rect 6141 -77 6333 -71
rect 6519 -37 6711 -31
rect 6519 -71 6531 -37
rect 6699 -71 6711 -37
rect 6519 -77 6711 -71
rect 6897 -37 7089 -31
rect 6897 -71 6909 -37
rect 7077 -71 7089 -37
rect 6897 -77 7089 -71
rect 7275 -37 7467 -31
rect 7275 -71 7287 -37
rect 7455 -71 7467 -37
rect 7275 -77 7467 -71
rect 7653 -37 7845 -31
rect 7653 -71 7665 -37
rect 7833 -71 7845 -37
rect 7653 -77 7845 -71
rect 8031 -37 8223 -31
rect 8031 -71 8043 -37
rect 8211 -71 8223 -37
rect 8031 -77 8223 -71
rect 8409 -37 8601 -31
rect 8409 -71 8421 -37
rect 8589 -71 8601 -37
rect 8409 -77 8601 -71
rect 8787 -37 8979 -31
rect 8787 -71 8799 -37
rect 8967 -71 8979 -37
rect 8787 -77 8979 -71
rect 9165 -37 9357 -31
rect 9165 -71 9177 -37
rect 9345 -71 9357 -37
rect 9165 -77 9357 -71
rect -9413 -121 -9367 -109
rect -9413 -1097 -9407 -121
rect -9373 -1097 -9367 -121
rect -9413 -1109 -9367 -1097
rect -9155 -121 -9109 -109
rect -9155 -1097 -9149 -121
rect -9115 -1097 -9109 -121
rect -9155 -1109 -9109 -1097
rect -9035 -121 -8989 -109
rect -9035 -1097 -9029 -121
rect -8995 -1097 -8989 -121
rect -9035 -1109 -8989 -1097
rect -8777 -121 -8731 -109
rect -8777 -1097 -8771 -121
rect -8737 -1097 -8731 -121
rect -8777 -1109 -8731 -1097
rect -8657 -121 -8611 -109
rect -8657 -1097 -8651 -121
rect -8617 -1097 -8611 -121
rect -8657 -1109 -8611 -1097
rect -8399 -121 -8353 -109
rect -8399 -1097 -8393 -121
rect -8359 -1097 -8353 -121
rect -8399 -1109 -8353 -1097
rect -8279 -121 -8233 -109
rect -8279 -1097 -8273 -121
rect -8239 -1097 -8233 -121
rect -8279 -1109 -8233 -1097
rect -8021 -121 -7975 -109
rect -8021 -1097 -8015 -121
rect -7981 -1097 -7975 -121
rect -8021 -1109 -7975 -1097
rect -7901 -121 -7855 -109
rect -7901 -1097 -7895 -121
rect -7861 -1097 -7855 -121
rect -7901 -1109 -7855 -1097
rect -7643 -121 -7597 -109
rect -7643 -1097 -7637 -121
rect -7603 -1097 -7597 -121
rect -7643 -1109 -7597 -1097
rect -7523 -121 -7477 -109
rect -7523 -1097 -7517 -121
rect -7483 -1097 -7477 -121
rect -7523 -1109 -7477 -1097
rect -7265 -121 -7219 -109
rect -7265 -1097 -7259 -121
rect -7225 -1097 -7219 -121
rect -7265 -1109 -7219 -1097
rect -7145 -121 -7099 -109
rect -7145 -1097 -7139 -121
rect -7105 -1097 -7099 -121
rect -7145 -1109 -7099 -1097
rect -6887 -121 -6841 -109
rect -6887 -1097 -6881 -121
rect -6847 -1097 -6841 -121
rect -6887 -1109 -6841 -1097
rect -6767 -121 -6721 -109
rect -6767 -1097 -6761 -121
rect -6727 -1097 -6721 -121
rect -6767 -1109 -6721 -1097
rect -6509 -121 -6463 -109
rect -6509 -1097 -6503 -121
rect -6469 -1097 -6463 -121
rect -6509 -1109 -6463 -1097
rect -6389 -121 -6343 -109
rect -6389 -1097 -6383 -121
rect -6349 -1097 -6343 -121
rect -6389 -1109 -6343 -1097
rect -6131 -121 -6085 -109
rect -6131 -1097 -6125 -121
rect -6091 -1097 -6085 -121
rect -6131 -1109 -6085 -1097
rect -6011 -121 -5965 -109
rect -6011 -1097 -6005 -121
rect -5971 -1097 -5965 -121
rect -6011 -1109 -5965 -1097
rect -5753 -121 -5707 -109
rect -5753 -1097 -5747 -121
rect -5713 -1097 -5707 -121
rect -5753 -1109 -5707 -1097
rect -5633 -121 -5587 -109
rect -5633 -1097 -5627 -121
rect -5593 -1097 -5587 -121
rect -5633 -1109 -5587 -1097
rect -5375 -121 -5329 -109
rect -5375 -1097 -5369 -121
rect -5335 -1097 -5329 -121
rect -5375 -1109 -5329 -1097
rect -5255 -121 -5209 -109
rect -5255 -1097 -5249 -121
rect -5215 -1097 -5209 -121
rect -5255 -1109 -5209 -1097
rect -4997 -121 -4951 -109
rect -4997 -1097 -4991 -121
rect -4957 -1097 -4951 -121
rect -4997 -1109 -4951 -1097
rect -4877 -121 -4831 -109
rect -4877 -1097 -4871 -121
rect -4837 -1097 -4831 -121
rect -4877 -1109 -4831 -1097
rect -4619 -121 -4573 -109
rect -4619 -1097 -4613 -121
rect -4579 -1097 -4573 -121
rect -4619 -1109 -4573 -1097
rect -4499 -121 -4453 -109
rect -4499 -1097 -4493 -121
rect -4459 -1097 -4453 -121
rect -4499 -1109 -4453 -1097
rect -4241 -121 -4195 -109
rect -4241 -1097 -4235 -121
rect -4201 -1097 -4195 -121
rect -4241 -1109 -4195 -1097
rect -4121 -121 -4075 -109
rect -4121 -1097 -4115 -121
rect -4081 -1097 -4075 -121
rect -4121 -1109 -4075 -1097
rect -3863 -121 -3817 -109
rect -3863 -1097 -3857 -121
rect -3823 -1097 -3817 -121
rect -3863 -1109 -3817 -1097
rect -3743 -121 -3697 -109
rect -3743 -1097 -3737 -121
rect -3703 -1097 -3697 -121
rect -3743 -1109 -3697 -1097
rect -3485 -121 -3439 -109
rect -3485 -1097 -3479 -121
rect -3445 -1097 -3439 -121
rect -3485 -1109 -3439 -1097
rect -3365 -121 -3319 -109
rect -3365 -1097 -3359 -121
rect -3325 -1097 -3319 -121
rect -3365 -1109 -3319 -1097
rect -3107 -121 -3061 -109
rect -3107 -1097 -3101 -121
rect -3067 -1097 -3061 -121
rect -3107 -1109 -3061 -1097
rect -2987 -121 -2941 -109
rect -2987 -1097 -2981 -121
rect -2947 -1097 -2941 -121
rect -2987 -1109 -2941 -1097
rect -2729 -121 -2683 -109
rect -2729 -1097 -2723 -121
rect -2689 -1097 -2683 -121
rect -2729 -1109 -2683 -1097
rect -2609 -121 -2563 -109
rect -2609 -1097 -2603 -121
rect -2569 -1097 -2563 -121
rect -2609 -1109 -2563 -1097
rect -2351 -121 -2305 -109
rect -2351 -1097 -2345 -121
rect -2311 -1097 -2305 -121
rect -2351 -1109 -2305 -1097
rect -2231 -121 -2185 -109
rect -2231 -1097 -2225 -121
rect -2191 -1097 -2185 -121
rect -2231 -1109 -2185 -1097
rect -1973 -121 -1927 -109
rect -1973 -1097 -1967 -121
rect -1933 -1097 -1927 -121
rect -1973 -1109 -1927 -1097
rect -1853 -121 -1807 -109
rect -1853 -1097 -1847 -121
rect -1813 -1097 -1807 -121
rect -1853 -1109 -1807 -1097
rect -1595 -121 -1549 -109
rect -1595 -1097 -1589 -121
rect -1555 -1097 -1549 -121
rect -1595 -1109 -1549 -1097
rect -1475 -121 -1429 -109
rect -1475 -1097 -1469 -121
rect -1435 -1097 -1429 -121
rect -1475 -1109 -1429 -1097
rect -1217 -121 -1171 -109
rect -1217 -1097 -1211 -121
rect -1177 -1097 -1171 -121
rect -1217 -1109 -1171 -1097
rect -1097 -121 -1051 -109
rect -1097 -1097 -1091 -121
rect -1057 -1097 -1051 -121
rect -1097 -1109 -1051 -1097
rect -839 -121 -793 -109
rect -839 -1097 -833 -121
rect -799 -1097 -793 -121
rect -839 -1109 -793 -1097
rect -719 -121 -673 -109
rect -719 -1097 -713 -121
rect -679 -1097 -673 -121
rect -719 -1109 -673 -1097
rect -461 -121 -415 -109
rect -461 -1097 -455 -121
rect -421 -1097 -415 -121
rect -461 -1109 -415 -1097
rect -341 -121 -295 -109
rect -341 -1097 -335 -121
rect -301 -1097 -295 -121
rect -341 -1109 -295 -1097
rect -83 -121 -37 -109
rect -83 -1097 -77 -121
rect -43 -1097 -37 -121
rect -83 -1109 -37 -1097
rect 37 -121 83 -109
rect 37 -1097 43 -121
rect 77 -1097 83 -121
rect 37 -1109 83 -1097
rect 295 -121 341 -109
rect 295 -1097 301 -121
rect 335 -1097 341 -121
rect 295 -1109 341 -1097
rect 415 -121 461 -109
rect 415 -1097 421 -121
rect 455 -1097 461 -121
rect 415 -1109 461 -1097
rect 673 -121 719 -109
rect 673 -1097 679 -121
rect 713 -1097 719 -121
rect 673 -1109 719 -1097
rect 793 -121 839 -109
rect 793 -1097 799 -121
rect 833 -1097 839 -121
rect 793 -1109 839 -1097
rect 1051 -121 1097 -109
rect 1051 -1097 1057 -121
rect 1091 -1097 1097 -121
rect 1051 -1109 1097 -1097
rect 1171 -121 1217 -109
rect 1171 -1097 1177 -121
rect 1211 -1097 1217 -121
rect 1171 -1109 1217 -1097
rect 1429 -121 1475 -109
rect 1429 -1097 1435 -121
rect 1469 -1097 1475 -121
rect 1429 -1109 1475 -1097
rect 1549 -121 1595 -109
rect 1549 -1097 1555 -121
rect 1589 -1097 1595 -121
rect 1549 -1109 1595 -1097
rect 1807 -121 1853 -109
rect 1807 -1097 1813 -121
rect 1847 -1097 1853 -121
rect 1807 -1109 1853 -1097
rect 1927 -121 1973 -109
rect 1927 -1097 1933 -121
rect 1967 -1097 1973 -121
rect 1927 -1109 1973 -1097
rect 2185 -121 2231 -109
rect 2185 -1097 2191 -121
rect 2225 -1097 2231 -121
rect 2185 -1109 2231 -1097
rect 2305 -121 2351 -109
rect 2305 -1097 2311 -121
rect 2345 -1097 2351 -121
rect 2305 -1109 2351 -1097
rect 2563 -121 2609 -109
rect 2563 -1097 2569 -121
rect 2603 -1097 2609 -121
rect 2563 -1109 2609 -1097
rect 2683 -121 2729 -109
rect 2683 -1097 2689 -121
rect 2723 -1097 2729 -121
rect 2683 -1109 2729 -1097
rect 2941 -121 2987 -109
rect 2941 -1097 2947 -121
rect 2981 -1097 2987 -121
rect 2941 -1109 2987 -1097
rect 3061 -121 3107 -109
rect 3061 -1097 3067 -121
rect 3101 -1097 3107 -121
rect 3061 -1109 3107 -1097
rect 3319 -121 3365 -109
rect 3319 -1097 3325 -121
rect 3359 -1097 3365 -121
rect 3319 -1109 3365 -1097
rect 3439 -121 3485 -109
rect 3439 -1097 3445 -121
rect 3479 -1097 3485 -121
rect 3439 -1109 3485 -1097
rect 3697 -121 3743 -109
rect 3697 -1097 3703 -121
rect 3737 -1097 3743 -121
rect 3697 -1109 3743 -1097
rect 3817 -121 3863 -109
rect 3817 -1097 3823 -121
rect 3857 -1097 3863 -121
rect 3817 -1109 3863 -1097
rect 4075 -121 4121 -109
rect 4075 -1097 4081 -121
rect 4115 -1097 4121 -121
rect 4075 -1109 4121 -1097
rect 4195 -121 4241 -109
rect 4195 -1097 4201 -121
rect 4235 -1097 4241 -121
rect 4195 -1109 4241 -1097
rect 4453 -121 4499 -109
rect 4453 -1097 4459 -121
rect 4493 -1097 4499 -121
rect 4453 -1109 4499 -1097
rect 4573 -121 4619 -109
rect 4573 -1097 4579 -121
rect 4613 -1097 4619 -121
rect 4573 -1109 4619 -1097
rect 4831 -121 4877 -109
rect 4831 -1097 4837 -121
rect 4871 -1097 4877 -121
rect 4831 -1109 4877 -1097
rect 4951 -121 4997 -109
rect 4951 -1097 4957 -121
rect 4991 -1097 4997 -121
rect 4951 -1109 4997 -1097
rect 5209 -121 5255 -109
rect 5209 -1097 5215 -121
rect 5249 -1097 5255 -121
rect 5209 -1109 5255 -1097
rect 5329 -121 5375 -109
rect 5329 -1097 5335 -121
rect 5369 -1097 5375 -121
rect 5329 -1109 5375 -1097
rect 5587 -121 5633 -109
rect 5587 -1097 5593 -121
rect 5627 -1097 5633 -121
rect 5587 -1109 5633 -1097
rect 5707 -121 5753 -109
rect 5707 -1097 5713 -121
rect 5747 -1097 5753 -121
rect 5707 -1109 5753 -1097
rect 5965 -121 6011 -109
rect 5965 -1097 5971 -121
rect 6005 -1097 6011 -121
rect 5965 -1109 6011 -1097
rect 6085 -121 6131 -109
rect 6085 -1097 6091 -121
rect 6125 -1097 6131 -121
rect 6085 -1109 6131 -1097
rect 6343 -121 6389 -109
rect 6343 -1097 6349 -121
rect 6383 -1097 6389 -121
rect 6343 -1109 6389 -1097
rect 6463 -121 6509 -109
rect 6463 -1097 6469 -121
rect 6503 -1097 6509 -121
rect 6463 -1109 6509 -1097
rect 6721 -121 6767 -109
rect 6721 -1097 6727 -121
rect 6761 -1097 6767 -121
rect 6721 -1109 6767 -1097
rect 6841 -121 6887 -109
rect 6841 -1097 6847 -121
rect 6881 -1097 6887 -121
rect 6841 -1109 6887 -1097
rect 7099 -121 7145 -109
rect 7099 -1097 7105 -121
rect 7139 -1097 7145 -121
rect 7099 -1109 7145 -1097
rect 7219 -121 7265 -109
rect 7219 -1097 7225 -121
rect 7259 -1097 7265 -121
rect 7219 -1109 7265 -1097
rect 7477 -121 7523 -109
rect 7477 -1097 7483 -121
rect 7517 -1097 7523 -121
rect 7477 -1109 7523 -1097
rect 7597 -121 7643 -109
rect 7597 -1097 7603 -121
rect 7637 -1097 7643 -121
rect 7597 -1109 7643 -1097
rect 7855 -121 7901 -109
rect 7855 -1097 7861 -121
rect 7895 -1097 7901 -121
rect 7855 -1109 7901 -1097
rect 7975 -121 8021 -109
rect 7975 -1097 7981 -121
rect 8015 -1097 8021 -121
rect 7975 -1109 8021 -1097
rect 8233 -121 8279 -109
rect 8233 -1097 8239 -121
rect 8273 -1097 8279 -121
rect 8233 -1109 8279 -1097
rect 8353 -121 8399 -109
rect 8353 -1097 8359 -121
rect 8393 -1097 8399 -121
rect 8353 -1109 8399 -1097
rect 8611 -121 8657 -109
rect 8611 -1097 8617 -121
rect 8651 -1097 8657 -121
rect 8611 -1109 8657 -1097
rect 8731 -121 8777 -109
rect 8731 -1097 8737 -121
rect 8771 -1097 8777 -121
rect 8731 -1109 8777 -1097
rect 8989 -121 9035 -109
rect 8989 -1097 8995 -121
rect 9029 -1097 9035 -121
rect 8989 -1109 9035 -1097
rect 9109 -121 9155 -109
rect 9109 -1097 9115 -121
rect 9149 -1097 9155 -121
rect 9109 -1109 9155 -1097
rect 9367 -121 9413 -109
rect 9367 -1097 9373 -121
rect 9407 -1097 9413 -121
rect 9367 -1109 9413 -1097
rect -9357 -1147 -9165 -1141
rect -9357 -1181 -9345 -1147
rect -9177 -1181 -9165 -1147
rect -9357 -1187 -9165 -1181
rect -8979 -1147 -8787 -1141
rect -8979 -1181 -8967 -1147
rect -8799 -1181 -8787 -1147
rect -8979 -1187 -8787 -1181
rect -8601 -1147 -8409 -1141
rect -8601 -1181 -8589 -1147
rect -8421 -1181 -8409 -1147
rect -8601 -1187 -8409 -1181
rect -8223 -1147 -8031 -1141
rect -8223 -1181 -8211 -1147
rect -8043 -1181 -8031 -1147
rect -8223 -1187 -8031 -1181
rect -7845 -1147 -7653 -1141
rect -7845 -1181 -7833 -1147
rect -7665 -1181 -7653 -1147
rect -7845 -1187 -7653 -1181
rect -7467 -1147 -7275 -1141
rect -7467 -1181 -7455 -1147
rect -7287 -1181 -7275 -1147
rect -7467 -1187 -7275 -1181
rect -7089 -1147 -6897 -1141
rect -7089 -1181 -7077 -1147
rect -6909 -1181 -6897 -1147
rect -7089 -1187 -6897 -1181
rect -6711 -1147 -6519 -1141
rect -6711 -1181 -6699 -1147
rect -6531 -1181 -6519 -1147
rect -6711 -1187 -6519 -1181
rect -6333 -1147 -6141 -1141
rect -6333 -1181 -6321 -1147
rect -6153 -1181 -6141 -1147
rect -6333 -1187 -6141 -1181
rect -5955 -1147 -5763 -1141
rect -5955 -1181 -5943 -1147
rect -5775 -1181 -5763 -1147
rect -5955 -1187 -5763 -1181
rect -5577 -1147 -5385 -1141
rect -5577 -1181 -5565 -1147
rect -5397 -1181 -5385 -1147
rect -5577 -1187 -5385 -1181
rect -5199 -1147 -5007 -1141
rect -5199 -1181 -5187 -1147
rect -5019 -1181 -5007 -1147
rect -5199 -1187 -5007 -1181
rect -4821 -1147 -4629 -1141
rect -4821 -1181 -4809 -1147
rect -4641 -1181 -4629 -1147
rect -4821 -1187 -4629 -1181
rect -4443 -1147 -4251 -1141
rect -4443 -1181 -4431 -1147
rect -4263 -1181 -4251 -1147
rect -4443 -1187 -4251 -1181
rect -4065 -1147 -3873 -1141
rect -4065 -1181 -4053 -1147
rect -3885 -1181 -3873 -1147
rect -4065 -1187 -3873 -1181
rect -3687 -1147 -3495 -1141
rect -3687 -1181 -3675 -1147
rect -3507 -1181 -3495 -1147
rect -3687 -1187 -3495 -1181
rect -3309 -1147 -3117 -1141
rect -3309 -1181 -3297 -1147
rect -3129 -1181 -3117 -1147
rect -3309 -1187 -3117 -1181
rect -2931 -1147 -2739 -1141
rect -2931 -1181 -2919 -1147
rect -2751 -1181 -2739 -1147
rect -2931 -1187 -2739 -1181
rect -2553 -1147 -2361 -1141
rect -2553 -1181 -2541 -1147
rect -2373 -1181 -2361 -1147
rect -2553 -1187 -2361 -1181
rect -2175 -1147 -1983 -1141
rect -2175 -1181 -2163 -1147
rect -1995 -1181 -1983 -1147
rect -2175 -1187 -1983 -1181
rect -1797 -1147 -1605 -1141
rect -1797 -1181 -1785 -1147
rect -1617 -1181 -1605 -1147
rect -1797 -1187 -1605 -1181
rect -1419 -1147 -1227 -1141
rect -1419 -1181 -1407 -1147
rect -1239 -1181 -1227 -1147
rect -1419 -1187 -1227 -1181
rect -1041 -1147 -849 -1141
rect -1041 -1181 -1029 -1147
rect -861 -1181 -849 -1147
rect -1041 -1187 -849 -1181
rect -663 -1147 -471 -1141
rect -663 -1181 -651 -1147
rect -483 -1181 -471 -1147
rect -663 -1187 -471 -1181
rect -285 -1147 -93 -1141
rect -285 -1181 -273 -1147
rect -105 -1181 -93 -1147
rect -285 -1187 -93 -1181
rect 93 -1147 285 -1141
rect 93 -1181 105 -1147
rect 273 -1181 285 -1147
rect 93 -1187 285 -1181
rect 471 -1147 663 -1141
rect 471 -1181 483 -1147
rect 651 -1181 663 -1147
rect 471 -1187 663 -1181
rect 849 -1147 1041 -1141
rect 849 -1181 861 -1147
rect 1029 -1181 1041 -1147
rect 849 -1187 1041 -1181
rect 1227 -1147 1419 -1141
rect 1227 -1181 1239 -1147
rect 1407 -1181 1419 -1147
rect 1227 -1187 1419 -1181
rect 1605 -1147 1797 -1141
rect 1605 -1181 1617 -1147
rect 1785 -1181 1797 -1147
rect 1605 -1187 1797 -1181
rect 1983 -1147 2175 -1141
rect 1983 -1181 1995 -1147
rect 2163 -1181 2175 -1147
rect 1983 -1187 2175 -1181
rect 2361 -1147 2553 -1141
rect 2361 -1181 2373 -1147
rect 2541 -1181 2553 -1147
rect 2361 -1187 2553 -1181
rect 2739 -1147 2931 -1141
rect 2739 -1181 2751 -1147
rect 2919 -1181 2931 -1147
rect 2739 -1187 2931 -1181
rect 3117 -1147 3309 -1141
rect 3117 -1181 3129 -1147
rect 3297 -1181 3309 -1147
rect 3117 -1187 3309 -1181
rect 3495 -1147 3687 -1141
rect 3495 -1181 3507 -1147
rect 3675 -1181 3687 -1147
rect 3495 -1187 3687 -1181
rect 3873 -1147 4065 -1141
rect 3873 -1181 3885 -1147
rect 4053 -1181 4065 -1147
rect 3873 -1187 4065 -1181
rect 4251 -1147 4443 -1141
rect 4251 -1181 4263 -1147
rect 4431 -1181 4443 -1147
rect 4251 -1187 4443 -1181
rect 4629 -1147 4821 -1141
rect 4629 -1181 4641 -1147
rect 4809 -1181 4821 -1147
rect 4629 -1187 4821 -1181
rect 5007 -1147 5199 -1141
rect 5007 -1181 5019 -1147
rect 5187 -1181 5199 -1147
rect 5007 -1187 5199 -1181
rect 5385 -1147 5577 -1141
rect 5385 -1181 5397 -1147
rect 5565 -1181 5577 -1147
rect 5385 -1187 5577 -1181
rect 5763 -1147 5955 -1141
rect 5763 -1181 5775 -1147
rect 5943 -1181 5955 -1147
rect 5763 -1187 5955 -1181
rect 6141 -1147 6333 -1141
rect 6141 -1181 6153 -1147
rect 6321 -1181 6333 -1147
rect 6141 -1187 6333 -1181
rect 6519 -1147 6711 -1141
rect 6519 -1181 6531 -1147
rect 6699 -1181 6711 -1147
rect 6519 -1187 6711 -1181
rect 6897 -1147 7089 -1141
rect 6897 -1181 6909 -1147
rect 7077 -1181 7089 -1147
rect 6897 -1187 7089 -1181
rect 7275 -1147 7467 -1141
rect 7275 -1181 7287 -1147
rect 7455 -1181 7467 -1147
rect 7275 -1187 7467 -1181
rect 7653 -1147 7845 -1141
rect 7653 -1181 7665 -1147
rect 7833 -1181 7845 -1147
rect 7653 -1187 7845 -1181
rect 8031 -1147 8223 -1141
rect 8031 -1181 8043 -1147
rect 8211 -1181 8223 -1147
rect 8031 -1187 8223 -1181
rect 8409 -1147 8601 -1141
rect 8409 -1181 8421 -1147
rect 8589 -1181 8601 -1147
rect 8409 -1187 8601 -1181
rect 8787 -1147 8979 -1141
rect 8787 -1181 8799 -1147
rect 8967 -1181 8979 -1147
rect 8787 -1187 8979 -1181
rect 9165 -1147 9357 -1141
rect 9165 -1181 9177 -1147
rect 9345 -1181 9357 -1147
rect 9165 -1187 9357 -1181
rect -9357 -1255 -9165 -1249
rect -9357 -1289 -9345 -1255
rect -9177 -1289 -9165 -1255
rect -9357 -1295 -9165 -1289
rect -8979 -1255 -8787 -1249
rect -8979 -1289 -8967 -1255
rect -8799 -1289 -8787 -1255
rect -8979 -1295 -8787 -1289
rect -8601 -1255 -8409 -1249
rect -8601 -1289 -8589 -1255
rect -8421 -1289 -8409 -1255
rect -8601 -1295 -8409 -1289
rect -8223 -1255 -8031 -1249
rect -8223 -1289 -8211 -1255
rect -8043 -1289 -8031 -1255
rect -8223 -1295 -8031 -1289
rect -7845 -1255 -7653 -1249
rect -7845 -1289 -7833 -1255
rect -7665 -1289 -7653 -1255
rect -7845 -1295 -7653 -1289
rect -7467 -1255 -7275 -1249
rect -7467 -1289 -7455 -1255
rect -7287 -1289 -7275 -1255
rect -7467 -1295 -7275 -1289
rect -7089 -1255 -6897 -1249
rect -7089 -1289 -7077 -1255
rect -6909 -1289 -6897 -1255
rect -7089 -1295 -6897 -1289
rect -6711 -1255 -6519 -1249
rect -6711 -1289 -6699 -1255
rect -6531 -1289 -6519 -1255
rect -6711 -1295 -6519 -1289
rect -6333 -1255 -6141 -1249
rect -6333 -1289 -6321 -1255
rect -6153 -1289 -6141 -1255
rect -6333 -1295 -6141 -1289
rect -5955 -1255 -5763 -1249
rect -5955 -1289 -5943 -1255
rect -5775 -1289 -5763 -1255
rect -5955 -1295 -5763 -1289
rect -5577 -1255 -5385 -1249
rect -5577 -1289 -5565 -1255
rect -5397 -1289 -5385 -1255
rect -5577 -1295 -5385 -1289
rect -5199 -1255 -5007 -1249
rect -5199 -1289 -5187 -1255
rect -5019 -1289 -5007 -1255
rect -5199 -1295 -5007 -1289
rect -4821 -1255 -4629 -1249
rect -4821 -1289 -4809 -1255
rect -4641 -1289 -4629 -1255
rect -4821 -1295 -4629 -1289
rect -4443 -1255 -4251 -1249
rect -4443 -1289 -4431 -1255
rect -4263 -1289 -4251 -1255
rect -4443 -1295 -4251 -1289
rect -4065 -1255 -3873 -1249
rect -4065 -1289 -4053 -1255
rect -3885 -1289 -3873 -1255
rect -4065 -1295 -3873 -1289
rect -3687 -1255 -3495 -1249
rect -3687 -1289 -3675 -1255
rect -3507 -1289 -3495 -1255
rect -3687 -1295 -3495 -1289
rect -3309 -1255 -3117 -1249
rect -3309 -1289 -3297 -1255
rect -3129 -1289 -3117 -1255
rect -3309 -1295 -3117 -1289
rect -2931 -1255 -2739 -1249
rect -2931 -1289 -2919 -1255
rect -2751 -1289 -2739 -1255
rect -2931 -1295 -2739 -1289
rect -2553 -1255 -2361 -1249
rect -2553 -1289 -2541 -1255
rect -2373 -1289 -2361 -1255
rect -2553 -1295 -2361 -1289
rect -2175 -1255 -1983 -1249
rect -2175 -1289 -2163 -1255
rect -1995 -1289 -1983 -1255
rect -2175 -1295 -1983 -1289
rect -1797 -1255 -1605 -1249
rect -1797 -1289 -1785 -1255
rect -1617 -1289 -1605 -1255
rect -1797 -1295 -1605 -1289
rect -1419 -1255 -1227 -1249
rect -1419 -1289 -1407 -1255
rect -1239 -1289 -1227 -1255
rect -1419 -1295 -1227 -1289
rect -1041 -1255 -849 -1249
rect -1041 -1289 -1029 -1255
rect -861 -1289 -849 -1255
rect -1041 -1295 -849 -1289
rect -663 -1255 -471 -1249
rect -663 -1289 -651 -1255
rect -483 -1289 -471 -1255
rect -663 -1295 -471 -1289
rect -285 -1255 -93 -1249
rect -285 -1289 -273 -1255
rect -105 -1289 -93 -1255
rect -285 -1295 -93 -1289
rect 93 -1255 285 -1249
rect 93 -1289 105 -1255
rect 273 -1289 285 -1255
rect 93 -1295 285 -1289
rect 471 -1255 663 -1249
rect 471 -1289 483 -1255
rect 651 -1289 663 -1255
rect 471 -1295 663 -1289
rect 849 -1255 1041 -1249
rect 849 -1289 861 -1255
rect 1029 -1289 1041 -1255
rect 849 -1295 1041 -1289
rect 1227 -1255 1419 -1249
rect 1227 -1289 1239 -1255
rect 1407 -1289 1419 -1255
rect 1227 -1295 1419 -1289
rect 1605 -1255 1797 -1249
rect 1605 -1289 1617 -1255
rect 1785 -1289 1797 -1255
rect 1605 -1295 1797 -1289
rect 1983 -1255 2175 -1249
rect 1983 -1289 1995 -1255
rect 2163 -1289 2175 -1255
rect 1983 -1295 2175 -1289
rect 2361 -1255 2553 -1249
rect 2361 -1289 2373 -1255
rect 2541 -1289 2553 -1255
rect 2361 -1295 2553 -1289
rect 2739 -1255 2931 -1249
rect 2739 -1289 2751 -1255
rect 2919 -1289 2931 -1255
rect 2739 -1295 2931 -1289
rect 3117 -1255 3309 -1249
rect 3117 -1289 3129 -1255
rect 3297 -1289 3309 -1255
rect 3117 -1295 3309 -1289
rect 3495 -1255 3687 -1249
rect 3495 -1289 3507 -1255
rect 3675 -1289 3687 -1255
rect 3495 -1295 3687 -1289
rect 3873 -1255 4065 -1249
rect 3873 -1289 3885 -1255
rect 4053 -1289 4065 -1255
rect 3873 -1295 4065 -1289
rect 4251 -1255 4443 -1249
rect 4251 -1289 4263 -1255
rect 4431 -1289 4443 -1255
rect 4251 -1295 4443 -1289
rect 4629 -1255 4821 -1249
rect 4629 -1289 4641 -1255
rect 4809 -1289 4821 -1255
rect 4629 -1295 4821 -1289
rect 5007 -1255 5199 -1249
rect 5007 -1289 5019 -1255
rect 5187 -1289 5199 -1255
rect 5007 -1295 5199 -1289
rect 5385 -1255 5577 -1249
rect 5385 -1289 5397 -1255
rect 5565 -1289 5577 -1255
rect 5385 -1295 5577 -1289
rect 5763 -1255 5955 -1249
rect 5763 -1289 5775 -1255
rect 5943 -1289 5955 -1255
rect 5763 -1295 5955 -1289
rect 6141 -1255 6333 -1249
rect 6141 -1289 6153 -1255
rect 6321 -1289 6333 -1255
rect 6141 -1295 6333 -1289
rect 6519 -1255 6711 -1249
rect 6519 -1289 6531 -1255
rect 6699 -1289 6711 -1255
rect 6519 -1295 6711 -1289
rect 6897 -1255 7089 -1249
rect 6897 -1289 6909 -1255
rect 7077 -1289 7089 -1255
rect 6897 -1295 7089 -1289
rect 7275 -1255 7467 -1249
rect 7275 -1289 7287 -1255
rect 7455 -1289 7467 -1255
rect 7275 -1295 7467 -1289
rect 7653 -1255 7845 -1249
rect 7653 -1289 7665 -1255
rect 7833 -1289 7845 -1255
rect 7653 -1295 7845 -1289
rect 8031 -1255 8223 -1249
rect 8031 -1289 8043 -1255
rect 8211 -1289 8223 -1255
rect 8031 -1295 8223 -1289
rect 8409 -1255 8601 -1249
rect 8409 -1289 8421 -1255
rect 8589 -1289 8601 -1255
rect 8409 -1295 8601 -1289
rect 8787 -1255 8979 -1249
rect 8787 -1289 8799 -1255
rect 8967 -1289 8979 -1255
rect 8787 -1295 8979 -1289
rect 9165 -1255 9357 -1249
rect 9165 -1289 9177 -1255
rect 9345 -1289 9357 -1255
rect 9165 -1295 9357 -1289
rect -9413 -1339 -9367 -1327
rect -9413 -2315 -9407 -1339
rect -9373 -2315 -9367 -1339
rect -9413 -2327 -9367 -2315
rect -9155 -1339 -9109 -1327
rect -9155 -2315 -9149 -1339
rect -9115 -2315 -9109 -1339
rect -9155 -2327 -9109 -2315
rect -9035 -1339 -8989 -1327
rect -9035 -2315 -9029 -1339
rect -8995 -2315 -8989 -1339
rect -9035 -2327 -8989 -2315
rect -8777 -1339 -8731 -1327
rect -8777 -2315 -8771 -1339
rect -8737 -2315 -8731 -1339
rect -8777 -2327 -8731 -2315
rect -8657 -1339 -8611 -1327
rect -8657 -2315 -8651 -1339
rect -8617 -2315 -8611 -1339
rect -8657 -2327 -8611 -2315
rect -8399 -1339 -8353 -1327
rect -8399 -2315 -8393 -1339
rect -8359 -2315 -8353 -1339
rect -8399 -2327 -8353 -2315
rect -8279 -1339 -8233 -1327
rect -8279 -2315 -8273 -1339
rect -8239 -2315 -8233 -1339
rect -8279 -2327 -8233 -2315
rect -8021 -1339 -7975 -1327
rect -8021 -2315 -8015 -1339
rect -7981 -2315 -7975 -1339
rect -8021 -2327 -7975 -2315
rect -7901 -1339 -7855 -1327
rect -7901 -2315 -7895 -1339
rect -7861 -2315 -7855 -1339
rect -7901 -2327 -7855 -2315
rect -7643 -1339 -7597 -1327
rect -7643 -2315 -7637 -1339
rect -7603 -2315 -7597 -1339
rect -7643 -2327 -7597 -2315
rect -7523 -1339 -7477 -1327
rect -7523 -2315 -7517 -1339
rect -7483 -2315 -7477 -1339
rect -7523 -2327 -7477 -2315
rect -7265 -1339 -7219 -1327
rect -7265 -2315 -7259 -1339
rect -7225 -2315 -7219 -1339
rect -7265 -2327 -7219 -2315
rect -7145 -1339 -7099 -1327
rect -7145 -2315 -7139 -1339
rect -7105 -2315 -7099 -1339
rect -7145 -2327 -7099 -2315
rect -6887 -1339 -6841 -1327
rect -6887 -2315 -6881 -1339
rect -6847 -2315 -6841 -1339
rect -6887 -2327 -6841 -2315
rect -6767 -1339 -6721 -1327
rect -6767 -2315 -6761 -1339
rect -6727 -2315 -6721 -1339
rect -6767 -2327 -6721 -2315
rect -6509 -1339 -6463 -1327
rect -6509 -2315 -6503 -1339
rect -6469 -2315 -6463 -1339
rect -6509 -2327 -6463 -2315
rect -6389 -1339 -6343 -1327
rect -6389 -2315 -6383 -1339
rect -6349 -2315 -6343 -1339
rect -6389 -2327 -6343 -2315
rect -6131 -1339 -6085 -1327
rect -6131 -2315 -6125 -1339
rect -6091 -2315 -6085 -1339
rect -6131 -2327 -6085 -2315
rect -6011 -1339 -5965 -1327
rect -6011 -2315 -6005 -1339
rect -5971 -2315 -5965 -1339
rect -6011 -2327 -5965 -2315
rect -5753 -1339 -5707 -1327
rect -5753 -2315 -5747 -1339
rect -5713 -2315 -5707 -1339
rect -5753 -2327 -5707 -2315
rect -5633 -1339 -5587 -1327
rect -5633 -2315 -5627 -1339
rect -5593 -2315 -5587 -1339
rect -5633 -2327 -5587 -2315
rect -5375 -1339 -5329 -1327
rect -5375 -2315 -5369 -1339
rect -5335 -2315 -5329 -1339
rect -5375 -2327 -5329 -2315
rect -5255 -1339 -5209 -1327
rect -5255 -2315 -5249 -1339
rect -5215 -2315 -5209 -1339
rect -5255 -2327 -5209 -2315
rect -4997 -1339 -4951 -1327
rect -4997 -2315 -4991 -1339
rect -4957 -2315 -4951 -1339
rect -4997 -2327 -4951 -2315
rect -4877 -1339 -4831 -1327
rect -4877 -2315 -4871 -1339
rect -4837 -2315 -4831 -1339
rect -4877 -2327 -4831 -2315
rect -4619 -1339 -4573 -1327
rect -4619 -2315 -4613 -1339
rect -4579 -2315 -4573 -1339
rect -4619 -2327 -4573 -2315
rect -4499 -1339 -4453 -1327
rect -4499 -2315 -4493 -1339
rect -4459 -2315 -4453 -1339
rect -4499 -2327 -4453 -2315
rect -4241 -1339 -4195 -1327
rect -4241 -2315 -4235 -1339
rect -4201 -2315 -4195 -1339
rect -4241 -2327 -4195 -2315
rect -4121 -1339 -4075 -1327
rect -4121 -2315 -4115 -1339
rect -4081 -2315 -4075 -1339
rect -4121 -2327 -4075 -2315
rect -3863 -1339 -3817 -1327
rect -3863 -2315 -3857 -1339
rect -3823 -2315 -3817 -1339
rect -3863 -2327 -3817 -2315
rect -3743 -1339 -3697 -1327
rect -3743 -2315 -3737 -1339
rect -3703 -2315 -3697 -1339
rect -3743 -2327 -3697 -2315
rect -3485 -1339 -3439 -1327
rect -3485 -2315 -3479 -1339
rect -3445 -2315 -3439 -1339
rect -3485 -2327 -3439 -2315
rect -3365 -1339 -3319 -1327
rect -3365 -2315 -3359 -1339
rect -3325 -2315 -3319 -1339
rect -3365 -2327 -3319 -2315
rect -3107 -1339 -3061 -1327
rect -3107 -2315 -3101 -1339
rect -3067 -2315 -3061 -1339
rect -3107 -2327 -3061 -2315
rect -2987 -1339 -2941 -1327
rect -2987 -2315 -2981 -1339
rect -2947 -2315 -2941 -1339
rect -2987 -2327 -2941 -2315
rect -2729 -1339 -2683 -1327
rect -2729 -2315 -2723 -1339
rect -2689 -2315 -2683 -1339
rect -2729 -2327 -2683 -2315
rect -2609 -1339 -2563 -1327
rect -2609 -2315 -2603 -1339
rect -2569 -2315 -2563 -1339
rect -2609 -2327 -2563 -2315
rect -2351 -1339 -2305 -1327
rect -2351 -2315 -2345 -1339
rect -2311 -2315 -2305 -1339
rect -2351 -2327 -2305 -2315
rect -2231 -1339 -2185 -1327
rect -2231 -2315 -2225 -1339
rect -2191 -2315 -2185 -1339
rect -2231 -2327 -2185 -2315
rect -1973 -1339 -1927 -1327
rect -1973 -2315 -1967 -1339
rect -1933 -2315 -1927 -1339
rect -1973 -2327 -1927 -2315
rect -1853 -1339 -1807 -1327
rect -1853 -2315 -1847 -1339
rect -1813 -2315 -1807 -1339
rect -1853 -2327 -1807 -2315
rect -1595 -1339 -1549 -1327
rect -1595 -2315 -1589 -1339
rect -1555 -2315 -1549 -1339
rect -1595 -2327 -1549 -2315
rect -1475 -1339 -1429 -1327
rect -1475 -2315 -1469 -1339
rect -1435 -2315 -1429 -1339
rect -1475 -2327 -1429 -2315
rect -1217 -1339 -1171 -1327
rect -1217 -2315 -1211 -1339
rect -1177 -2315 -1171 -1339
rect -1217 -2327 -1171 -2315
rect -1097 -1339 -1051 -1327
rect -1097 -2315 -1091 -1339
rect -1057 -2315 -1051 -1339
rect -1097 -2327 -1051 -2315
rect -839 -1339 -793 -1327
rect -839 -2315 -833 -1339
rect -799 -2315 -793 -1339
rect -839 -2327 -793 -2315
rect -719 -1339 -673 -1327
rect -719 -2315 -713 -1339
rect -679 -2315 -673 -1339
rect -719 -2327 -673 -2315
rect -461 -1339 -415 -1327
rect -461 -2315 -455 -1339
rect -421 -2315 -415 -1339
rect -461 -2327 -415 -2315
rect -341 -1339 -295 -1327
rect -341 -2315 -335 -1339
rect -301 -2315 -295 -1339
rect -341 -2327 -295 -2315
rect -83 -1339 -37 -1327
rect -83 -2315 -77 -1339
rect -43 -2315 -37 -1339
rect -83 -2327 -37 -2315
rect 37 -1339 83 -1327
rect 37 -2315 43 -1339
rect 77 -2315 83 -1339
rect 37 -2327 83 -2315
rect 295 -1339 341 -1327
rect 295 -2315 301 -1339
rect 335 -2315 341 -1339
rect 295 -2327 341 -2315
rect 415 -1339 461 -1327
rect 415 -2315 421 -1339
rect 455 -2315 461 -1339
rect 415 -2327 461 -2315
rect 673 -1339 719 -1327
rect 673 -2315 679 -1339
rect 713 -2315 719 -1339
rect 673 -2327 719 -2315
rect 793 -1339 839 -1327
rect 793 -2315 799 -1339
rect 833 -2315 839 -1339
rect 793 -2327 839 -2315
rect 1051 -1339 1097 -1327
rect 1051 -2315 1057 -1339
rect 1091 -2315 1097 -1339
rect 1051 -2327 1097 -2315
rect 1171 -1339 1217 -1327
rect 1171 -2315 1177 -1339
rect 1211 -2315 1217 -1339
rect 1171 -2327 1217 -2315
rect 1429 -1339 1475 -1327
rect 1429 -2315 1435 -1339
rect 1469 -2315 1475 -1339
rect 1429 -2327 1475 -2315
rect 1549 -1339 1595 -1327
rect 1549 -2315 1555 -1339
rect 1589 -2315 1595 -1339
rect 1549 -2327 1595 -2315
rect 1807 -1339 1853 -1327
rect 1807 -2315 1813 -1339
rect 1847 -2315 1853 -1339
rect 1807 -2327 1853 -2315
rect 1927 -1339 1973 -1327
rect 1927 -2315 1933 -1339
rect 1967 -2315 1973 -1339
rect 1927 -2327 1973 -2315
rect 2185 -1339 2231 -1327
rect 2185 -2315 2191 -1339
rect 2225 -2315 2231 -1339
rect 2185 -2327 2231 -2315
rect 2305 -1339 2351 -1327
rect 2305 -2315 2311 -1339
rect 2345 -2315 2351 -1339
rect 2305 -2327 2351 -2315
rect 2563 -1339 2609 -1327
rect 2563 -2315 2569 -1339
rect 2603 -2315 2609 -1339
rect 2563 -2327 2609 -2315
rect 2683 -1339 2729 -1327
rect 2683 -2315 2689 -1339
rect 2723 -2315 2729 -1339
rect 2683 -2327 2729 -2315
rect 2941 -1339 2987 -1327
rect 2941 -2315 2947 -1339
rect 2981 -2315 2987 -1339
rect 2941 -2327 2987 -2315
rect 3061 -1339 3107 -1327
rect 3061 -2315 3067 -1339
rect 3101 -2315 3107 -1339
rect 3061 -2327 3107 -2315
rect 3319 -1339 3365 -1327
rect 3319 -2315 3325 -1339
rect 3359 -2315 3365 -1339
rect 3319 -2327 3365 -2315
rect 3439 -1339 3485 -1327
rect 3439 -2315 3445 -1339
rect 3479 -2315 3485 -1339
rect 3439 -2327 3485 -2315
rect 3697 -1339 3743 -1327
rect 3697 -2315 3703 -1339
rect 3737 -2315 3743 -1339
rect 3697 -2327 3743 -2315
rect 3817 -1339 3863 -1327
rect 3817 -2315 3823 -1339
rect 3857 -2315 3863 -1339
rect 3817 -2327 3863 -2315
rect 4075 -1339 4121 -1327
rect 4075 -2315 4081 -1339
rect 4115 -2315 4121 -1339
rect 4075 -2327 4121 -2315
rect 4195 -1339 4241 -1327
rect 4195 -2315 4201 -1339
rect 4235 -2315 4241 -1339
rect 4195 -2327 4241 -2315
rect 4453 -1339 4499 -1327
rect 4453 -2315 4459 -1339
rect 4493 -2315 4499 -1339
rect 4453 -2327 4499 -2315
rect 4573 -1339 4619 -1327
rect 4573 -2315 4579 -1339
rect 4613 -2315 4619 -1339
rect 4573 -2327 4619 -2315
rect 4831 -1339 4877 -1327
rect 4831 -2315 4837 -1339
rect 4871 -2315 4877 -1339
rect 4831 -2327 4877 -2315
rect 4951 -1339 4997 -1327
rect 4951 -2315 4957 -1339
rect 4991 -2315 4997 -1339
rect 4951 -2327 4997 -2315
rect 5209 -1339 5255 -1327
rect 5209 -2315 5215 -1339
rect 5249 -2315 5255 -1339
rect 5209 -2327 5255 -2315
rect 5329 -1339 5375 -1327
rect 5329 -2315 5335 -1339
rect 5369 -2315 5375 -1339
rect 5329 -2327 5375 -2315
rect 5587 -1339 5633 -1327
rect 5587 -2315 5593 -1339
rect 5627 -2315 5633 -1339
rect 5587 -2327 5633 -2315
rect 5707 -1339 5753 -1327
rect 5707 -2315 5713 -1339
rect 5747 -2315 5753 -1339
rect 5707 -2327 5753 -2315
rect 5965 -1339 6011 -1327
rect 5965 -2315 5971 -1339
rect 6005 -2315 6011 -1339
rect 5965 -2327 6011 -2315
rect 6085 -1339 6131 -1327
rect 6085 -2315 6091 -1339
rect 6125 -2315 6131 -1339
rect 6085 -2327 6131 -2315
rect 6343 -1339 6389 -1327
rect 6343 -2315 6349 -1339
rect 6383 -2315 6389 -1339
rect 6343 -2327 6389 -2315
rect 6463 -1339 6509 -1327
rect 6463 -2315 6469 -1339
rect 6503 -2315 6509 -1339
rect 6463 -2327 6509 -2315
rect 6721 -1339 6767 -1327
rect 6721 -2315 6727 -1339
rect 6761 -2315 6767 -1339
rect 6721 -2327 6767 -2315
rect 6841 -1339 6887 -1327
rect 6841 -2315 6847 -1339
rect 6881 -2315 6887 -1339
rect 6841 -2327 6887 -2315
rect 7099 -1339 7145 -1327
rect 7099 -2315 7105 -1339
rect 7139 -2315 7145 -1339
rect 7099 -2327 7145 -2315
rect 7219 -1339 7265 -1327
rect 7219 -2315 7225 -1339
rect 7259 -2315 7265 -1339
rect 7219 -2327 7265 -2315
rect 7477 -1339 7523 -1327
rect 7477 -2315 7483 -1339
rect 7517 -2315 7523 -1339
rect 7477 -2327 7523 -2315
rect 7597 -1339 7643 -1327
rect 7597 -2315 7603 -1339
rect 7637 -2315 7643 -1339
rect 7597 -2327 7643 -2315
rect 7855 -1339 7901 -1327
rect 7855 -2315 7861 -1339
rect 7895 -2315 7901 -1339
rect 7855 -2327 7901 -2315
rect 7975 -1339 8021 -1327
rect 7975 -2315 7981 -1339
rect 8015 -2315 8021 -1339
rect 7975 -2327 8021 -2315
rect 8233 -1339 8279 -1327
rect 8233 -2315 8239 -1339
rect 8273 -2315 8279 -1339
rect 8233 -2327 8279 -2315
rect 8353 -1339 8399 -1327
rect 8353 -2315 8359 -1339
rect 8393 -2315 8399 -1339
rect 8353 -2327 8399 -2315
rect 8611 -1339 8657 -1327
rect 8611 -2315 8617 -1339
rect 8651 -2315 8657 -1339
rect 8611 -2327 8657 -2315
rect 8731 -1339 8777 -1327
rect 8731 -2315 8737 -1339
rect 8771 -2315 8777 -1339
rect 8731 -2327 8777 -2315
rect 8989 -1339 9035 -1327
rect 8989 -2315 8995 -1339
rect 9029 -2315 9035 -1339
rect 8989 -2327 9035 -2315
rect 9109 -1339 9155 -1327
rect 9109 -2315 9115 -1339
rect 9149 -2315 9155 -1339
rect 9109 -2327 9155 -2315
rect 9367 -1339 9413 -1327
rect 9367 -2315 9373 -1339
rect 9407 -2315 9413 -1339
rect 9367 -2327 9413 -2315
rect -9357 -2365 -9165 -2359
rect -9357 -2399 -9345 -2365
rect -9177 -2399 -9165 -2365
rect -9357 -2405 -9165 -2399
rect -8979 -2365 -8787 -2359
rect -8979 -2399 -8967 -2365
rect -8799 -2399 -8787 -2365
rect -8979 -2405 -8787 -2399
rect -8601 -2365 -8409 -2359
rect -8601 -2399 -8589 -2365
rect -8421 -2399 -8409 -2365
rect -8601 -2405 -8409 -2399
rect -8223 -2365 -8031 -2359
rect -8223 -2399 -8211 -2365
rect -8043 -2399 -8031 -2365
rect -8223 -2405 -8031 -2399
rect -7845 -2365 -7653 -2359
rect -7845 -2399 -7833 -2365
rect -7665 -2399 -7653 -2365
rect -7845 -2405 -7653 -2399
rect -7467 -2365 -7275 -2359
rect -7467 -2399 -7455 -2365
rect -7287 -2399 -7275 -2365
rect -7467 -2405 -7275 -2399
rect -7089 -2365 -6897 -2359
rect -7089 -2399 -7077 -2365
rect -6909 -2399 -6897 -2365
rect -7089 -2405 -6897 -2399
rect -6711 -2365 -6519 -2359
rect -6711 -2399 -6699 -2365
rect -6531 -2399 -6519 -2365
rect -6711 -2405 -6519 -2399
rect -6333 -2365 -6141 -2359
rect -6333 -2399 -6321 -2365
rect -6153 -2399 -6141 -2365
rect -6333 -2405 -6141 -2399
rect -5955 -2365 -5763 -2359
rect -5955 -2399 -5943 -2365
rect -5775 -2399 -5763 -2365
rect -5955 -2405 -5763 -2399
rect -5577 -2365 -5385 -2359
rect -5577 -2399 -5565 -2365
rect -5397 -2399 -5385 -2365
rect -5577 -2405 -5385 -2399
rect -5199 -2365 -5007 -2359
rect -5199 -2399 -5187 -2365
rect -5019 -2399 -5007 -2365
rect -5199 -2405 -5007 -2399
rect -4821 -2365 -4629 -2359
rect -4821 -2399 -4809 -2365
rect -4641 -2399 -4629 -2365
rect -4821 -2405 -4629 -2399
rect -4443 -2365 -4251 -2359
rect -4443 -2399 -4431 -2365
rect -4263 -2399 -4251 -2365
rect -4443 -2405 -4251 -2399
rect -4065 -2365 -3873 -2359
rect -4065 -2399 -4053 -2365
rect -3885 -2399 -3873 -2365
rect -4065 -2405 -3873 -2399
rect -3687 -2365 -3495 -2359
rect -3687 -2399 -3675 -2365
rect -3507 -2399 -3495 -2365
rect -3687 -2405 -3495 -2399
rect -3309 -2365 -3117 -2359
rect -3309 -2399 -3297 -2365
rect -3129 -2399 -3117 -2365
rect -3309 -2405 -3117 -2399
rect -2931 -2365 -2739 -2359
rect -2931 -2399 -2919 -2365
rect -2751 -2399 -2739 -2365
rect -2931 -2405 -2739 -2399
rect -2553 -2365 -2361 -2359
rect -2553 -2399 -2541 -2365
rect -2373 -2399 -2361 -2365
rect -2553 -2405 -2361 -2399
rect -2175 -2365 -1983 -2359
rect -2175 -2399 -2163 -2365
rect -1995 -2399 -1983 -2365
rect -2175 -2405 -1983 -2399
rect -1797 -2365 -1605 -2359
rect -1797 -2399 -1785 -2365
rect -1617 -2399 -1605 -2365
rect -1797 -2405 -1605 -2399
rect -1419 -2365 -1227 -2359
rect -1419 -2399 -1407 -2365
rect -1239 -2399 -1227 -2365
rect -1419 -2405 -1227 -2399
rect -1041 -2365 -849 -2359
rect -1041 -2399 -1029 -2365
rect -861 -2399 -849 -2365
rect -1041 -2405 -849 -2399
rect -663 -2365 -471 -2359
rect -663 -2399 -651 -2365
rect -483 -2399 -471 -2365
rect -663 -2405 -471 -2399
rect -285 -2365 -93 -2359
rect -285 -2399 -273 -2365
rect -105 -2399 -93 -2365
rect -285 -2405 -93 -2399
rect 93 -2365 285 -2359
rect 93 -2399 105 -2365
rect 273 -2399 285 -2365
rect 93 -2405 285 -2399
rect 471 -2365 663 -2359
rect 471 -2399 483 -2365
rect 651 -2399 663 -2365
rect 471 -2405 663 -2399
rect 849 -2365 1041 -2359
rect 849 -2399 861 -2365
rect 1029 -2399 1041 -2365
rect 849 -2405 1041 -2399
rect 1227 -2365 1419 -2359
rect 1227 -2399 1239 -2365
rect 1407 -2399 1419 -2365
rect 1227 -2405 1419 -2399
rect 1605 -2365 1797 -2359
rect 1605 -2399 1617 -2365
rect 1785 -2399 1797 -2365
rect 1605 -2405 1797 -2399
rect 1983 -2365 2175 -2359
rect 1983 -2399 1995 -2365
rect 2163 -2399 2175 -2365
rect 1983 -2405 2175 -2399
rect 2361 -2365 2553 -2359
rect 2361 -2399 2373 -2365
rect 2541 -2399 2553 -2365
rect 2361 -2405 2553 -2399
rect 2739 -2365 2931 -2359
rect 2739 -2399 2751 -2365
rect 2919 -2399 2931 -2365
rect 2739 -2405 2931 -2399
rect 3117 -2365 3309 -2359
rect 3117 -2399 3129 -2365
rect 3297 -2399 3309 -2365
rect 3117 -2405 3309 -2399
rect 3495 -2365 3687 -2359
rect 3495 -2399 3507 -2365
rect 3675 -2399 3687 -2365
rect 3495 -2405 3687 -2399
rect 3873 -2365 4065 -2359
rect 3873 -2399 3885 -2365
rect 4053 -2399 4065 -2365
rect 3873 -2405 4065 -2399
rect 4251 -2365 4443 -2359
rect 4251 -2399 4263 -2365
rect 4431 -2399 4443 -2365
rect 4251 -2405 4443 -2399
rect 4629 -2365 4821 -2359
rect 4629 -2399 4641 -2365
rect 4809 -2399 4821 -2365
rect 4629 -2405 4821 -2399
rect 5007 -2365 5199 -2359
rect 5007 -2399 5019 -2365
rect 5187 -2399 5199 -2365
rect 5007 -2405 5199 -2399
rect 5385 -2365 5577 -2359
rect 5385 -2399 5397 -2365
rect 5565 -2399 5577 -2365
rect 5385 -2405 5577 -2399
rect 5763 -2365 5955 -2359
rect 5763 -2399 5775 -2365
rect 5943 -2399 5955 -2365
rect 5763 -2405 5955 -2399
rect 6141 -2365 6333 -2359
rect 6141 -2399 6153 -2365
rect 6321 -2399 6333 -2365
rect 6141 -2405 6333 -2399
rect 6519 -2365 6711 -2359
rect 6519 -2399 6531 -2365
rect 6699 -2399 6711 -2365
rect 6519 -2405 6711 -2399
rect 6897 -2365 7089 -2359
rect 6897 -2399 6909 -2365
rect 7077 -2399 7089 -2365
rect 6897 -2405 7089 -2399
rect 7275 -2365 7467 -2359
rect 7275 -2399 7287 -2365
rect 7455 -2399 7467 -2365
rect 7275 -2405 7467 -2399
rect 7653 -2365 7845 -2359
rect 7653 -2399 7665 -2365
rect 7833 -2399 7845 -2365
rect 7653 -2405 7845 -2399
rect 8031 -2365 8223 -2359
rect 8031 -2399 8043 -2365
rect 8211 -2399 8223 -2365
rect 8031 -2405 8223 -2399
rect 8409 -2365 8601 -2359
rect 8409 -2399 8421 -2365
rect 8589 -2399 8601 -2365
rect 8409 -2405 8601 -2399
rect 8787 -2365 8979 -2359
rect 8787 -2399 8799 -2365
rect 8967 -2399 8979 -2365
rect 8787 -2405 8979 -2399
rect 9165 -2365 9357 -2359
rect 9165 -2399 9177 -2365
rect 9345 -2399 9357 -2365
rect 9165 -2405 9357 -2399
<< properties >>
string FIXED_BBOX -9524 -2520 9524 2520
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 1.0 m 4 nf 50 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
