magic
tech sky130A
magscale 1 2
timestamp 1730737834
<< pwell >>
rect -7294 -2423 7294 2423
<< mvnmos >>
rect -7066 1165 -6866 2165
rect -6808 1165 -6608 2165
rect -6550 1165 -6350 2165
rect -6292 1165 -6092 2165
rect -6034 1165 -5834 2165
rect -5776 1165 -5576 2165
rect -5518 1165 -5318 2165
rect -5260 1165 -5060 2165
rect -5002 1165 -4802 2165
rect -4744 1165 -4544 2165
rect -4486 1165 -4286 2165
rect -4228 1165 -4028 2165
rect -3970 1165 -3770 2165
rect -3712 1165 -3512 2165
rect -3454 1165 -3254 2165
rect -3196 1165 -2996 2165
rect -2938 1165 -2738 2165
rect -2680 1165 -2480 2165
rect -2422 1165 -2222 2165
rect -2164 1165 -1964 2165
rect -1906 1165 -1706 2165
rect -1648 1165 -1448 2165
rect -1390 1165 -1190 2165
rect -1132 1165 -932 2165
rect -874 1165 -674 2165
rect -616 1165 -416 2165
rect -358 1165 -158 2165
rect -100 1165 100 2165
rect 158 1165 358 2165
rect 416 1165 616 2165
rect 674 1165 874 2165
rect 932 1165 1132 2165
rect 1190 1165 1390 2165
rect 1448 1165 1648 2165
rect 1706 1165 1906 2165
rect 1964 1165 2164 2165
rect 2222 1165 2422 2165
rect 2480 1165 2680 2165
rect 2738 1165 2938 2165
rect 2996 1165 3196 2165
rect 3254 1165 3454 2165
rect 3512 1165 3712 2165
rect 3770 1165 3970 2165
rect 4028 1165 4228 2165
rect 4286 1165 4486 2165
rect 4544 1165 4744 2165
rect 4802 1165 5002 2165
rect 5060 1165 5260 2165
rect 5318 1165 5518 2165
rect 5576 1165 5776 2165
rect 5834 1165 6034 2165
rect 6092 1165 6292 2165
rect 6350 1165 6550 2165
rect 6608 1165 6808 2165
rect 6866 1165 7066 2165
rect -7066 55 -6866 1055
rect -6808 55 -6608 1055
rect -6550 55 -6350 1055
rect -6292 55 -6092 1055
rect -6034 55 -5834 1055
rect -5776 55 -5576 1055
rect -5518 55 -5318 1055
rect -5260 55 -5060 1055
rect -5002 55 -4802 1055
rect -4744 55 -4544 1055
rect -4486 55 -4286 1055
rect -4228 55 -4028 1055
rect -3970 55 -3770 1055
rect -3712 55 -3512 1055
rect -3454 55 -3254 1055
rect -3196 55 -2996 1055
rect -2938 55 -2738 1055
rect -2680 55 -2480 1055
rect -2422 55 -2222 1055
rect -2164 55 -1964 1055
rect -1906 55 -1706 1055
rect -1648 55 -1448 1055
rect -1390 55 -1190 1055
rect -1132 55 -932 1055
rect -874 55 -674 1055
rect -616 55 -416 1055
rect -358 55 -158 1055
rect -100 55 100 1055
rect 158 55 358 1055
rect 416 55 616 1055
rect 674 55 874 1055
rect 932 55 1132 1055
rect 1190 55 1390 1055
rect 1448 55 1648 1055
rect 1706 55 1906 1055
rect 1964 55 2164 1055
rect 2222 55 2422 1055
rect 2480 55 2680 1055
rect 2738 55 2938 1055
rect 2996 55 3196 1055
rect 3254 55 3454 1055
rect 3512 55 3712 1055
rect 3770 55 3970 1055
rect 4028 55 4228 1055
rect 4286 55 4486 1055
rect 4544 55 4744 1055
rect 4802 55 5002 1055
rect 5060 55 5260 1055
rect 5318 55 5518 1055
rect 5576 55 5776 1055
rect 5834 55 6034 1055
rect 6092 55 6292 1055
rect 6350 55 6550 1055
rect 6608 55 6808 1055
rect 6866 55 7066 1055
rect -7066 -1055 -6866 -55
rect -6808 -1055 -6608 -55
rect -6550 -1055 -6350 -55
rect -6292 -1055 -6092 -55
rect -6034 -1055 -5834 -55
rect -5776 -1055 -5576 -55
rect -5518 -1055 -5318 -55
rect -5260 -1055 -5060 -55
rect -5002 -1055 -4802 -55
rect -4744 -1055 -4544 -55
rect -4486 -1055 -4286 -55
rect -4228 -1055 -4028 -55
rect -3970 -1055 -3770 -55
rect -3712 -1055 -3512 -55
rect -3454 -1055 -3254 -55
rect -3196 -1055 -2996 -55
rect -2938 -1055 -2738 -55
rect -2680 -1055 -2480 -55
rect -2422 -1055 -2222 -55
rect -2164 -1055 -1964 -55
rect -1906 -1055 -1706 -55
rect -1648 -1055 -1448 -55
rect -1390 -1055 -1190 -55
rect -1132 -1055 -932 -55
rect -874 -1055 -674 -55
rect -616 -1055 -416 -55
rect -358 -1055 -158 -55
rect -100 -1055 100 -55
rect 158 -1055 358 -55
rect 416 -1055 616 -55
rect 674 -1055 874 -55
rect 932 -1055 1132 -55
rect 1190 -1055 1390 -55
rect 1448 -1055 1648 -55
rect 1706 -1055 1906 -55
rect 1964 -1055 2164 -55
rect 2222 -1055 2422 -55
rect 2480 -1055 2680 -55
rect 2738 -1055 2938 -55
rect 2996 -1055 3196 -55
rect 3254 -1055 3454 -55
rect 3512 -1055 3712 -55
rect 3770 -1055 3970 -55
rect 4028 -1055 4228 -55
rect 4286 -1055 4486 -55
rect 4544 -1055 4744 -55
rect 4802 -1055 5002 -55
rect 5060 -1055 5260 -55
rect 5318 -1055 5518 -55
rect 5576 -1055 5776 -55
rect 5834 -1055 6034 -55
rect 6092 -1055 6292 -55
rect 6350 -1055 6550 -55
rect 6608 -1055 6808 -55
rect 6866 -1055 7066 -55
rect -7066 -2165 -6866 -1165
rect -6808 -2165 -6608 -1165
rect -6550 -2165 -6350 -1165
rect -6292 -2165 -6092 -1165
rect -6034 -2165 -5834 -1165
rect -5776 -2165 -5576 -1165
rect -5518 -2165 -5318 -1165
rect -5260 -2165 -5060 -1165
rect -5002 -2165 -4802 -1165
rect -4744 -2165 -4544 -1165
rect -4486 -2165 -4286 -1165
rect -4228 -2165 -4028 -1165
rect -3970 -2165 -3770 -1165
rect -3712 -2165 -3512 -1165
rect -3454 -2165 -3254 -1165
rect -3196 -2165 -2996 -1165
rect -2938 -2165 -2738 -1165
rect -2680 -2165 -2480 -1165
rect -2422 -2165 -2222 -1165
rect -2164 -2165 -1964 -1165
rect -1906 -2165 -1706 -1165
rect -1648 -2165 -1448 -1165
rect -1390 -2165 -1190 -1165
rect -1132 -2165 -932 -1165
rect -874 -2165 -674 -1165
rect -616 -2165 -416 -1165
rect -358 -2165 -158 -1165
rect -100 -2165 100 -1165
rect 158 -2165 358 -1165
rect 416 -2165 616 -1165
rect 674 -2165 874 -1165
rect 932 -2165 1132 -1165
rect 1190 -2165 1390 -1165
rect 1448 -2165 1648 -1165
rect 1706 -2165 1906 -1165
rect 1964 -2165 2164 -1165
rect 2222 -2165 2422 -1165
rect 2480 -2165 2680 -1165
rect 2738 -2165 2938 -1165
rect 2996 -2165 3196 -1165
rect 3254 -2165 3454 -1165
rect 3512 -2165 3712 -1165
rect 3770 -2165 3970 -1165
rect 4028 -2165 4228 -1165
rect 4286 -2165 4486 -1165
rect 4544 -2165 4744 -1165
rect 4802 -2165 5002 -1165
rect 5060 -2165 5260 -1165
rect 5318 -2165 5518 -1165
rect 5576 -2165 5776 -1165
rect 5834 -2165 6034 -1165
rect 6092 -2165 6292 -1165
rect 6350 -2165 6550 -1165
rect 6608 -2165 6808 -1165
rect 6866 -2165 7066 -1165
<< mvndiff >>
rect -7124 2153 -7066 2165
rect -7124 1177 -7112 2153
rect -7078 1177 -7066 2153
rect -7124 1165 -7066 1177
rect -6866 2153 -6808 2165
rect -6866 1177 -6854 2153
rect -6820 1177 -6808 2153
rect -6866 1165 -6808 1177
rect -6608 2153 -6550 2165
rect -6608 1177 -6596 2153
rect -6562 1177 -6550 2153
rect -6608 1165 -6550 1177
rect -6350 2153 -6292 2165
rect -6350 1177 -6338 2153
rect -6304 1177 -6292 2153
rect -6350 1165 -6292 1177
rect -6092 2153 -6034 2165
rect -6092 1177 -6080 2153
rect -6046 1177 -6034 2153
rect -6092 1165 -6034 1177
rect -5834 2153 -5776 2165
rect -5834 1177 -5822 2153
rect -5788 1177 -5776 2153
rect -5834 1165 -5776 1177
rect -5576 2153 -5518 2165
rect -5576 1177 -5564 2153
rect -5530 1177 -5518 2153
rect -5576 1165 -5518 1177
rect -5318 2153 -5260 2165
rect -5318 1177 -5306 2153
rect -5272 1177 -5260 2153
rect -5318 1165 -5260 1177
rect -5060 2153 -5002 2165
rect -5060 1177 -5048 2153
rect -5014 1177 -5002 2153
rect -5060 1165 -5002 1177
rect -4802 2153 -4744 2165
rect -4802 1177 -4790 2153
rect -4756 1177 -4744 2153
rect -4802 1165 -4744 1177
rect -4544 2153 -4486 2165
rect -4544 1177 -4532 2153
rect -4498 1177 -4486 2153
rect -4544 1165 -4486 1177
rect -4286 2153 -4228 2165
rect -4286 1177 -4274 2153
rect -4240 1177 -4228 2153
rect -4286 1165 -4228 1177
rect -4028 2153 -3970 2165
rect -4028 1177 -4016 2153
rect -3982 1177 -3970 2153
rect -4028 1165 -3970 1177
rect -3770 2153 -3712 2165
rect -3770 1177 -3758 2153
rect -3724 1177 -3712 2153
rect -3770 1165 -3712 1177
rect -3512 2153 -3454 2165
rect -3512 1177 -3500 2153
rect -3466 1177 -3454 2153
rect -3512 1165 -3454 1177
rect -3254 2153 -3196 2165
rect -3254 1177 -3242 2153
rect -3208 1177 -3196 2153
rect -3254 1165 -3196 1177
rect -2996 2153 -2938 2165
rect -2996 1177 -2984 2153
rect -2950 1177 -2938 2153
rect -2996 1165 -2938 1177
rect -2738 2153 -2680 2165
rect -2738 1177 -2726 2153
rect -2692 1177 -2680 2153
rect -2738 1165 -2680 1177
rect -2480 2153 -2422 2165
rect -2480 1177 -2468 2153
rect -2434 1177 -2422 2153
rect -2480 1165 -2422 1177
rect -2222 2153 -2164 2165
rect -2222 1177 -2210 2153
rect -2176 1177 -2164 2153
rect -2222 1165 -2164 1177
rect -1964 2153 -1906 2165
rect -1964 1177 -1952 2153
rect -1918 1177 -1906 2153
rect -1964 1165 -1906 1177
rect -1706 2153 -1648 2165
rect -1706 1177 -1694 2153
rect -1660 1177 -1648 2153
rect -1706 1165 -1648 1177
rect -1448 2153 -1390 2165
rect -1448 1177 -1436 2153
rect -1402 1177 -1390 2153
rect -1448 1165 -1390 1177
rect -1190 2153 -1132 2165
rect -1190 1177 -1178 2153
rect -1144 1177 -1132 2153
rect -1190 1165 -1132 1177
rect -932 2153 -874 2165
rect -932 1177 -920 2153
rect -886 1177 -874 2153
rect -932 1165 -874 1177
rect -674 2153 -616 2165
rect -674 1177 -662 2153
rect -628 1177 -616 2153
rect -674 1165 -616 1177
rect -416 2153 -358 2165
rect -416 1177 -404 2153
rect -370 1177 -358 2153
rect -416 1165 -358 1177
rect -158 2153 -100 2165
rect -158 1177 -146 2153
rect -112 1177 -100 2153
rect -158 1165 -100 1177
rect 100 2153 158 2165
rect 100 1177 112 2153
rect 146 1177 158 2153
rect 100 1165 158 1177
rect 358 2153 416 2165
rect 358 1177 370 2153
rect 404 1177 416 2153
rect 358 1165 416 1177
rect 616 2153 674 2165
rect 616 1177 628 2153
rect 662 1177 674 2153
rect 616 1165 674 1177
rect 874 2153 932 2165
rect 874 1177 886 2153
rect 920 1177 932 2153
rect 874 1165 932 1177
rect 1132 2153 1190 2165
rect 1132 1177 1144 2153
rect 1178 1177 1190 2153
rect 1132 1165 1190 1177
rect 1390 2153 1448 2165
rect 1390 1177 1402 2153
rect 1436 1177 1448 2153
rect 1390 1165 1448 1177
rect 1648 2153 1706 2165
rect 1648 1177 1660 2153
rect 1694 1177 1706 2153
rect 1648 1165 1706 1177
rect 1906 2153 1964 2165
rect 1906 1177 1918 2153
rect 1952 1177 1964 2153
rect 1906 1165 1964 1177
rect 2164 2153 2222 2165
rect 2164 1177 2176 2153
rect 2210 1177 2222 2153
rect 2164 1165 2222 1177
rect 2422 2153 2480 2165
rect 2422 1177 2434 2153
rect 2468 1177 2480 2153
rect 2422 1165 2480 1177
rect 2680 2153 2738 2165
rect 2680 1177 2692 2153
rect 2726 1177 2738 2153
rect 2680 1165 2738 1177
rect 2938 2153 2996 2165
rect 2938 1177 2950 2153
rect 2984 1177 2996 2153
rect 2938 1165 2996 1177
rect 3196 2153 3254 2165
rect 3196 1177 3208 2153
rect 3242 1177 3254 2153
rect 3196 1165 3254 1177
rect 3454 2153 3512 2165
rect 3454 1177 3466 2153
rect 3500 1177 3512 2153
rect 3454 1165 3512 1177
rect 3712 2153 3770 2165
rect 3712 1177 3724 2153
rect 3758 1177 3770 2153
rect 3712 1165 3770 1177
rect 3970 2153 4028 2165
rect 3970 1177 3982 2153
rect 4016 1177 4028 2153
rect 3970 1165 4028 1177
rect 4228 2153 4286 2165
rect 4228 1177 4240 2153
rect 4274 1177 4286 2153
rect 4228 1165 4286 1177
rect 4486 2153 4544 2165
rect 4486 1177 4498 2153
rect 4532 1177 4544 2153
rect 4486 1165 4544 1177
rect 4744 2153 4802 2165
rect 4744 1177 4756 2153
rect 4790 1177 4802 2153
rect 4744 1165 4802 1177
rect 5002 2153 5060 2165
rect 5002 1177 5014 2153
rect 5048 1177 5060 2153
rect 5002 1165 5060 1177
rect 5260 2153 5318 2165
rect 5260 1177 5272 2153
rect 5306 1177 5318 2153
rect 5260 1165 5318 1177
rect 5518 2153 5576 2165
rect 5518 1177 5530 2153
rect 5564 1177 5576 2153
rect 5518 1165 5576 1177
rect 5776 2153 5834 2165
rect 5776 1177 5788 2153
rect 5822 1177 5834 2153
rect 5776 1165 5834 1177
rect 6034 2153 6092 2165
rect 6034 1177 6046 2153
rect 6080 1177 6092 2153
rect 6034 1165 6092 1177
rect 6292 2153 6350 2165
rect 6292 1177 6304 2153
rect 6338 1177 6350 2153
rect 6292 1165 6350 1177
rect 6550 2153 6608 2165
rect 6550 1177 6562 2153
rect 6596 1177 6608 2153
rect 6550 1165 6608 1177
rect 6808 2153 6866 2165
rect 6808 1177 6820 2153
rect 6854 1177 6866 2153
rect 6808 1165 6866 1177
rect 7066 2153 7124 2165
rect 7066 1177 7078 2153
rect 7112 1177 7124 2153
rect 7066 1165 7124 1177
rect -7124 1043 -7066 1055
rect -7124 67 -7112 1043
rect -7078 67 -7066 1043
rect -7124 55 -7066 67
rect -6866 1043 -6808 1055
rect -6866 67 -6854 1043
rect -6820 67 -6808 1043
rect -6866 55 -6808 67
rect -6608 1043 -6550 1055
rect -6608 67 -6596 1043
rect -6562 67 -6550 1043
rect -6608 55 -6550 67
rect -6350 1043 -6292 1055
rect -6350 67 -6338 1043
rect -6304 67 -6292 1043
rect -6350 55 -6292 67
rect -6092 1043 -6034 1055
rect -6092 67 -6080 1043
rect -6046 67 -6034 1043
rect -6092 55 -6034 67
rect -5834 1043 -5776 1055
rect -5834 67 -5822 1043
rect -5788 67 -5776 1043
rect -5834 55 -5776 67
rect -5576 1043 -5518 1055
rect -5576 67 -5564 1043
rect -5530 67 -5518 1043
rect -5576 55 -5518 67
rect -5318 1043 -5260 1055
rect -5318 67 -5306 1043
rect -5272 67 -5260 1043
rect -5318 55 -5260 67
rect -5060 1043 -5002 1055
rect -5060 67 -5048 1043
rect -5014 67 -5002 1043
rect -5060 55 -5002 67
rect -4802 1043 -4744 1055
rect -4802 67 -4790 1043
rect -4756 67 -4744 1043
rect -4802 55 -4744 67
rect -4544 1043 -4486 1055
rect -4544 67 -4532 1043
rect -4498 67 -4486 1043
rect -4544 55 -4486 67
rect -4286 1043 -4228 1055
rect -4286 67 -4274 1043
rect -4240 67 -4228 1043
rect -4286 55 -4228 67
rect -4028 1043 -3970 1055
rect -4028 67 -4016 1043
rect -3982 67 -3970 1043
rect -4028 55 -3970 67
rect -3770 1043 -3712 1055
rect -3770 67 -3758 1043
rect -3724 67 -3712 1043
rect -3770 55 -3712 67
rect -3512 1043 -3454 1055
rect -3512 67 -3500 1043
rect -3466 67 -3454 1043
rect -3512 55 -3454 67
rect -3254 1043 -3196 1055
rect -3254 67 -3242 1043
rect -3208 67 -3196 1043
rect -3254 55 -3196 67
rect -2996 1043 -2938 1055
rect -2996 67 -2984 1043
rect -2950 67 -2938 1043
rect -2996 55 -2938 67
rect -2738 1043 -2680 1055
rect -2738 67 -2726 1043
rect -2692 67 -2680 1043
rect -2738 55 -2680 67
rect -2480 1043 -2422 1055
rect -2480 67 -2468 1043
rect -2434 67 -2422 1043
rect -2480 55 -2422 67
rect -2222 1043 -2164 1055
rect -2222 67 -2210 1043
rect -2176 67 -2164 1043
rect -2222 55 -2164 67
rect -1964 1043 -1906 1055
rect -1964 67 -1952 1043
rect -1918 67 -1906 1043
rect -1964 55 -1906 67
rect -1706 1043 -1648 1055
rect -1706 67 -1694 1043
rect -1660 67 -1648 1043
rect -1706 55 -1648 67
rect -1448 1043 -1390 1055
rect -1448 67 -1436 1043
rect -1402 67 -1390 1043
rect -1448 55 -1390 67
rect -1190 1043 -1132 1055
rect -1190 67 -1178 1043
rect -1144 67 -1132 1043
rect -1190 55 -1132 67
rect -932 1043 -874 1055
rect -932 67 -920 1043
rect -886 67 -874 1043
rect -932 55 -874 67
rect -674 1043 -616 1055
rect -674 67 -662 1043
rect -628 67 -616 1043
rect -674 55 -616 67
rect -416 1043 -358 1055
rect -416 67 -404 1043
rect -370 67 -358 1043
rect -416 55 -358 67
rect -158 1043 -100 1055
rect -158 67 -146 1043
rect -112 67 -100 1043
rect -158 55 -100 67
rect 100 1043 158 1055
rect 100 67 112 1043
rect 146 67 158 1043
rect 100 55 158 67
rect 358 1043 416 1055
rect 358 67 370 1043
rect 404 67 416 1043
rect 358 55 416 67
rect 616 1043 674 1055
rect 616 67 628 1043
rect 662 67 674 1043
rect 616 55 674 67
rect 874 1043 932 1055
rect 874 67 886 1043
rect 920 67 932 1043
rect 874 55 932 67
rect 1132 1043 1190 1055
rect 1132 67 1144 1043
rect 1178 67 1190 1043
rect 1132 55 1190 67
rect 1390 1043 1448 1055
rect 1390 67 1402 1043
rect 1436 67 1448 1043
rect 1390 55 1448 67
rect 1648 1043 1706 1055
rect 1648 67 1660 1043
rect 1694 67 1706 1043
rect 1648 55 1706 67
rect 1906 1043 1964 1055
rect 1906 67 1918 1043
rect 1952 67 1964 1043
rect 1906 55 1964 67
rect 2164 1043 2222 1055
rect 2164 67 2176 1043
rect 2210 67 2222 1043
rect 2164 55 2222 67
rect 2422 1043 2480 1055
rect 2422 67 2434 1043
rect 2468 67 2480 1043
rect 2422 55 2480 67
rect 2680 1043 2738 1055
rect 2680 67 2692 1043
rect 2726 67 2738 1043
rect 2680 55 2738 67
rect 2938 1043 2996 1055
rect 2938 67 2950 1043
rect 2984 67 2996 1043
rect 2938 55 2996 67
rect 3196 1043 3254 1055
rect 3196 67 3208 1043
rect 3242 67 3254 1043
rect 3196 55 3254 67
rect 3454 1043 3512 1055
rect 3454 67 3466 1043
rect 3500 67 3512 1043
rect 3454 55 3512 67
rect 3712 1043 3770 1055
rect 3712 67 3724 1043
rect 3758 67 3770 1043
rect 3712 55 3770 67
rect 3970 1043 4028 1055
rect 3970 67 3982 1043
rect 4016 67 4028 1043
rect 3970 55 4028 67
rect 4228 1043 4286 1055
rect 4228 67 4240 1043
rect 4274 67 4286 1043
rect 4228 55 4286 67
rect 4486 1043 4544 1055
rect 4486 67 4498 1043
rect 4532 67 4544 1043
rect 4486 55 4544 67
rect 4744 1043 4802 1055
rect 4744 67 4756 1043
rect 4790 67 4802 1043
rect 4744 55 4802 67
rect 5002 1043 5060 1055
rect 5002 67 5014 1043
rect 5048 67 5060 1043
rect 5002 55 5060 67
rect 5260 1043 5318 1055
rect 5260 67 5272 1043
rect 5306 67 5318 1043
rect 5260 55 5318 67
rect 5518 1043 5576 1055
rect 5518 67 5530 1043
rect 5564 67 5576 1043
rect 5518 55 5576 67
rect 5776 1043 5834 1055
rect 5776 67 5788 1043
rect 5822 67 5834 1043
rect 5776 55 5834 67
rect 6034 1043 6092 1055
rect 6034 67 6046 1043
rect 6080 67 6092 1043
rect 6034 55 6092 67
rect 6292 1043 6350 1055
rect 6292 67 6304 1043
rect 6338 67 6350 1043
rect 6292 55 6350 67
rect 6550 1043 6608 1055
rect 6550 67 6562 1043
rect 6596 67 6608 1043
rect 6550 55 6608 67
rect 6808 1043 6866 1055
rect 6808 67 6820 1043
rect 6854 67 6866 1043
rect 6808 55 6866 67
rect 7066 1043 7124 1055
rect 7066 67 7078 1043
rect 7112 67 7124 1043
rect 7066 55 7124 67
rect -7124 -67 -7066 -55
rect -7124 -1043 -7112 -67
rect -7078 -1043 -7066 -67
rect -7124 -1055 -7066 -1043
rect -6866 -67 -6808 -55
rect -6866 -1043 -6854 -67
rect -6820 -1043 -6808 -67
rect -6866 -1055 -6808 -1043
rect -6608 -67 -6550 -55
rect -6608 -1043 -6596 -67
rect -6562 -1043 -6550 -67
rect -6608 -1055 -6550 -1043
rect -6350 -67 -6292 -55
rect -6350 -1043 -6338 -67
rect -6304 -1043 -6292 -67
rect -6350 -1055 -6292 -1043
rect -6092 -67 -6034 -55
rect -6092 -1043 -6080 -67
rect -6046 -1043 -6034 -67
rect -6092 -1055 -6034 -1043
rect -5834 -67 -5776 -55
rect -5834 -1043 -5822 -67
rect -5788 -1043 -5776 -67
rect -5834 -1055 -5776 -1043
rect -5576 -67 -5518 -55
rect -5576 -1043 -5564 -67
rect -5530 -1043 -5518 -67
rect -5576 -1055 -5518 -1043
rect -5318 -67 -5260 -55
rect -5318 -1043 -5306 -67
rect -5272 -1043 -5260 -67
rect -5318 -1055 -5260 -1043
rect -5060 -67 -5002 -55
rect -5060 -1043 -5048 -67
rect -5014 -1043 -5002 -67
rect -5060 -1055 -5002 -1043
rect -4802 -67 -4744 -55
rect -4802 -1043 -4790 -67
rect -4756 -1043 -4744 -67
rect -4802 -1055 -4744 -1043
rect -4544 -67 -4486 -55
rect -4544 -1043 -4532 -67
rect -4498 -1043 -4486 -67
rect -4544 -1055 -4486 -1043
rect -4286 -67 -4228 -55
rect -4286 -1043 -4274 -67
rect -4240 -1043 -4228 -67
rect -4286 -1055 -4228 -1043
rect -4028 -67 -3970 -55
rect -4028 -1043 -4016 -67
rect -3982 -1043 -3970 -67
rect -4028 -1055 -3970 -1043
rect -3770 -67 -3712 -55
rect -3770 -1043 -3758 -67
rect -3724 -1043 -3712 -67
rect -3770 -1055 -3712 -1043
rect -3512 -67 -3454 -55
rect -3512 -1043 -3500 -67
rect -3466 -1043 -3454 -67
rect -3512 -1055 -3454 -1043
rect -3254 -67 -3196 -55
rect -3254 -1043 -3242 -67
rect -3208 -1043 -3196 -67
rect -3254 -1055 -3196 -1043
rect -2996 -67 -2938 -55
rect -2996 -1043 -2984 -67
rect -2950 -1043 -2938 -67
rect -2996 -1055 -2938 -1043
rect -2738 -67 -2680 -55
rect -2738 -1043 -2726 -67
rect -2692 -1043 -2680 -67
rect -2738 -1055 -2680 -1043
rect -2480 -67 -2422 -55
rect -2480 -1043 -2468 -67
rect -2434 -1043 -2422 -67
rect -2480 -1055 -2422 -1043
rect -2222 -67 -2164 -55
rect -2222 -1043 -2210 -67
rect -2176 -1043 -2164 -67
rect -2222 -1055 -2164 -1043
rect -1964 -67 -1906 -55
rect -1964 -1043 -1952 -67
rect -1918 -1043 -1906 -67
rect -1964 -1055 -1906 -1043
rect -1706 -67 -1648 -55
rect -1706 -1043 -1694 -67
rect -1660 -1043 -1648 -67
rect -1706 -1055 -1648 -1043
rect -1448 -67 -1390 -55
rect -1448 -1043 -1436 -67
rect -1402 -1043 -1390 -67
rect -1448 -1055 -1390 -1043
rect -1190 -67 -1132 -55
rect -1190 -1043 -1178 -67
rect -1144 -1043 -1132 -67
rect -1190 -1055 -1132 -1043
rect -932 -67 -874 -55
rect -932 -1043 -920 -67
rect -886 -1043 -874 -67
rect -932 -1055 -874 -1043
rect -674 -67 -616 -55
rect -674 -1043 -662 -67
rect -628 -1043 -616 -67
rect -674 -1055 -616 -1043
rect -416 -67 -358 -55
rect -416 -1043 -404 -67
rect -370 -1043 -358 -67
rect -416 -1055 -358 -1043
rect -158 -67 -100 -55
rect -158 -1043 -146 -67
rect -112 -1043 -100 -67
rect -158 -1055 -100 -1043
rect 100 -67 158 -55
rect 100 -1043 112 -67
rect 146 -1043 158 -67
rect 100 -1055 158 -1043
rect 358 -67 416 -55
rect 358 -1043 370 -67
rect 404 -1043 416 -67
rect 358 -1055 416 -1043
rect 616 -67 674 -55
rect 616 -1043 628 -67
rect 662 -1043 674 -67
rect 616 -1055 674 -1043
rect 874 -67 932 -55
rect 874 -1043 886 -67
rect 920 -1043 932 -67
rect 874 -1055 932 -1043
rect 1132 -67 1190 -55
rect 1132 -1043 1144 -67
rect 1178 -1043 1190 -67
rect 1132 -1055 1190 -1043
rect 1390 -67 1448 -55
rect 1390 -1043 1402 -67
rect 1436 -1043 1448 -67
rect 1390 -1055 1448 -1043
rect 1648 -67 1706 -55
rect 1648 -1043 1660 -67
rect 1694 -1043 1706 -67
rect 1648 -1055 1706 -1043
rect 1906 -67 1964 -55
rect 1906 -1043 1918 -67
rect 1952 -1043 1964 -67
rect 1906 -1055 1964 -1043
rect 2164 -67 2222 -55
rect 2164 -1043 2176 -67
rect 2210 -1043 2222 -67
rect 2164 -1055 2222 -1043
rect 2422 -67 2480 -55
rect 2422 -1043 2434 -67
rect 2468 -1043 2480 -67
rect 2422 -1055 2480 -1043
rect 2680 -67 2738 -55
rect 2680 -1043 2692 -67
rect 2726 -1043 2738 -67
rect 2680 -1055 2738 -1043
rect 2938 -67 2996 -55
rect 2938 -1043 2950 -67
rect 2984 -1043 2996 -67
rect 2938 -1055 2996 -1043
rect 3196 -67 3254 -55
rect 3196 -1043 3208 -67
rect 3242 -1043 3254 -67
rect 3196 -1055 3254 -1043
rect 3454 -67 3512 -55
rect 3454 -1043 3466 -67
rect 3500 -1043 3512 -67
rect 3454 -1055 3512 -1043
rect 3712 -67 3770 -55
rect 3712 -1043 3724 -67
rect 3758 -1043 3770 -67
rect 3712 -1055 3770 -1043
rect 3970 -67 4028 -55
rect 3970 -1043 3982 -67
rect 4016 -1043 4028 -67
rect 3970 -1055 4028 -1043
rect 4228 -67 4286 -55
rect 4228 -1043 4240 -67
rect 4274 -1043 4286 -67
rect 4228 -1055 4286 -1043
rect 4486 -67 4544 -55
rect 4486 -1043 4498 -67
rect 4532 -1043 4544 -67
rect 4486 -1055 4544 -1043
rect 4744 -67 4802 -55
rect 4744 -1043 4756 -67
rect 4790 -1043 4802 -67
rect 4744 -1055 4802 -1043
rect 5002 -67 5060 -55
rect 5002 -1043 5014 -67
rect 5048 -1043 5060 -67
rect 5002 -1055 5060 -1043
rect 5260 -67 5318 -55
rect 5260 -1043 5272 -67
rect 5306 -1043 5318 -67
rect 5260 -1055 5318 -1043
rect 5518 -67 5576 -55
rect 5518 -1043 5530 -67
rect 5564 -1043 5576 -67
rect 5518 -1055 5576 -1043
rect 5776 -67 5834 -55
rect 5776 -1043 5788 -67
rect 5822 -1043 5834 -67
rect 5776 -1055 5834 -1043
rect 6034 -67 6092 -55
rect 6034 -1043 6046 -67
rect 6080 -1043 6092 -67
rect 6034 -1055 6092 -1043
rect 6292 -67 6350 -55
rect 6292 -1043 6304 -67
rect 6338 -1043 6350 -67
rect 6292 -1055 6350 -1043
rect 6550 -67 6608 -55
rect 6550 -1043 6562 -67
rect 6596 -1043 6608 -67
rect 6550 -1055 6608 -1043
rect 6808 -67 6866 -55
rect 6808 -1043 6820 -67
rect 6854 -1043 6866 -67
rect 6808 -1055 6866 -1043
rect 7066 -67 7124 -55
rect 7066 -1043 7078 -67
rect 7112 -1043 7124 -67
rect 7066 -1055 7124 -1043
rect -7124 -1177 -7066 -1165
rect -7124 -2153 -7112 -1177
rect -7078 -2153 -7066 -1177
rect -7124 -2165 -7066 -2153
rect -6866 -1177 -6808 -1165
rect -6866 -2153 -6854 -1177
rect -6820 -2153 -6808 -1177
rect -6866 -2165 -6808 -2153
rect -6608 -1177 -6550 -1165
rect -6608 -2153 -6596 -1177
rect -6562 -2153 -6550 -1177
rect -6608 -2165 -6550 -2153
rect -6350 -1177 -6292 -1165
rect -6350 -2153 -6338 -1177
rect -6304 -2153 -6292 -1177
rect -6350 -2165 -6292 -2153
rect -6092 -1177 -6034 -1165
rect -6092 -2153 -6080 -1177
rect -6046 -2153 -6034 -1177
rect -6092 -2165 -6034 -2153
rect -5834 -1177 -5776 -1165
rect -5834 -2153 -5822 -1177
rect -5788 -2153 -5776 -1177
rect -5834 -2165 -5776 -2153
rect -5576 -1177 -5518 -1165
rect -5576 -2153 -5564 -1177
rect -5530 -2153 -5518 -1177
rect -5576 -2165 -5518 -2153
rect -5318 -1177 -5260 -1165
rect -5318 -2153 -5306 -1177
rect -5272 -2153 -5260 -1177
rect -5318 -2165 -5260 -2153
rect -5060 -1177 -5002 -1165
rect -5060 -2153 -5048 -1177
rect -5014 -2153 -5002 -1177
rect -5060 -2165 -5002 -2153
rect -4802 -1177 -4744 -1165
rect -4802 -2153 -4790 -1177
rect -4756 -2153 -4744 -1177
rect -4802 -2165 -4744 -2153
rect -4544 -1177 -4486 -1165
rect -4544 -2153 -4532 -1177
rect -4498 -2153 -4486 -1177
rect -4544 -2165 -4486 -2153
rect -4286 -1177 -4228 -1165
rect -4286 -2153 -4274 -1177
rect -4240 -2153 -4228 -1177
rect -4286 -2165 -4228 -2153
rect -4028 -1177 -3970 -1165
rect -4028 -2153 -4016 -1177
rect -3982 -2153 -3970 -1177
rect -4028 -2165 -3970 -2153
rect -3770 -1177 -3712 -1165
rect -3770 -2153 -3758 -1177
rect -3724 -2153 -3712 -1177
rect -3770 -2165 -3712 -2153
rect -3512 -1177 -3454 -1165
rect -3512 -2153 -3500 -1177
rect -3466 -2153 -3454 -1177
rect -3512 -2165 -3454 -2153
rect -3254 -1177 -3196 -1165
rect -3254 -2153 -3242 -1177
rect -3208 -2153 -3196 -1177
rect -3254 -2165 -3196 -2153
rect -2996 -1177 -2938 -1165
rect -2996 -2153 -2984 -1177
rect -2950 -2153 -2938 -1177
rect -2996 -2165 -2938 -2153
rect -2738 -1177 -2680 -1165
rect -2738 -2153 -2726 -1177
rect -2692 -2153 -2680 -1177
rect -2738 -2165 -2680 -2153
rect -2480 -1177 -2422 -1165
rect -2480 -2153 -2468 -1177
rect -2434 -2153 -2422 -1177
rect -2480 -2165 -2422 -2153
rect -2222 -1177 -2164 -1165
rect -2222 -2153 -2210 -1177
rect -2176 -2153 -2164 -1177
rect -2222 -2165 -2164 -2153
rect -1964 -1177 -1906 -1165
rect -1964 -2153 -1952 -1177
rect -1918 -2153 -1906 -1177
rect -1964 -2165 -1906 -2153
rect -1706 -1177 -1648 -1165
rect -1706 -2153 -1694 -1177
rect -1660 -2153 -1648 -1177
rect -1706 -2165 -1648 -2153
rect -1448 -1177 -1390 -1165
rect -1448 -2153 -1436 -1177
rect -1402 -2153 -1390 -1177
rect -1448 -2165 -1390 -2153
rect -1190 -1177 -1132 -1165
rect -1190 -2153 -1178 -1177
rect -1144 -2153 -1132 -1177
rect -1190 -2165 -1132 -2153
rect -932 -1177 -874 -1165
rect -932 -2153 -920 -1177
rect -886 -2153 -874 -1177
rect -932 -2165 -874 -2153
rect -674 -1177 -616 -1165
rect -674 -2153 -662 -1177
rect -628 -2153 -616 -1177
rect -674 -2165 -616 -2153
rect -416 -1177 -358 -1165
rect -416 -2153 -404 -1177
rect -370 -2153 -358 -1177
rect -416 -2165 -358 -2153
rect -158 -1177 -100 -1165
rect -158 -2153 -146 -1177
rect -112 -2153 -100 -1177
rect -158 -2165 -100 -2153
rect 100 -1177 158 -1165
rect 100 -2153 112 -1177
rect 146 -2153 158 -1177
rect 100 -2165 158 -2153
rect 358 -1177 416 -1165
rect 358 -2153 370 -1177
rect 404 -2153 416 -1177
rect 358 -2165 416 -2153
rect 616 -1177 674 -1165
rect 616 -2153 628 -1177
rect 662 -2153 674 -1177
rect 616 -2165 674 -2153
rect 874 -1177 932 -1165
rect 874 -2153 886 -1177
rect 920 -2153 932 -1177
rect 874 -2165 932 -2153
rect 1132 -1177 1190 -1165
rect 1132 -2153 1144 -1177
rect 1178 -2153 1190 -1177
rect 1132 -2165 1190 -2153
rect 1390 -1177 1448 -1165
rect 1390 -2153 1402 -1177
rect 1436 -2153 1448 -1177
rect 1390 -2165 1448 -2153
rect 1648 -1177 1706 -1165
rect 1648 -2153 1660 -1177
rect 1694 -2153 1706 -1177
rect 1648 -2165 1706 -2153
rect 1906 -1177 1964 -1165
rect 1906 -2153 1918 -1177
rect 1952 -2153 1964 -1177
rect 1906 -2165 1964 -2153
rect 2164 -1177 2222 -1165
rect 2164 -2153 2176 -1177
rect 2210 -2153 2222 -1177
rect 2164 -2165 2222 -2153
rect 2422 -1177 2480 -1165
rect 2422 -2153 2434 -1177
rect 2468 -2153 2480 -1177
rect 2422 -2165 2480 -2153
rect 2680 -1177 2738 -1165
rect 2680 -2153 2692 -1177
rect 2726 -2153 2738 -1177
rect 2680 -2165 2738 -2153
rect 2938 -1177 2996 -1165
rect 2938 -2153 2950 -1177
rect 2984 -2153 2996 -1177
rect 2938 -2165 2996 -2153
rect 3196 -1177 3254 -1165
rect 3196 -2153 3208 -1177
rect 3242 -2153 3254 -1177
rect 3196 -2165 3254 -2153
rect 3454 -1177 3512 -1165
rect 3454 -2153 3466 -1177
rect 3500 -2153 3512 -1177
rect 3454 -2165 3512 -2153
rect 3712 -1177 3770 -1165
rect 3712 -2153 3724 -1177
rect 3758 -2153 3770 -1177
rect 3712 -2165 3770 -2153
rect 3970 -1177 4028 -1165
rect 3970 -2153 3982 -1177
rect 4016 -2153 4028 -1177
rect 3970 -2165 4028 -2153
rect 4228 -1177 4286 -1165
rect 4228 -2153 4240 -1177
rect 4274 -2153 4286 -1177
rect 4228 -2165 4286 -2153
rect 4486 -1177 4544 -1165
rect 4486 -2153 4498 -1177
rect 4532 -2153 4544 -1177
rect 4486 -2165 4544 -2153
rect 4744 -1177 4802 -1165
rect 4744 -2153 4756 -1177
rect 4790 -2153 4802 -1177
rect 4744 -2165 4802 -2153
rect 5002 -1177 5060 -1165
rect 5002 -2153 5014 -1177
rect 5048 -2153 5060 -1177
rect 5002 -2165 5060 -2153
rect 5260 -1177 5318 -1165
rect 5260 -2153 5272 -1177
rect 5306 -2153 5318 -1177
rect 5260 -2165 5318 -2153
rect 5518 -1177 5576 -1165
rect 5518 -2153 5530 -1177
rect 5564 -2153 5576 -1177
rect 5518 -2165 5576 -2153
rect 5776 -1177 5834 -1165
rect 5776 -2153 5788 -1177
rect 5822 -2153 5834 -1177
rect 5776 -2165 5834 -2153
rect 6034 -1177 6092 -1165
rect 6034 -2153 6046 -1177
rect 6080 -2153 6092 -1177
rect 6034 -2165 6092 -2153
rect 6292 -1177 6350 -1165
rect 6292 -2153 6304 -1177
rect 6338 -2153 6350 -1177
rect 6292 -2165 6350 -2153
rect 6550 -1177 6608 -1165
rect 6550 -2153 6562 -1177
rect 6596 -2153 6608 -1177
rect 6550 -2165 6608 -2153
rect 6808 -1177 6866 -1165
rect 6808 -2153 6820 -1177
rect 6854 -2153 6866 -1177
rect 6808 -2165 6866 -2153
rect 7066 -1177 7124 -1165
rect 7066 -2153 7078 -1177
rect 7112 -2153 7124 -1177
rect 7066 -2165 7124 -2153
<< mvndiffc >>
rect -7112 1177 -7078 2153
rect -6854 1177 -6820 2153
rect -6596 1177 -6562 2153
rect -6338 1177 -6304 2153
rect -6080 1177 -6046 2153
rect -5822 1177 -5788 2153
rect -5564 1177 -5530 2153
rect -5306 1177 -5272 2153
rect -5048 1177 -5014 2153
rect -4790 1177 -4756 2153
rect -4532 1177 -4498 2153
rect -4274 1177 -4240 2153
rect -4016 1177 -3982 2153
rect -3758 1177 -3724 2153
rect -3500 1177 -3466 2153
rect -3242 1177 -3208 2153
rect -2984 1177 -2950 2153
rect -2726 1177 -2692 2153
rect -2468 1177 -2434 2153
rect -2210 1177 -2176 2153
rect -1952 1177 -1918 2153
rect -1694 1177 -1660 2153
rect -1436 1177 -1402 2153
rect -1178 1177 -1144 2153
rect -920 1177 -886 2153
rect -662 1177 -628 2153
rect -404 1177 -370 2153
rect -146 1177 -112 2153
rect 112 1177 146 2153
rect 370 1177 404 2153
rect 628 1177 662 2153
rect 886 1177 920 2153
rect 1144 1177 1178 2153
rect 1402 1177 1436 2153
rect 1660 1177 1694 2153
rect 1918 1177 1952 2153
rect 2176 1177 2210 2153
rect 2434 1177 2468 2153
rect 2692 1177 2726 2153
rect 2950 1177 2984 2153
rect 3208 1177 3242 2153
rect 3466 1177 3500 2153
rect 3724 1177 3758 2153
rect 3982 1177 4016 2153
rect 4240 1177 4274 2153
rect 4498 1177 4532 2153
rect 4756 1177 4790 2153
rect 5014 1177 5048 2153
rect 5272 1177 5306 2153
rect 5530 1177 5564 2153
rect 5788 1177 5822 2153
rect 6046 1177 6080 2153
rect 6304 1177 6338 2153
rect 6562 1177 6596 2153
rect 6820 1177 6854 2153
rect 7078 1177 7112 2153
rect -7112 67 -7078 1043
rect -6854 67 -6820 1043
rect -6596 67 -6562 1043
rect -6338 67 -6304 1043
rect -6080 67 -6046 1043
rect -5822 67 -5788 1043
rect -5564 67 -5530 1043
rect -5306 67 -5272 1043
rect -5048 67 -5014 1043
rect -4790 67 -4756 1043
rect -4532 67 -4498 1043
rect -4274 67 -4240 1043
rect -4016 67 -3982 1043
rect -3758 67 -3724 1043
rect -3500 67 -3466 1043
rect -3242 67 -3208 1043
rect -2984 67 -2950 1043
rect -2726 67 -2692 1043
rect -2468 67 -2434 1043
rect -2210 67 -2176 1043
rect -1952 67 -1918 1043
rect -1694 67 -1660 1043
rect -1436 67 -1402 1043
rect -1178 67 -1144 1043
rect -920 67 -886 1043
rect -662 67 -628 1043
rect -404 67 -370 1043
rect -146 67 -112 1043
rect 112 67 146 1043
rect 370 67 404 1043
rect 628 67 662 1043
rect 886 67 920 1043
rect 1144 67 1178 1043
rect 1402 67 1436 1043
rect 1660 67 1694 1043
rect 1918 67 1952 1043
rect 2176 67 2210 1043
rect 2434 67 2468 1043
rect 2692 67 2726 1043
rect 2950 67 2984 1043
rect 3208 67 3242 1043
rect 3466 67 3500 1043
rect 3724 67 3758 1043
rect 3982 67 4016 1043
rect 4240 67 4274 1043
rect 4498 67 4532 1043
rect 4756 67 4790 1043
rect 5014 67 5048 1043
rect 5272 67 5306 1043
rect 5530 67 5564 1043
rect 5788 67 5822 1043
rect 6046 67 6080 1043
rect 6304 67 6338 1043
rect 6562 67 6596 1043
rect 6820 67 6854 1043
rect 7078 67 7112 1043
rect -7112 -1043 -7078 -67
rect -6854 -1043 -6820 -67
rect -6596 -1043 -6562 -67
rect -6338 -1043 -6304 -67
rect -6080 -1043 -6046 -67
rect -5822 -1043 -5788 -67
rect -5564 -1043 -5530 -67
rect -5306 -1043 -5272 -67
rect -5048 -1043 -5014 -67
rect -4790 -1043 -4756 -67
rect -4532 -1043 -4498 -67
rect -4274 -1043 -4240 -67
rect -4016 -1043 -3982 -67
rect -3758 -1043 -3724 -67
rect -3500 -1043 -3466 -67
rect -3242 -1043 -3208 -67
rect -2984 -1043 -2950 -67
rect -2726 -1043 -2692 -67
rect -2468 -1043 -2434 -67
rect -2210 -1043 -2176 -67
rect -1952 -1043 -1918 -67
rect -1694 -1043 -1660 -67
rect -1436 -1043 -1402 -67
rect -1178 -1043 -1144 -67
rect -920 -1043 -886 -67
rect -662 -1043 -628 -67
rect -404 -1043 -370 -67
rect -146 -1043 -112 -67
rect 112 -1043 146 -67
rect 370 -1043 404 -67
rect 628 -1043 662 -67
rect 886 -1043 920 -67
rect 1144 -1043 1178 -67
rect 1402 -1043 1436 -67
rect 1660 -1043 1694 -67
rect 1918 -1043 1952 -67
rect 2176 -1043 2210 -67
rect 2434 -1043 2468 -67
rect 2692 -1043 2726 -67
rect 2950 -1043 2984 -67
rect 3208 -1043 3242 -67
rect 3466 -1043 3500 -67
rect 3724 -1043 3758 -67
rect 3982 -1043 4016 -67
rect 4240 -1043 4274 -67
rect 4498 -1043 4532 -67
rect 4756 -1043 4790 -67
rect 5014 -1043 5048 -67
rect 5272 -1043 5306 -67
rect 5530 -1043 5564 -67
rect 5788 -1043 5822 -67
rect 6046 -1043 6080 -67
rect 6304 -1043 6338 -67
rect 6562 -1043 6596 -67
rect 6820 -1043 6854 -67
rect 7078 -1043 7112 -67
rect -7112 -2153 -7078 -1177
rect -6854 -2153 -6820 -1177
rect -6596 -2153 -6562 -1177
rect -6338 -2153 -6304 -1177
rect -6080 -2153 -6046 -1177
rect -5822 -2153 -5788 -1177
rect -5564 -2153 -5530 -1177
rect -5306 -2153 -5272 -1177
rect -5048 -2153 -5014 -1177
rect -4790 -2153 -4756 -1177
rect -4532 -2153 -4498 -1177
rect -4274 -2153 -4240 -1177
rect -4016 -2153 -3982 -1177
rect -3758 -2153 -3724 -1177
rect -3500 -2153 -3466 -1177
rect -3242 -2153 -3208 -1177
rect -2984 -2153 -2950 -1177
rect -2726 -2153 -2692 -1177
rect -2468 -2153 -2434 -1177
rect -2210 -2153 -2176 -1177
rect -1952 -2153 -1918 -1177
rect -1694 -2153 -1660 -1177
rect -1436 -2153 -1402 -1177
rect -1178 -2153 -1144 -1177
rect -920 -2153 -886 -1177
rect -662 -2153 -628 -1177
rect -404 -2153 -370 -1177
rect -146 -2153 -112 -1177
rect 112 -2153 146 -1177
rect 370 -2153 404 -1177
rect 628 -2153 662 -1177
rect 886 -2153 920 -1177
rect 1144 -2153 1178 -1177
rect 1402 -2153 1436 -1177
rect 1660 -2153 1694 -1177
rect 1918 -2153 1952 -1177
rect 2176 -2153 2210 -1177
rect 2434 -2153 2468 -1177
rect 2692 -2153 2726 -1177
rect 2950 -2153 2984 -1177
rect 3208 -2153 3242 -1177
rect 3466 -2153 3500 -1177
rect 3724 -2153 3758 -1177
rect 3982 -2153 4016 -1177
rect 4240 -2153 4274 -1177
rect 4498 -2153 4532 -1177
rect 4756 -2153 4790 -1177
rect 5014 -2153 5048 -1177
rect 5272 -2153 5306 -1177
rect 5530 -2153 5564 -1177
rect 5788 -2153 5822 -1177
rect 6046 -2153 6080 -1177
rect 6304 -2153 6338 -1177
rect 6562 -2153 6596 -1177
rect 6820 -2153 6854 -1177
rect 7078 -2153 7112 -1177
<< mvpsubdiff >>
rect -7258 2375 7258 2387
rect -7258 2341 -7150 2375
rect 7150 2341 7258 2375
rect -7258 2329 7258 2341
rect -7258 2279 -7200 2329
rect -7258 -2279 -7246 2279
rect -7212 -2279 -7200 2279
rect 7200 2279 7258 2329
rect -7258 -2329 -7200 -2279
rect 7200 -2279 7212 2279
rect 7246 -2279 7258 2279
rect 7200 -2329 7258 -2279
rect -7258 -2341 7258 -2329
rect -7258 -2375 -7150 -2341
rect 7150 -2375 7258 -2341
rect -7258 -2387 7258 -2375
<< mvpsubdiffcont >>
rect -7150 2341 7150 2375
rect -7246 -2279 -7212 2279
rect 7212 -2279 7246 2279
rect -7150 -2375 7150 -2341
<< poly >>
rect -7066 2237 -6866 2253
rect -7066 2203 -7050 2237
rect -6882 2203 -6866 2237
rect -7066 2165 -6866 2203
rect -6808 2237 -6608 2253
rect -6808 2203 -6792 2237
rect -6624 2203 -6608 2237
rect -6808 2165 -6608 2203
rect -6550 2237 -6350 2253
rect -6550 2203 -6534 2237
rect -6366 2203 -6350 2237
rect -6550 2165 -6350 2203
rect -6292 2237 -6092 2253
rect -6292 2203 -6276 2237
rect -6108 2203 -6092 2237
rect -6292 2165 -6092 2203
rect -6034 2237 -5834 2253
rect -6034 2203 -6018 2237
rect -5850 2203 -5834 2237
rect -6034 2165 -5834 2203
rect -5776 2237 -5576 2253
rect -5776 2203 -5760 2237
rect -5592 2203 -5576 2237
rect -5776 2165 -5576 2203
rect -5518 2237 -5318 2253
rect -5518 2203 -5502 2237
rect -5334 2203 -5318 2237
rect -5518 2165 -5318 2203
rect -5260 2237 -5060 2253
rect -5260 2203 -5244 2237
rect -5076 2203 -5060 2237
rect -5260 2165 -5060 2203
rect -5002 2237 -4802 2253
rect -5002 2203 -4986 2237
rect -4818 2203 -4802 2237
rect -5002 2165 -4802 2203
rect -4744 2237 -4544 2253
rect -4744 2203 -4728 2237
rect -4560 2203 -4544 2237
rect -4744 2165 -4544 2203
rect -4486 2237 -4286 2253
rect -4486 2203 -4470 2237
rect -4302 2203 -4286 2237
rect -4486 2165 -4286 2203
rect -4228 2237 -4028 2253
rect -4228 2203 -4212 2237
rect -4044 2203 -4028 2237
rect -4228 2165 -4028 2203
rect -3970 2237 -3770 2253
rect -3970 2203 -3954 2237
rect -3786 2203 -3770 2237
rect -3970 2165 -3770 2203
rect -3712 2237 -3512 2253
rect -3712 2203 -3696 2237
rect -3528 2203 -3512 2237
rect -3712 2165 -3512 2203
rect -3454 2237 -3254 2253
rect -3454 2203 -3438 2237
rect -3270 2203 -3254 2237
rect -3454 2165 -3254 2203
rect -3196 2237 -2996 2253
rect -3196 2203 -3180 2237
rect -3012 2203 -2996 2237
rect -3196 2165 -2996 2203
rect -2938 2237 -2738 2253
rect -2938 2203 -2922 2237
rect -2754 2203 -2738 2237
rect -2938 2165 -2738 2203
rect -2680 2237 -2480 2253
rect -2680 2203 -2664 2237
rect -2496 2203 -2480 2237
rect -2680 2165 -2480 2203
rect -2422 2237 -2222 2253
rect -2422 2203 -2406 2237
rect -2238 2203 -2222 2237
rect -2422 2165 -2222 2203
rect -2164 2237 -1964 2253
rect -2164 2203 -2148 2237
rect -1980 2203 -1964 2237
rect -2164 2165 -1964 2203
rect -1906 2237 -1706 2253
rect -1906 2203 -1890 2237
rect -1722 2203 -1706 2237
rect -1906 2165 -1706 2203
rect -1648 2237 -1448 2253
rect -1648 2203 -1632 2237
rect -1464 2203 -1448 2237
rect -1648 2165 -1448 2203
rect -1390 2237 -1190 2253
rect -1390 2203 -1374 2237
rect -1206 2203 -1190 2237
rect -1390 2165 -1190 2203
rect -1132 2237 -932 2253
rect -1132 2203 -1116 2237
rect -948 2203 -932 2237
rect -1132 2165 -932 2203
rect -874 2237 -674 2253
rect -874 2203 -858 2237
rect -690 2203 -674 2237
rect -874 2165 -674 2203
rect -616 2237 -416 2253
rect -616 2203 -600 2237
rect -432 2203 -416 2237
rect -616 2165 -416 2203
rect -358 2237 -158 2253
rect -358 2203 -342 2237
rect -174 2203 -158 2237
rect -358 2165 -158 2203
rect -100 2237 100 2253
rect -100 2203 -84 2237
rect 84 2203 100 2237
rect -100 2165 100 2203
rect 158 2237 358 2253
rect 158 2203 174 2237
rect 342 2203 358 2237
rect 158 2165 358 2203
rect 416 2237 616 2253
rect 416 2203 432 2237
rect 600 2203 616 2237
rect 416 2165 616 2203
rect 674 2237 874 2253
rect 674 2203 690 2237
rect 858 2203 874 2237
rect 674 2165 874 2203
rect 932 2237 1132 2253
rect 932 2203 948 2237
rect 1116 2203 1132 2237
rect 932 2165 1132 2203
rect 1190 2237 1390 2253
rect 1190 2203 1206 2237
rect 1374 2203 1390 2237
rect 1190 2165 1390 2203
rect 1448 2237 1648 2253
rect 1448 2203 1464 2237
rect 1632 2203 1648 2237
rect 1448 2165 1648 2203
rect 1706 2237 1906 2253
rect 1706 2203 1722 2237
rect 1890 2203 1906 2237
rect 1706 2165 1906 2203
rect 1964 2237 2164 2253
rect 1964 2203 1980 2237
rect 2148 2203 2164 2237
rect 1964 2165 2164 2203
rect 2222 2237 2422 2253
rect 2222 2203 2238 2237
rect 2406 2203 2422 2237
rect 2222 2165 2422 2203
rect 2480 2237 2680 2253
rect 2480 2203 2496 2237
rect 2664 2203 2680 2237
rect 2480 2165 2680 2203
rect 2738 2237 2938 2253
rect 2738 2203 2754 2237
rect 2922 2203 2938 2237
rect 2738 2165 2938 2203
rect 2996 2237 3196 2253
rect 2996 2203 3012 2237
rect 3180 2203 3196 2237
rect 2996 2165 3196 2203
rect 3254 2237 3454 2253
rect 3254 2203 3270 2237
rect 3438 2203 3454 2237
rect 3254 2165 3454 2203
rect 3512 2237 3712 2253
rect 3512 2203 3528 2237
rect 3696 2203 3712 2237
rect 3512 2165 3712 2203
rect 3770 2237 3970 2253
rect 3770 2203 3786 2237
rect 3954 2203 3970 2237
rect 3770 2165 3970 2203
rect 4028 2237 4228 2253
rect 4028 2203 4044 2237
rect 4212 2203 4228 2237
rect 4028 2165 4228 2203
rect 4286 2237 4486 2253
rect 4286 2203 4302 2237
rect 4470 2203 4486 2237
rect 4286 2165 4486 2203
rect 4544 2237 4744 2253
rect 4544 2203 4560 2237
rect 4728 2203 4744 2237
rect 4544 2165 4744 2203
rect 4802 2237 5002 2253
rect 4802 2203 4818 2237
rect 4986 2203 5002 2237
rect 4802 2165 5002 2203
rect 5060 2237 5260 2253
rect 5060 2203 5076 2237
rect 5244 2203 5260 2237
rect 5060 2165 5260 2203
rect 5318 2237 5518 2253
rect 5318 2203 5334 2237
rect 5502 2203 5518 2237
rect 5318 2165 5518 2203
rect 5576 2237 5776 2253
rect 5576 2203 5592 2237
rect 5760 2203 5776 2237
rect 5576 2165 5776 2203
rect 5834 2237 6034 2253
rect 5834 2203 5850 2237
rect 6018 2203 6034 2237
rect 5834 2165 6034 2203
rect 6092 2237 6292 2253
rect 6092 2203 6108 2237
rect 6276 2203 6292 2237
rect 6092 2165 6292 2203
rect 6350 2237 6550 2253
rect 6350 2203 6366 2237
rect 6534 2203 6550 2237
rect 6350 2165 6550 2203
rect 6608 2237 6808 2253
rect 6608 2203 6624 2237
rect 6792 2203 6808 2237
rect 6608 2165 6808 2203
rect 6866 2237 7066 2253
rect 6866 2203 6882 2237
rect 7050 2203 7066 2237
rect 6866 2165 7066 2203
rect -7066 1127 -6866 1165
rect -7066 1093 -7050 1127
rect -6882 1093 -6866 1127
rect -7066 1055 -6866 1093
rect -6808 1127 -6608 1165
rect -6808 1093 -6792 1127
rect -6624 1093 -6608 1127
rect -6808 1055 -6608 1093
rect -6550 1127 -6350 1165
rect -6550 1093 -6534 1127
rect -6366 1093 -6350 1127
rect -6550 1055 -6350 1093
rect -6292 1127 -6092 1165
rect -6292 1093 -6276 1127
rect -6108 1093 -6092 1127
rect -6292 1055 -6092 1093
rect -6034 1127 -5834 1165
rect -6034 1093 -6018 1127
rect -5850 1093 -5834 1127
rect -6034 1055 -5834 1093
rect -5776 1127 -5576 1165
rect -5776 1093 -5760 1127
rect -5592 1093 -5576 1127
rect -5776 1055 -5576 1093
rect -5518 1127 -5318 1165
rect -5518 1093 -5502 1127
rect -5334 1093 -5318 1127
rect -5518 1055 -5318 1093
rect -5260 1127 -5060 1165
rect -5260 1093 -5244 1127
rect -5076 1093 -5060 1127
rect -5260 1055 -5060 1093
rect -5002 1127 -4802 1165
rect -5002 1093 -4986 1127
rect -4818 1093 -4802 1127
rect -5002 1055 -4802 1093
rect -4744 1127 -4544 1165
rect -4744 1093 -4728 1127
rect -4560 1093 -4544 1127
rect -4744 1055 -4544 1093
rect -4486 1127 -4286 1165
rect -4486 1093 -4470 1127
rect -4302 1093 -4286 1127
rect -4486 1055 -4286 1093
rect -4228 1127 -4028 1165
rect -4228 1093 -4212 1127
rect -4044 1093 -4028 1127
rect -4228 1055 -4028 1093
rect -3970 1127 -3770 1165
rect -3970 1093 -3954 1127
rect -3786 1093 -3770 1127
rect -3970 1055 -3770 1093
rect -3712 1127 -3512 1165
rect -3712 1093 -3696 1127
rect -3528 1093 -3512 1127
rect -3712 1055 -3512 1093
rect -3454 1127 -3254 1165
rect -3454 1093 -3438 1127
rect -3270 1093 -3254 1127
rect -3454 1055 -3254 1093
rect -3196 1127 -2996 1165
rect -3196 1093 -3180 1127
rect -3012 1093 -2996 1127
rect -3196 1055 -2996 1093
rect -2938 1127 -2738 1165
rect -2938 1093 -2922 1127
rect -2754 1093 -2738 1127
rect -2938 1055 -2738 1093
rect -2680 1127 -2480 1165
rect -2680 1093 -2664 1127
rect -2496 1093 -2480 1127
rect -2680 1055 -2480 1093
rect -2422 1127 -2222 1165
rect -2422 1093 -2406 1127
rect -2238 1093 -2222 1127
rect -2422 1055 -2222 1093
rect -2164 1127 -1964 1165
rect -2164 1093 -2148 1127
rect -1980 1093 -1964 1127
rect -2164 1055 -1964 1093
rect -1906 1127 -1706 1165
rect -1906 1093 -1890 1127
rect -1722 1093 -1706 1127
rect -1906 1055 -1706 1093
rect -1648 1127 -1448 1165
rect -1648 1093 -1632 1127
rect -1464 1093 -1448 1127
rect -1648 1055 -1448 1093
rect -1390 1127 -1190 1165
rect -1390 1093 -1374 1127
rect -1206 1093 -1190 1127
rect -1390 1055 -1190 1093
rect -1132 1127 -932 1165
rect -1132 1093 -1116 1127
rect -948 1093 -932 1127
rect -1132 1055 -932 1093
rect -874 1127 -674 1165
rect -874 1093 -858 1127
rect -690 1093 -674 1127
rect -874 1055 -674 1093
rect -616 1127 -416 1165
rect -616 1093 -600 1127
rect -432 1093 -416 1127
rect -616 1055 -416 1093
rect -358 1127 -158 1165
rect -358 1093 -342 1127
rect -174 1093 -158 1127
rect -358 1055 -158 1093
rect -100 1127 100 1165
rect -100 1093 -84 1127
rect 84 1093 100 1127
rect -100 1055 100 1093
rect 158 1127 358 1165
rect 158 1093 174 1127
rect 342 1093 358 1127
rect 158 1055 358 1093
rect 416 1127 616 1165
rect 416 1093 432 1127
rect 600 1093 616 1127
rect 416 1055 616 1093
rect 674 1127 874 1165
rect 674 1093 690 1127
rect 858 1093 874 1127
rect 674 1055 874 1093
rect 932 1127 1132 1165
rect 932 1093 948 1127
rect 1116 1093 1132 1127
rect 932 1055 1132 1093
rect 1190 1127 1390 1165
rect 1190 1093 1206 1127
rect 1374 1093 1390 1127
rect 1190 1055 1390 1093
rect 1448 1127 1648 1165
rect 1448 1093 1464 1127
rect 1632 1093 1648 1127
rect 1448 1055 1648 1093
rect 1706 1127 1906 1165
rect 1706 1093 1722 1127
rect 1890 1093 1906 1127
rect 1706 1055 1906 1093
rect 1964 1127 2164 1165
rect 1964 1093 1980 1127
rect 2148 1093 2164 1127
rect 1964 1055 2164 1093
rect 2222 1127 2422 1165
rect 2222 1093 2238 1127
rect 2406 1093 2422 1127
rect 2222 1055 2422 1093
rect 2480 1127 2680 1165
rect 2480 1093 2496 1127
rect 2664 1093 2680 1127
rect 2480 1055 2680 1093
rect 2738 1127 2938 1165
rect 2738 1093 2754 1127
rect 2922 1093 2938 1127
rect 2738 1055 2938 1093
rect 2996 1127 3196 1165
rect 2996 1093 3012 1127
rect 3180 1093 3196 1127
rect 2996 1055 3196 1093
rect 3254 1127 3454 1165
rect 3254 1093 3270 1127
rect 3438 1093 3454 1127
rect 3254 1055 3454 1093
rect 3512 1127 3712 1165
rect 3512 1093 3528 1127
rect 3696 1093 3712 1127
rect 3512 1055 3712 1093
rect 3770 1127 3970 1165
rect 3770 1093 3786 1127
rect 3954 1093 3970 1127
rect 3770 1055 3970 1093
rect 4028 1127 4228 1165
rect 4028 1093 4044 1127
rect 4212 1093 4228 1127
rect 4028 1055 4228 1093
rect 4286 1127 4486 1165
rect 4286 1093 4302 1127
rect 4470 1093 4486 1127
rect 4286 1055 4486 1093
rect 4544 1127 4744 1165
rect 4544 1093 4560 1127
rect 4728 1093 4744 1127
rect 4544 1055 4744 1093
rect 4802 1127 5002 1165
rect 4802 1093 4818 1127
rect 4986 1093 5002 1127
rect 4802 1055 5002 1093
rect 5060 1127 5260 1165
rect 5060 1093 5076 1127
rect 5244 1093 5260 1127
rect 5060 1055 5260 1093
rect 5318 1127 5518 1165
rect 5318 1093 5334 1127
rect 5502 1093 5518 1127
rect 5318 1055 5518 1093
rect 5576 1127 5776 1165
rect 5576 1093 5592 1127
rect 5760 1093 5776 1127
rect 5576 1055 5776 1093
rect 5834 1127 6034 1165
rect 5834 1093 5850 1127
rect 6018 1093 6034 1127
rect 5834 1055 6034 1093
rect 6092 1127 6292 1165
rect 6092 1093 6108 1127
rect 6276 1093 6292 1127
rect 6092 1055 6292 1093
rect 6350 1127 6550 1165
rect 6350 1093 6366 1127
rect 6534 1093 6550 1127
rect 6350 1055 6550 1093
rect 6608 1127 6808 1165
rect 6608 1093 6624 1127
rect 6792 1093 6808 1127
rect 6608 1055 6808 1093
rect 6866 1127 7066 1165
rect 6866 1093 6882 1127
rect 7050 1093 7066 1127
rect 6866 1055 7066 1093
rect -7066 17 -6866 55
rect -7066 -17 -7050 17
rect -6882 -17 -6866 17
rect -7066 -55 -6866 -17
rect -6808 17 -6608 55
rect -6808 -17 -6792 17
rect -6624 -17 -6608 17
rect -6808 -55 -6608 -17
rect -6550 17 -6350 55
rect -6550 -17 -6534 17
rect -6366 -17 -6350 17
rect -6550 -55 -6350 -17
rect -6292 17 -6092 55
rect -6292 -17 -6276 17
rect -6108 -17 -6092 17
rect -6292 -55 -6092 -17
rect -6034 17 -5834 55
rect -6034 -17 -6018 17
rect -5850 -17 -5834 17
rect -6034 -55 -5834 -17
rect -5776 17 -5576 55
rect -5776 -17 -5760 17
rect -5592 -17 -5576 17
rect -5776 -55 -5576 -17
rect -5518 17 -5318 55
rect -5518 -17 -5502 17
rect -5334 -17 -5318 17
rect -5518 -55 -5318 -17
rect -5260 17 -5060 55
rect -5260 -17 -5244 17
rect -5076 -17 -5060 17
rect -5260 -55 -5060 -17
rect -5002 17 -4802 55
rect -5002 -17 -4986 17
rect -4818 -17 -4802 17
rect -5002 -55 -4802 -17
rect -4744 17 -4544 55
rect -4744 -17 -4728 17
rect -4560 -17 -4544 17
rect -4744 -55 -4544 -17
rect -4486 17 -4286 55
rect -4486 -17 -4470 17
rect -4302 -17 -4286 17
rect -4486 -55 -4286 -17
rect -4228 17 -4028 55
rect -4228 -17 -4212 17
rect -4044 -17 -4028 17
rect -4228 -55 -4028 -17
rect -3970 17 -3770 55
rect -3970 -17 -3954 17
rect -3786 -17 -3770 17
rect -3970 -55 -3770 -17
rect -3712 17 -3512 55
rect -3712 -17 -3696 17
rect -3528 -17 -3512 17
rect -3712 -55 -3512 -17
rect -3454 17 -3254 55
rect -3454 -17 -3438 17
rect -3270 -17 -3254 17
rect -3454 -55 -3254 -17
rect -3196 17 -2996 55
rect -3196 -17 -3180 17
rect -3012 -17 -2996 17
rect -3196 -55 -2996 -17
rect -2938 17 -2738 55
rect -2938 -17 -2922 17
rect -2754 -17 -2738 17
rect -2938 -55 -2738 -17
rect -2680 17 -2480 55
rect -2680 -17 -2664 17
rect -2496 -17 -2480 17
rect -2680 -55 -2480 -17
rect -2422 17 -2222 55
rect -2422 -17 -2406 17
rect -2238 -17 -2222 17
rect -2422 -55 -2222 -17
rect -2164 17 -1964 55
rect -2164 -17 -2148 17
rect -1980 -17 -1964 17
rect -2164 -55 -1964 -17
rect -1906 17 -1706 55
rect -1906 -17 -1890 17
rect -1722 -17 -1706 17
rect -1906 -55 -1706 -17
rect -1648 17 -1448 55
rect -1648 -17 -1632 17
rect -1464 -17 -1448 17
rect -1648 -55 -1448 -17
rect -1390 17 -1190 55
rect -1390 -17 -1374 17
rect -1206 -17 -1190 17
rect -1390 -55 -1190 -17
rect -1132 17 -932 55
rect -1132 -17 -1116 17
rect -948 -17 -932 17
rect -1132 -55 -932 -17
rect -874 17 -674 55
rect -874 -17 -858 17
rect -690 -17 -674 17
rect -874 -55 -674 -17
rect -616 17 -416 55
rect -616 -17 -600 17
rect -432 -17 -416 17
rect -616 -55 -416 -17
rect -358 17 -158 55
rect -358 -17 -342 17
rect -174 -17 -158 17
rect -358 -55 -158 -17
rect -100 17 100 55
rect -100 -17 -84 17
rect 84 -17 100 17
rect -100 -55 100 -17
rect 158 17 358 55
rect 158 -17 174 17
rect 342 -17 358 17
rect 158 -55 358 -17
rect 416 17 616 55
rect 416 -17 432 17
rect 600 -17 616 17
rect 416 -55 616 -17
rect 674 17 874 55
rect 674 -17 690 17
rect 858 -17 874 17
rect 674 -55 874 -17
rect 932 17 1132 55
rect 932 -17 948 17
rect 1116 -17 1132 17
rect 932 -55 1132 -17
rect 1190 17 1390 55
rect 1190 -17 1206 17
rect 1374 -17 1390 17
rect 1190 -55 1390 -17
rect 1448 17 1648 55
rect 1448 -17 1464 17
rect 1632 -17 1648 17
rect 1448 -55 1648 -17
rect 1706 17 1906 55
rect 1706 -17 1722 17
rect 1890 -17 1906 17
rect 1706 -55 1906 -17
rect 1964 17 2164 55
rect 1964 -17 1980 17
rect 2148 -17 2164 17
rect 1964 -55 2164 -17
rect 2222 17 2422 55
rect 2222 -17 2238 17
rect 2406 -17 2422 17
rect 2222 -55 2422 -17
rect 2480 17 2680 55
rect 2480 -17 2496 17
rect 2664 -17 2680 17
rect 2480 -55 2680 -17
rect 2738 17 2938 55
rect 2738 -17 2754 17
rect 2922 -17 2938 17
rect 2738 -55 2938 -17
rect 2996 17 3196 55
rect 2996 -17 3012 17
rect 3180 -17 3196 17
rect 2996 -55 3196 -17
rect 3254 17 3454 55
rect 3254 -17 3270 17
rect 3438 -17 3454 17
rect 3254 -55 3454 -17
rect 3512 17 3712 55
rect 3512 -17 3528 17
rect 3696 -17 3712 17
rect 3512 -55 3712 -17
rect 3770 17 3970 55
rect 3770 -17 3786 17
rect 3954 -17 3970 17
rect 3770 -55 3970 -17
rect 4028 17 4228 55
rect 4028 -17 4044 17
rect 4212 -17 4228 17
rect 4028 -55 4228 -17
rect 4286 17 4486 55
rect 4286 -17 4302 17
rect 4470 -17 4486 17
rect 4286 -55 4486 -17
rect 4544 17 4744 55
rect 4544 -17 4560 17
rect 4728 -17 4744 17
rect 4544 -55 4744 -17
rect 4802 17 5002 55
rect 4802 -17 4818 17
rect 4986 -17 5002 17
rect 4802 -55 5002 -17
rect 5060 17 5260 55
rect 5060 -17 5076 17
rect 5244 -17 5260 17
rect 5060 -55 5260 -17
rect 5318 17 5518 55
rect 5318 -17 5334 17
rect 5502 -17 5518 17
rect 5318 -55 5518 -17
rect 5576 17 5776 55
rect 5576 -17 5592 17
rect 5760 -17 5776 17
rect 5576 -55 5776 -17
rect 5834 17 6034 55
rect 5834 -17 5850 17
rect 6018 -17 6034 17
rect 5834 -55 6034 -17
rect 6092 17 6292 55
rect 6092 -17 6108 17
rect 6276 -17 6292 17
rect 6092 -55 6292 -17
rect 6350 17 6550 55
rect 6350 -17 6366 17
rect 6534 -17 6550 17
rect 6350 -55 6550 -17
rect 6608 17 6808 55
rect 6608 -17 6624 17
rect 6792 -17 6808 17
rect 6608 -55 6808 -17
rect 6866 17 7066 55
rect 6866 -17 6882 17
rect 7050 -17 7066 17
rect 6866 -55 7066 -17
rect -7066 -1093 -6866 -1055
rect -7066 -1127 -7050 -1093
rect -6882 -1127 -6866 -1093
rect -7066 -1165 -6866 -1127
rect -6808 -1093 -6608 -1055
rect -6808 -1127 -6792 -1093
rect -6624 -1127 -6608 -1093
rect -6808 -1165 -6608 -1127
rect -6550 -1093 -6350 -1055
rect -6550 -1127 -6534 -1093
rect -6366 -1127 -6350 -1093
rect -6550 -1165 -6350 -1127
rect -6292 -1093 -6092 -1055
rect -6292 -1127 -6276 -1093
rect -6108 -1127 -6092 -1093
rect -6292 -1165 -6092 -1127
rect -6034 -1093 -5834 -1055
rect -6034 -1127 -6018 -1093
rect -5850 -1127 -5834 -1093
rect -6034 -1165 -5834 -1127
rect -5776 -1093 -5576 -1055
rect -5776 -1127 -5760 -1093
rect -5592 -1127 -5576 -1093
rect -5776 -1165 -5576 -1127
rect -5518 -1093 -5318 -1055
rect -5518 -1127 -5502 -1093
rect -5334 -1127 -5318 -1093
rect -5518 -1165 -5318 -1127
rect -5260 -1093 -5060 -1055
rect -5260 -1127 -5244 -1093
rect -5076 -1127 -5060 -1093
rect -5260 -1165 -5060 -1127
rect -5002 -1093 -4802 -1055
rect -5002 -1127 -4986 -1093
rect -4818 -1127 -4802 -1093
rect -5002 -1165 -4802 -1127
rect -4744 -1093 -4544 -1055
rect -4744 -1127 -4728 -1093
rect -4560 -1127 -4544 -1093
rect -4744 -1165 -4544 -1127
rect -4486 -1093 -4286 -1055
rect -4486 -1127 -4470 -1093
rect -4302 -1127 -4286 -1093
rect -4486 -1165 -4286 -1127
rect -4228 -1093 -4028 -1055
rect -4228 -1127 -4212 -1093
rect -4044 -1127 -4028 -1093
rect -4228 -1165 -4028 -1127
rect -3970 -1093 -3770 -1055
rect -3970 -1127 -3954 -1093
rect -3786 -1127 -3770 -1093
rect -3970 -1165 -3770 -1127
rect -3712 -1093 -3512 -1055
rect -3712 -1127 -3696 -1093
rect -3528 -1127 -3512 -1093
rect -3712 -1165 -3512 -1127
rect -3454 -1093 -3254 -1055
rect -3454 -1127 -3438 -1093
rect -3270 -1127 -3254 -1093
rect -3454 -1165 -3254 -1127
rect -3196 -1093 -2996 -1055
rect -3196 -1127 -3180 -1093
rect -3012 -1127 -2996 -1093
rect -3196 -1165 -2996 -1127
rect -2938 -1093 -2738 -1055
rect -2938 -1127 -2922 -1093
rect -2754 -1127 -2738 -1093
rect -2938 -1165 -2738 -1127
rect -2680 -1093 -2480 -1055
rect -2680 -1127 -2664 -1093
rect -2496 -1127 -2480 -1093
rect -2680 -1165 -2480 -1127
rect -2422 -1093 -2222 -1055
rect -2422 -1127 -2406 -1093
rect -2238 -1127 -2222 -1093
rect -2422 -1165 -2222 -1127
rect -2164 -1093 -1964 -1055
rect -2164 -1127 -2148 -1093
rect -1980 -1127 -1964 -1093
rect -2164 -1165 -1964 -1127
rect -1906 -1093 -1706 -1055
rect -1906 -1127 -1890 -1093
rect -1722 -1127 -1706 -1093
rect -1906 -1165 -1706 -1127
rect -1648 -1093 -1448 -1055
rect -1648 -1127 -1632 -1093
rect -1464 -1127 -1448 -1093
rect -1648 -1165 -1448 -1127
rect -1390 -1093 -1190 -1055
rect -1390 -1127 -1374 -1093
rect -1206 -1127 -1190 -1093
rect -1390 -1165 -1190 -1127
rect -1132 -1093 -932 -1055
rect -1132 -1127 -1116 -1093
rect -948 -1127 -932 -1093
rect -1132 -1165 -932 -1127
rect -874 -1093 -674 -1055
rect -874 -1127 -858 -1093
rect -690 -1127 -674 -1093
rect -874 -1165 -674 -1127
rect -616 -1093 -416 -1055
rect -616 -1127 -600 -1093
rect -432 -1127 -416 -1093
rect -616 -1165 -416 -1127
rect -358 -1093 -158 -1055
rect -358 -1127 -342 -1093
rect -174 -1127 -158 -1093
rect -358 -1165 -158 -1127
rect -100 -1093 100 -1055
rect -100 -1127 -84 -1093
rect 84 -1127 100 -1093
rect -100 -1165 100 -1127
rect 158 -1093 358 -1055
rect 158 -1127 174 -1093
rect 342 -1127 358 -1093
rect 158 -1165 358 -1127
rect 416 -1093 616 -1055
rect 416 -1127 432 -1093
rect 600 -1127 616 -1093
rect 416 -1165 616 -1127
rect 674 -1093 874 -1055
rect 674 -1127 690 -1093
rect 858 -1127 874 -1093
rect 674 -1165 874 -1127
rect 932 -1093 1132 -1055
rect 932 -1127 948 -1093
rect 1116 -1127 1132 -1093
rect 932 -1165 1132 -1127
rect 1190 -1093 1390 -1055
rect 1190 -1127 1206 -1093
rect 1374 -1127 1390 -1093
rect 1190 -1165 1390 -1127
rect 1448 -1093 1648 -1055
rect 1448 -1127 1464 -1093
rect 1632 -1127 1648 -1093
rect 1448 -1165 1648 -1127
rect 1706 -1093 1906 -1055
rect 1706 -1127 1722 -1093
rect 1890 -1127 1906 -1093
rect 1706 -1165 1906 -1127
rect 1964 -1093 2164 -1055
rect 1964 -1127 1980 -1093
rect 2148 -1127 2164 -1093
rect 1964 -1165 2164 -1127
rect 2222 -1093 2422 -1055
rect 2222 -1127 2238 -1093
rect 2406 -1127 2422 -1093
rect 2222 -1165 2422 -1127
rect 2480 -1093 2680 -1055
rect 2480 -1127 2496 -1093
rect 2664 -1127 2680 -1093
rect 2480 -1165 2680 -1127
rect 2738 -1093 2938 -1055
rect 2738 -1127 2754 -1093
rect 2922 -1127 2938 -1093
rect 2738 -1165 2938 -1127
rect 2996 -1093 3196 -1055
rect 2996 -1127 3012 -1093
rect 3180 -1127 3196 -1093
rect 2996 -1165 3196 -1127
rect 3254 -1093 3454 -1055
rect 3254 -1127 3270 -1093
rect 3438 -1127 3454 -1093
rect 3254 -1165 3454 -1127
rect 3512 -1093 3712 -1055
rect 3512 -1127 3528 -1093
rect 3696 -1127 3712 -1093
rect 3512 -1165 3712 -1127
rect 3770 -1093 3970 -1055
rect 3770 -1127 3786 -1093
rect 3954 -1127 3970 -1093
rect 3770 -1165 3970 -1127
rect 4028 -1093 4228 -1055
rect 4028 -1127 4044 -1093
rect 4212 -1127 4228 -1093
rect 4028 -1165 4228 -1127
rect 4286 -1093 4486 -1055
rect 4286 -1127 4302 -1093
rect 4470 -1127 4486 -1093
rect 4286 -1165 4486 -1127
rect 4544 -1093 4744 -1055
rect 4544 -1127 4560 -1093
rect 4728 -1127 4744 -1093
rect 4544 -1165 4744 -1127
rect 4802 -1093 5002 -1055
rect 4802 -1127 4818 -1093
rect 4986 -1127 5002 -1093
rect 4802 -1165 5002 -1127
rect 5060 -1093 5260 -1055
rect 5060 -1127 5076 -1093
rect 5244 -1127 5260 -1093
rect 5060 -1165 5260 -1127
rect 5318 -1093 5518 -1055
rect 5318 -1127 5334 -1093
rect 5502 -1127 5518 -1093
rect 5318 -1165 5518 -1127
rect 5576 -1093 5776 -1055
rect 5576 -1127 5592 -1093
rect 5760 -1127 5776 -1093
rect 5576 -1165 5776 -1127
rect 5834 -1093 6034 -1055
rect 5834 -1127 5850 -1093
rect 6018 -1127 6034 -1093
rect 5834 -1165 6034 -1127
rect 6092 -1093 6292 -1055
rect 6092 -1127 6108 -1093
rect 6276 -1127 6292 -1093
rect 6092 -1165 6292 -1127
rect 6350 -1093 6550 -1055
rect 6350 -1127 6366 -1093
rect 6534 -1127 6550 -1093
rect 6350 -1165 6550 -1127
rect 6608 -1093 6808 -1055
rect 6608 -1127 6624 -1093
rect 6792 -1127 6808 -1093
rect 6608 -1165 6808 -1127
rect 6866 -1093 7066 -1055
rect 6866 -1127 6882 -1093
rect 7050 -1127 7066 -1093
rect 6866 -1165 7066 -1127
rect -7066 -2203 -6866 -2165
rect -7066 -2237 -7050 -2203
rect -6882 -2237 -6866 -2203
rect -7066 -2253 -6866 -2237
rect -6808 -2203 -6608 -2165
rect -6808 -2237 -6792 -2203
rect -6624 -2237 -6608 -2203
rect -6808 -2253 -6608 -2237
rect -6550 -2203 -6350 -2165
rect -6550 -2237 -6534 -2203
rect -6366 -2237 -6350 -2203
rect -6550 -2253 -6350 -2237
rect -6292 -2203 -6092 -2165
rect -6292 -2237 -6276 -2203
rect -6108 -2237 -6092 -2203
rect -6292 -2253 -6092 -2237
rect -6034 -2203 -5834 -2165
rect -6034 -2237 -6018 -2203
rect -5850 -2237 -5834 -2203
rect -6034 -2253 -5834 -2237
rect -5776 -2203 -5576 -2165
rect -5776 -2237 -5760 -2203
rect -5592 -2237 -5576 -2203
rect -5776 -2253 -5576 -2237
rect -5518 -2203 -5318 -2165
rect -5518 -2237 -5502 -2203
rect -5334 -2237 -5318 -2203
rect -5518 -2253 -5318 -2237
rect -5260 -2203 -5060 -2165
rect -5260 -2237 -5244 -2203
rect -5076 -2237 -5060 -2203
rect -5260 -2253 -5060 -2237
rect -5002 -2203 -4802 -2165
rect -5002 -2237 -4986 -2203
rect -4818 -2237 -4802 -2203
rect -5002 -2253 -4802 -2237
rect -4744 -2203 -4544 -2165
rect -4744 -2237 -4728 -2203
rect -4560 -2237 -4544 -2203
rect -4744 -2253 -4544 -2237
rect -4486 -2203 -4286 -2165
rect -4486 -2237 -4470 -2203
rect -4302 -2237 -4286 -2203
rect -4486 -2253 -4286 -2237
rect -4228 -2203 -4028 -2165
rect -4228 -2237 -4212 -2203
rect -4044 -2237 -4028 -2203
rect -4228 -2253 -4028 -2237
rect -3970 -2203 -3770 -2165
rect -3970 -2237 -3954 -2203
rect -3786 -2237 -3770 -2203
rect -3970 -2253 -3770 -2237
rect -3712 -2203 -3512 -2165
rect -3712 -2237 -3696 -2203
rect -3528 -2237 -3512 -2203
rect -3712 -2253 -3512 -2237
rect -3454 -2203 -3254 -2165
rect -3454 -2237 -3438 -2203
rect -3270 -2237 -3254 -2203
rect -3454 -2253 -3254 -2237
rect -3196 -2203 -2996 -2165
rect -3196 -2237 -3180 -2203
rect -3012 -2237 -2996 -2203
rect -3196 -2253 -2996 -2237
rect -2938 -2203 -2738 -2165
rect -2938 -2237 -2922 -2203
rect -2754 -2237 -2738 -2203
rect -2938 -2253 -2738 -2237
rect -2680 -2203 -2480 -2165
rect -2680 -2237 -2664 -2203
rect -2496 -2237 -2480 -2203
rect -2680 -2253 -2480 -2237
rect -2422 -2203 -2222 -2165
rect -2422 -2237 -2406 -2203
rect -2238 -2237 -2222 -2203
rect -2422 -2253 -2222 -2237
rect -2164 -2203 -1964 -2165
rect -2164 -2237 -2148 -2203
rect -1980 -2237 -1964 -2203
rect -2164 -2253 -1964 -2237
rect -1906 -2203 -1706 -2165
rect -1906 -2237 -1890 -2203
rect -1722 -2237 -1706 -2203
rect -1906 -2253 -1706 -2237
rect -1648 -2203 -1448 -2165
rect -1648 -2237 -1632 -2203
rect -1464 -2237 -1448 -2203
rect -1648 -2253 -1448 -2237
rect -1390 -2203 -1190 -2165
rect -1390 -2237 -1374 -2203
rect -1206 -2237 -1190 -2203
rect -1390 -2253 -1190 -2237
rect -1132 -2203 -932 -2165
rect -1132 -2237 -1116 -2203
rect -948 -2237 -932 -2203
rect -1132 -2253 -932 -2237
rect -874 -2203 -674 -2165
rect -874 -2237 -858 -2203
rect -690 -2237 -674 -2203
rect -874 -2253 -674 -2237
rect -616 -2203 -416 -2165
rect -616 -2237 -600 -2203
rect -432 -2237 -416 -2203
rect -616 -2253 -416 -2237
rect -358 -2203 -158 -2165
rect -358 -2237 -342 -2203
rect -174 -2237 -158 -2203
rect -358 -2253 -158 -2237
rect -100 -2203 100 -2165
rect -100 -2237 -84 -2203
rect 84 -2237 100 -2203
rect -100 -2253 100 -2237
rect 158 -2203 358 -2165
rect 158 -2237 174 -2203
rect 342 -2237 358 -2203
rect 158 -2253 358 -2237
rect 416 -2203 616 -2165
rect 416 -2237 432 -2203
rect 600 -2237 616 -2203
rect 416 -2253 616 -2237
rect 674 -2203 874 -2165
rect 674 -2237 690 -2203
rect 858 -2237 874 -2203
rect 674 -2253 874 -2237
rect 932 -2203 1132 -2165
rect 932 -2237 948 -2203
rect 1116 -2237 1132 -2203
rect 932 -2253 1132 -2237
rect 1190 -2203 1390 -2165
rect 1190 -2237 1206 -2203
rect 1374 -2237 1390 -2203
rect 1190 -2253 1390 -2237
rect 1448 -2203 1648 -2165
rect 1448 -2237 1464 -2203
rect 1632 -2237 1648 -2203
rect 1448 -2253 1648 -2237
rect 1706 -2203 1906 -2165
rect 1706 -2237 1722 -2203
rect 1890 -2237 1906 -2203
rect 1706 -2253 1906 -2237
rect 1964 -2203 2164 -2165
rect 1964 -2237 1980 -2203
rect 2148 -2237 2164 -2203
rect 1964 -2253 2164 -2237
rect 2222 -2203 2422 -2165
rect 2222 -2237 2238 -2203
rect 2406 -2237 2422 -2203
rect 2222 -2253 2422 -2237
rect 2480 -2203 2680 -2165
rect 2480 -2237 2496 -2203
rect 2664 -2237 2680 -2203
rect 2480 -2253 2680 -2237
rect 2738 -2203 2938 -2165
rect 2738 -2237 2754 -2203
rect 2922 -2237 2938 -2203
rect 2738 -2253 2938 -2237
rect 2996 -2203 3196 -2165
rect 2996 -2237 3012 -2203
rect 3180 -2237 3196 -2203
rect 2996 -2253 3196 -2237
rect 3254 -2203 3454 -2165
rect 3254 -2237 3270 -2203
rect 3438 -2237 3454 -2203
rect 3254 -2253 3454 -2237
rect 3512 -2203 3712 -2165
rect 3512 -2237 3528 -2203
rect 3696 -2237 3712 -2203
rect 3512 -2253 3712 -2237
rect 3770 -2203 3970 -2165
rect 3770 -2237 3786 -2203
rect 3954 -2237 3970 -2203
rect 3770 -2253 3970 -2237
rect 4028 -2203 4228 -2165
rect 4028 -2237 4044 -2203
rect 4212 -2237 4228 -2203
rect 4028 -2253 4228 -2237
rect 4286 -2203 4486 -2165
rect 4286 -2237 4302 -2203
rect 4470 -2237 4486 -2203
rect 4286 -2253 4486 -2237
rect 4544 -2203 4744 -2165
rect 4544 -2237 4560 -2203
rect 4728 -2237 4744 -2203
rect 4544 -2253 4744 -2237
rect 4802 -2203 5002 -2165
rect 4802 -2237 4818 -2203
rect 4986 -2237 5002 -2203
rect 4802 -2253 5002 -2237
rect 5060 -2203 5260 -2165
rect 5060 -2237 5076 -2203
rect 5244 -2237 5260 -2203
rect 5060 -2253 5260 -2237
rect 5318 -2203 5518 -2165
rect 5318 -2237 5334 -2203
rect 5502 -2237 5518 -2203
rect 5318 -2253 5518 -2237
rect 5576 -2203 5776 -2165
rect 5576 -2237 5592 -2203
rect 5760 -2237 5776 -2203
rect 5576 -2253 5776 -2237
rect 5834 -2203 6034 -2165
rect 5834 -2237 5850 -2203
rect 6018 -2237 6034 -2203
rect 5834 -2253 6034 -2237
rect 6092 -2203 6292 -2165
rect 6092 -2237 6108 -2203
rect 6276 -2237 6292 -2203
rect 6092 -2253 6292 -2237
rect 6350 -2203 6550 -2165
rect 6350 -2237 6366 -2203
rect 6534 -2237 6550 -2203
rect 6350 -2253 6550 -2237
rect 6608 -2203 6808 -2165
rect 6608 -2237 6624 -2203
rect 6792 -2237 6808 -2203
rect 6608 -2253 6808 -2237
rect 6866 -2203 7066 -2165
rect 6866 -2237 6882 -2203
rect 7050 -2237 7066 -2203
rect 6866 -2253 7066 -2237
<< polycont >>
rect -7050 2203 -6882 2237
rect -6792 2203 -6624 2237
rect -6534 2203 -6366 2237
rect -6276 2203 -6108 2237
rect -6018 2203 -5850 2237
rect -5760 2203 -5592 2237
rect -5502 2203 -5334 2237
rect -5244 2203 -5076 2237
rect -4986 2203 -4818 2237
rect -4728 2203 -4560 2237
rect -4470 2203 -4302 2237
rect -4212 2203 -4044 2237
rect -3954 2203 -3786 2237
rect -3696 2203 -3528 2237
rect -3438 2203 -3270 2237
rect -3180 2203 -3012 2237
rect -2922 2203 -2754 2237
rect -2664 2203 -2496 2237
rect -2406 2203 -2238 2237
rect -2148 2203 -1980 2237
rect -1890 2203 -1722 2237
rect -1632 2203 -1464 2237
rect -1374 2203 -1206 2237
rect -1116 2203 -948 2237
rect -858 2203 -690 2237
rect -600 2203 -432 2237
rect -342 2203 -174 2237
rect -84 2203 84 2237
rect 174 2203 342 2237
rect 432 2203 600 2237
rect 690 2203 858 2237
rect 948 2203 1116 2237
rect 1206 2203 1374 2237
rect 1464 2203 1632 2237
rect 1722 2203 1890 2237
rect 1980 2203 2148 2237
rect 2238 2203 2406 2237
rect 2496 2203 2664 2237
rect 2754 2203 2922 2237
rect 3012 2203 3180 2237
rect 3270 2203 3438 2237
rect 3528 2203 3696 2237
rect 3786 2203 3954 2237
rect 4044 2203 4212 2237
rect 4302 2203 4470 2237
rect 4560 2203 4728 2237
rect 4818 2203 4986 2237
rect 5076 2203 5244 2237
rect 5334 2203 5502 2237
rect 5592 2203 5760 2237
rect 5850 2203 6018 2237
rect 6108 2203 6276 2237
rect 6366 2203 6534 2237
rect 6624 2203 6792 2237
rect 6882 2203 7050 2237
rect -7050 1093 -6882 1127
rect -6792 1093 -6624 1127
rect -6534 1093 -6366 1127
rect -6276 1093 -6108 1127
rect -6018 1093 -5850 1127
rect -5760 1093 -5592 1127
rect -5502 1093 -5334 1127
rect -5244 1093 -5076 1127
rect -4986 1093 -4818 1127
rect -4728 1093 -4560 1127
rect -4470 1093 -4302 1127
rect -4212 1093 -4044 1127
rect -3954 1093 -3786 1127
rect -3696 1093 -3528 1127
rect -3438 1093 -3270 1127
rect -3180 1093 -3012 1127
rect -2922 1093 -2754 1127
rect -2664 1093 -2496 1127
rect -2406 1093 -2238 1127
rect -2148 1093 -1980 1127
rect -1890 1093 -1722 1127
rect -1632 1093 -1464 1127
rect -1374 1093 -1206 1127
rect -1116 1093 -948 1127
rect -858 1093 -690 1127
rect -600 1093 -432 1127
rect -342 1093 -174 1127
rect -84 1093 84 1127
rect 174 1093 342 1127
rect 432 1093 600 1127
rect 690 1093 858 1127
rect 948 1093 1116 1127
rect 1206 1093 1374 1127
rect 1464 1093 1632 1127
rect 1722 1093 1890 1127
rect 1980 1093 2148 1127
rect 2238 1093 2406 1127
rect 2496 1093 2664 1127
rect 2754 1093 2922 1127
rect 3012 1093 3180 1127
rect 3270 1093 3438 1127
rect 3528 1093 3696 1127
rect 3786 1093 3954 1127
rect 4044 1093 4212 1127
rect 4302 1093 4470 1127
rect 4560 1093 4728 1127
rect 4818 1093 4986 1127
rect 5076 1093 5244 1127
rect 5334 1093 5502 1127
rect 5592 1093 5760 1127
rect 5850 1093 6018 1127
rect 6108 1093 6276 1127
rect 6366 1093 6534 1127
rect 6624 1093 6792 1127
rect 6882 1093 7050 1127
rect -7050 -17 -6882 17
rect -6792 -17 -6624 17
rect -6534 -17 -6366 17
rect -6276 -17 -6108 17
rect -6018 -17 -5850 17
rect -5760 -17 -5592 17
rect -5502 -17 -5334 17
rect -5244 -17 -5076 17
rect -4986 -17 -4818 17
rect -4728 -17 -4560 17
rect -4470 -17 -4302 17
rect -4212 -17 -4044 17
rect -3954 -17 -3786 17
rect -3696 -17 -3528 17
rect -3438 -17 -3270 17
rect -3180 -17 -3012 17
rect -2922 -17 -2754 17
rect -2664 -17 -2496 17
rect -2406 -17 -2238 17
rect -2148 -17 -1980 17
rect -1890 -17 -1722 17
rect -1632 -17 -1464 17
rect -1374 -17 -1206 17
rect -1116 -17 -948 17
rect -858 -17 -690 17
rect -600 -17 -432 17
rect -342 -17 -174 17
rect -84 -17 84 17
rect 174 -17 342 17
rect 432 -17 600 17
rect 690 -17 858 17
rect 948 -17 1116 17
rect 1206 -17 1374 17
rect 1464 -17 1632 17
rect 1722 -17 1890 17
rect 1980 -17 2148 17
rect 2238 -17 2406 17
rect 2496 -17 2664 17
rect 2754 -17 2922 17
rect 3012 -17 3180 17
rect 3270 -17 3438 17
rect 3528 -17 3696 17
rect 3786 -17 3954 17
rect 4044 -17 4212 17
rect 4302 -17 4470 17
rect 4560 -17 4728 17
rect 4818 -17 4986 17
rect 5076 -17 5244 17
rect 5334 -17 5502 17
rect 5592 -17 5760 17
rect 5850 -17 6018 17
rect 6108 -17 6276 17
rect 6366 -17 6534 17
rect 6624 -17 6792 17
rect 6882 -17 7050 17
rect -7050 -1127 -6882 -1093
rect -6792 -1127 -6624 -1093
rect -6534 -1127 -6366 -1093
rect -6276 -1127 -6108 -1093
rect -6018 -1127 -5850 -1093
rect -5760 -1127 -5592 -1093
rect -5502 -1127 -5334 -1093
rect -5244 -1127 -5076 -1093
rect -4986 -1127 -4818 -1093
rect -4728 -1127 -4560 -1093
rect -4470 -1127 -4302 -1093
rect -4212 -1127 -4044 -1093
rect -3954 -1127 -3786 -1093
rect -3696 -1127 -3528 -1093
rect -3438 -1127 -3270 -1093
rect -3180 -1127 -3012 -1093
rect -2922 -1127 -2754 -1093
rect -2664 -1127 -2496 -1093
rect -2406 -1127 -2238 -1093
rect -2148 -1127 -1980 -1093
rect -1890 -1127 -1722 -1093
rect -1632 -1127 -1464 -1093
rect -1374 -1127 -1206 -1093
rect -1116 -1127 -948 -1093
rect -858 -1127 -690 -1093
rect -600 -1127 -432 -1093
rect -342 -1127 -174 -1093
rect -84 -1127 84 -1093
rect 174 -1127 342 -1093
rect 432 -1127 600 -1093
rect 690 -1127 858 -1093
rect 948 -1127 1116 -1093
rect 1206 -1127 1374 -1093
rect 1464 -1127 1632 -1093
rect 1722 -1127 1890 -1093
rect 1980 -1127 2148 -1093
rect 2238 -1127 2406 -1093
rect 2496 -1127 2664 -1093
rect 2754 -1127 2922 -1093
rect 3012 -1127 3180 -1093
rect 3270 -1127 3438 -1093
rect 3528 -1127 3696 -1093
rect 3786 -1127 3954 -1093
rect 4044 -1127 4212 -1093
rect 4302 -1127 4470 -1093
rect 4560 -1127 4728 -1093
rect 4818 -1127 4986 -1093
rect 5076 -1127 5244 -1093
rect 5334 -1127 5502 -1093
rect 5592 -1127 5760 -1093
rect 5850 -1127 6018 -1093
rect 6108 -1127 6276 -1093
rect 6366 -1127 6534 -1093
rect 6624 -1127 6792 -1093
rect 6882 -1127 7050 -1093
rect -7050 -2237 -6882 -2203
rect -6792 -2237 -6624 -2203
rect -6534 -2237 -6366 -2203
rect -6276 -2237 -6108 -2203
rect -6018 -2237 -5850 -2203
rect -5760 -2237 -5592 -2203
rect -5502 -2237 -5334 -2203
rect -5244 -2237 -5076 -2203
rect -4986 -2237 -4818 -2203
rect -4728 -2237 -4560 -2203
rect -4470 -2237 -4302 -2203
rect -4212 -2237 -4044 -2203
rect -3954 -2237 -3786 -2203
rect -3696 -2237 -3528 -2203
rect -3438 -2237 -3270 -2203
rect -3180 -2237 -3012 -2203
rect -2922 -2237 -2754 -2203
rect -2664 -2237 -2496 -2203
rect -2406 -2237 -2238 -2203
rect -2148 -2237 -1980 -2203
rect -1890 -2237 -1722 -2203
rect -1632 -2237 -1464 -2203
rect -1374 -2237 -1206 -2203
rect -1116 -2237 -948 -2203
rect -858 -2237 -690 -2203
rect -600 -2237 -432 -2203
rect -342 -2237 -174 -2203
rect -84 -2237 84 -2203
rect 174 -2237 342 -2203
rect 432 -2237 600 -2203
rect 690 -2237 858 -2203
rect 948 -2237 1116 -2203
rect 1206 -2237 1374 -2203
rect 1464 -2237 1632 -2203
rect 1722 -2237 1890 -2203
rect 1980 -2237 2148 -2203
rect 2238 -2237 2406 -2203
rect 2496 -2237 2664 -2203
rect 2754 -2237 2922 -2203
rect 3012 -2237 3180 -2203
rect 3270 -2237 3438 -2203
rect 3528 -2237 3696 -2203
rect 3786 -2237 3954 -2203
rect 4044 -2237 4212 -2203
rect 4302 -2237 4470 -2203
rect 4560 -2237 4728 -2203
rect 4818 -2237 4986 -2203
rect 5076 -2237 5244 -2203
rect 5334 -2237 5502 -2203
rect 5592 -2237 5760 -2203
rect 5850 -2237 6018 -2203
rect 6108 -2237 6276 -2203
rect 6366 -2237 6534 -2203
rect 6624 -2237 6792 -2203
rect 6882 -2237 7050 -2203
<< locali >>
rect -7246 2341 -7150 2375
rect 7150 2341 7246 2375
rect -7246 2279 -7212 2341
rect 7212 2279 7246 2341
rect -7066 2203 -7050 2237
rect -6882 2203 -6866 2237
rect -6808 2203 -6792 2237
rect -6624 2203 -6608 2237
rect -6550 2203 -6534 2237
rect -6366 2203 -6350 2237
rect -6292 2203 -6276 2237
rect -6108 2203 -6092 2237
rect -6034 2203 -6018 2237
rect -5850 2203 -5834 2237
rect -5776 2203 -5760 2237
rect -5592 2203 -5576 2237
rect -5518 2203 -5502 2237
rect -5334 2203 -5318 2237
rect -5260 2203 -5244 2237
rect -5076 2203 -5060 2237
rect -5002 2203 -4986 2237
rect -4818 2203 -4802 2237
rect -4744 2203 -4728 2237
rect -4560 2203 -4544 2237
rect -4486 2203 -4470 2237
rect -4302 2203 -4286 2237
rect -4228 2203 -4212 2237
rect -4044 2203 -4028 2237
rect -3970 2203 -3954 2237
rect -3786 2203 -3770 2237
rect -3712 2203 -3696 2237
rect -3528 2203 -3512 2237
rect -3454 2203 -3438 2237
rect -3270 2203 -3254 2237
rect -3196 2203 -3180 2237
rect -3012 2203 -2996 2237
rect -2938 2203 -2922 2237
rect -2754 2203 -2738 2237
rect -2680 2203 -2664 2237
rect -2496 2203 -2480 2237
rect -2422 2203 -2406 2237
rect -2238 2203 -2222 2237
rect -2164 2203 -2148 2237
rect -1980 2203 -1964 2237
rect -1906 2203 -1890 2237
rect -1722 2203 -1706 2237
rect -1648 2203 -1632 2237
rect -1464 2203 -1448 2237
rect -1390 2203 -1374 2237
rect -1206 2203 -1190 2237
rect -1132 2203 -1116 2237
rect -948 2203 -932 2237
rect -874 2203 -858 2237
rect -690 2203 -674 2237
rect -616 2203 -600 2237
rect -432 2203 -416 2237
rect -358 2203 -342 2237
rect -174 2203 -158 2237
rect -100 2203 -84 2237
rect 84 2203 100 2237
rect 158 2203 174 2237
rect 342 2203 358 2237
rect 416 2203 432 2237
rect 600 2203 616 2237
rect 674 2203 690 2237
rect 858 2203 874 2237
rect 932 2203 948 2237
rect 1116 2203 1132 2237
rect 1190 2203 1206 2237
rect 1374 2203 1390 2237
rect 1448 2203 1464 2237
rect 1632 2203 1648 2237
rect 1706 2203 1722 2237
rect 1890 2203 1906 2237
rect 1964 2203 1980 2237
rect 2148 2203 2164 2237
rect 2222 2203 2238 2237
rect 2406 2203 2422 2237
rect 2480 2203 2496 2237
rect 2664 2203 2680 2237
rect 2738 2203 2754 2237
rect 2922 2203 2938 2237
rect 2996 2203 3012 2237
rect 3180 2203 3196 2237
rect 3254 2203 3270 2237
rect 3438 2203 3454 2237
rect 3512 2203 3528 2237
rect 3696 2203 3712 2237
rect 3770 2203 3786 2237
rect 3954 2203 3970 2237
rect 4028 2203 4044 2237
rect 4212 2203 4228 2237
rect 4286 2203 4302 2237
rect 4470 2203 4486 2237
rect 4544 2203 4560 2237
rect 4728 2203 4744 2237
rect 4802 2203 4818 2237
rect 4986 2203 5002 2237
rect 5060 2203 5076 2237
rect 5244 2203 5260 2237
rect 5318 2203 5334 2237
rect 5502 2203 5518 2237
rect 5576 2203 5592 2237
rect 5760 2203 5776 2237
rect 5834 2203 5850 2237
rect 6018 2203 6034 2237
rect 6092 2203 6108 2237
rect 6276 2203 6292 2237
rect 6350 2203 6366 2237
rect 6534 2203 6550 2237
rect 6608 2203 6624 2237
rect 6792 2203 6808 2237
rect 6866 2203 6882 2237
rect 7050 2203 7066 2237
rect -7112 2153 -7078 2169
rect -7112 1161 -7078 1177
rect -6854 2153 -6820 2169
rect -6854 1161 -6820 1177
rect -6596 2153 -6562 2169
rect -6596 1161 -6562 1177
rect -6338 2153 -6304 2169
rect -6338 1161 -6304 1177
rect -6080 2153 -6046 2169
rect -6080 1161 -6046 1177
rect -5822 2153 -5788 2169
rect -5822 1161 -5788 1177
rect -5564 2153 -5530 2169
rect -5564 1161 -5530 1177
rect -5306 2153 -5272 2169
rect -5306 1161 -5272 1177
rect -5048 2153 -5014 2169
rect -5048 1161 -5014 1177
rect -4790 2153 -4756 2169
rect -4790 1161 -4756 1177
rect -4532 2153 -4498 2169
rect -4532 1161 -4498 1177
rect -4274 2153 -4240 2169
rect -4274 1161 -4240 1177
rect -4016 2153 -3982 2169
rect -4016 1161 -3982 1177
rect -3758 2153 -3724 2169
rect -3758 1161 -3724 1177
rect -3500 2153 -3466 2169
rect -3500 1161 -3466 1177
rect -3242 2153 -3208 2169
rect -3242 1161 -3208 1177
rect -2984 2153 -2950 2169
rect -2984 1161 -2950 1177
rect -2726 2153 -2692 2169
rect -2726 1161 -2692 1177
rect -2468 2153 -2434 2169
rect -2468 1161 -2434 1177
rect -2210 2153 -2176 2169
rect -2210 1161 -2176 1177
rect -1952 2153 -1918 2169
rect -1952 1161 -1918 1177
rect -1694 2153 -1660 2169
rect -1694 1161 -1660 1177
rect -1436 2153 -1402 2169
rect -1436 1161 -1402 1177
rect -1178 2153 -1144 2169
rect -1178 1161 -1144 1177
rect -920 2153 -886 2169
rect -920 1161 -886 1177
rect -662 2153 -628 2169
rect -662 1161 -628 1177
rect -404 2153 -370 2169
rect -404 1161 -370 1177
rect -146 2153 -112 2169
rect -146 1161 -112 1177
rect 112 2153 146 2169
rect 112 1161 146 1177
rect 370 2153 404 2169
rect 370 1161 404 1177
rect 628 2153 662 2169
rect 628 1161 662 1177
rect 886 2153 920 2169
rect 886 1161 920 1177
rect 1144 2153 1178 2169
rect 1144 1161 1178 1177
rect 1402 2153 1436 2169
rect 1402 1161 1436 1177
rect 1660 2153 1694 2169
rect 1660 1161 1694 1177
rect 1918 2153 1952 2169
rect 1918 1161 1952 1177
rect 2176 2153 2210 2169
rect 2176 1161 2210 1177
rect 2434 2153 2468 2169
rect 2434 1161 2468 1177
rect 2692 2153 2726 2169
rect 2692 1161 2726 1177
rect 2950 2153 2984 2169
rect 2950 1161 2984 1177
rect 3208 2153 3242 2169
rect 3208 1161 3242 1177
rect 3466 2153 3500 2169
rect 3466 1161 3500 1177
rect 3724 2153 3758 2169
rect 3724 1161 3758 1177
rect 3982 2153 4016 2169
rect 3982 1161 4016 1177
rect 4240 2153 4274 2169
rect 4240 1161 4274 1177
rect 4498 2153 4532 2169
rect 4498 1161 4532 1177
rect 4756 2153 4790 2169
rect 4756 1161 4790 1177
rect 5014 2153 5048 2169
rect 5014 1161 5048 1177
rect 5272 2153 5306 2169
rect 5272 1161 5306 1177
rect 5530 2153 5564 2169
rect 5530 1161 5564 1177
rect 5788 2153 5822 2169
rect 5788 1161 5822 1177
rect 6046 2153 6080 2169
rect 6046 1161 6080 1177
rect 6304 2153 6338 2169
rect 6304 1161 6338 1177
rect 6562 2153 6596 2169
rect 6562 1161 6596 1177
rect 6820 2153 6854 2169
rect 6820 1161 6854 1177
rect 7078 2153 7112 2169
rect 7078 1161 7112 1177
rect -7066 1093 -7050 1127
rect -6882 1093 -6866 1127
rect -6808 1093 -6792 1127
rect -6624 1093 -6608 1127
rect -6550 1093 -6534 1127
rect -6366 1093 -6350 1127
rect -6292 1093 -6276 1127
rect -6108 1093 -6092 1127
rect -6034 1093 -6018 1127
rect -5850 1093 -5834 1127
rect -5776 1093 -5760 1127
rect -5592 1093 -5576 1127
rect -5518 1093 -5502 1127
rect -5334 1093 -5318 1127
rect -5260 1093 -5244 1127
rect -5076 1093 -5060 1127
rect -5002 1093 -4986 1127
rect -4818 1093 -4802 1127
rect -4744 1093 -4728 1127
rect -4560 1093 -4544 1127
rect -4486 1093 -4470 1127
rect -4302 1093 -4286 1127
rect -4228 1093 -4212 1127
rect -4044 1093 -4028 1127
rect -3970 1093 -3954 1127
rect -3786 1093 -3770 1127
rect -3712 1093 -3696 1127
rect -3528 1093 -3512 1127
rect -3454 1093 -3438 1127
rect -3270 1093 -3254 1127
rect -3196 1093 -3180 1127
rect -3012 1093 -2996 1127
rect -2938 1093 -2922 1127
rect -2754 1093 -2738 1127
rect -2680 1093 -2664 1127
rect -2496 1093 -2480 1127
rect -2422 1093 -2406 1127
rect -2238 1093 -2222 1127
rect -2164 1093 -2148 1127
rect -1980 1093 -1964 1127
rect -1906 1093 -1890 1127
rect -1722 1093 -1706 1127
rect -1648 1093 -1632 1127
rect -1464 1093 -1448 1127
rect -1390 1093 -1374 1127
rect -1206 1093 -1190 1127
rect -1132 1093 -1116 1127
rect -948 1093 -932 1127
rect -874 1093 -858 1127
rect -690 1093 -674 1127
rect -616 1093 -600 1127
rect -432 1093 -416 1127
rect -358 1093 -342 1127
rect -174 1093 -158 1127
rect -100 1093 -84 1127
rect 84 1093 100 1127
rect 158 1093 174 1127
rect 342 1093 358 1127
rect 416 1093 432 1127
rect 600 1093 616 1127
rect 674 1093 690 1127
rect 858 1093 874 1127
rect 932 1093 948 1127
rect 1116 1093 1132 1127
rect 1190 1093 1206 1127
rect 1374 1093 1390 1127
rect 1448 1093 1464 1127
rect 1632 1093 1648 1127
rect 1706 1093 1722 1127
rect 1890 1093 1906 1127
rect 1964 1093 1980 1127
rect 2148 1093 2164 1127
rect 2222 1093 2238 1127
rect 2406 1093 2422 1127
rect 2480 1093 2496 1127
rect 2664 1093 2680 1127
rect 2738 1093 2754 1127
rect 2922 1093 2938 1127
rect 2996 1093 3012 1127
rect 3180 1093 3196 1127
rect 3254 1093 3270 1127
rect 3438 1093 3454 1127
rect 3512 1093 3528 1127
rect 3696 1093 3712 1127
rect 3770 1093 3786 1127
rect 3954 1093 3970 1127
rect 4028 1093 4044 1127
rect 4212 1093 4228 1127
rect 4286 1093 4302 1127
rect 4470 1093 4486 1127
rect 4544 1093 4560 1127
rect 4728 1093 4744 1127
rect 4802 1093 4818 1127
rect 4986 1093 5002 1127
rect 5060 1093 5076 1127
rect 5244 1093 5260 1127
rect 5318 1093 5334 1127
rect 5502 1093 5518 1127
rect 5576 1093 5592 1127
rect 5760 1093 5776 1127
rect 5834 1093 5850 1127
rect 6018 1093 6034 1127
rect 6092 1093 6108 1127
rect 6276 1093 6292 1127
rect 6350 1093 6366 1127
rect 6534 1093 6550 1127
rect 6608 1093 6624 1127
rect 6792 1093 6808 1127
rect 6866 1093 6882 1127
rect 7050 1093 7066 1127
rect -7112 1043 -7078 1059
rect -7112 51 -7078 67
rect -6854 1043 -6820 1059
rect -6854 51 -6820 67
rect -6596 1043 -6562 1059
rect -6596 51 -6562 67
rect -6338 1043 -6304 1059
rect -6338 51 -6304 67
rect -6080 1043 -6046 1059
rect -6080 51 -6046 67
rect -5822 1043 -5788 1059
rect -5822 51 -5788 67
rect -5564 1043 -5530 1059
rect -5564 51 -5530 67
rect -5306 1043 -5272 1059
rect -5306 51 -5272 67
rect -5048 1043 -5014 1059
rect -5048 51 -5014 67
rect -4790 1043 -4756 1059
rect -4790 51 -4756 67
rect -4532 1043 -4498 1059
rect -4532 51 -4498 67
rect -4274 1043 -4240 1059
rect -4274 51 -4240 67
rect -4016 1043 -3982 1059
rect -4016 51 -3982 67
rect -3758 1043 -3724 1059
rect -3758 51 -3724 67
rect -3500 1043 -3466 1059
rect -3500 51 -3466 67
rect -3242 1043 -3208 1059
rect -3242 51 -3208 67
rect -2984 1043 -2950 1059
rect -2984 51 -2950 67
rect -2726 1043 -2692 1059
rect -2726 51 -2692 67
rect -2468 1043 -2434 1059
rect -2468 51 -2434 67
rect -2210 1043 -2176 1059
rect -2210 51 -2176 67
rect -1952 1043 -1918 1059
rect -1952 51 -1918 67
rect -1694 1043 -1660 1059
rect -1694 51 -1660 67
rect -1436 1043 -1402 1059
rect -1436 51 -1402 67
rect -1178 1043 -1144 1059
rect -1178 51 -1144 67
rect -920 1043 -886 1059
rect -920 51 -886 67
rect -662 1043 -628 1059
rect -662 51 -628 67
rect -404 1043 -370 1059
rect -404 51 -370 67
rect -146 1043 -112 1059
rect -146 51 -112 67
rect 112 1043 146 1059
rect 112 51 146 67
rect 370 1043 404 1059
rect 370 51 404 67
rect 628 1043 662 1059
rect 628 51 662 67
rect 886 1043 920 1059
rect 886 51 920 67
rect 1144 1043 1178 1059
rect 1144 51 1178 67
rect 1402 1043 1436 1059
rect 1402 51 1436 67
rect 1660 1043 1694 1059
rect 1660 51 1694 67
rect 1918 1043 1952 1059
rect 1918 51 1952 67
rect 2176 1043 2210 1059
rect 2176 51 2210 67
rect 2434 1043 2468 1059
rect 2434 51 2468 67
rect 2692 1043 2726 1059
rect 2692 51 2726 67
rect 2950 1043 2984 1059
rect 2950 51 2984 67
rect 3208 1043 3242 1059
rect 3208 51 3242 67
rect 3466 1043 3500 1059
rect 3466 51 3500 67
rect 3724 1043 3758 1059
rect 3724 51 3758 67
rect 3982 1043 4016 1059
rect 3982 51 4016 67
rect 4240 1043 4274 1059
rect 4240 51 4274 67
rect 4498 1043 4532 1059
rect 4498 51 4532 67
rect 4756 1043 4790 1059
rect 4756 51 4790 67
rect 5014 1043 5048 1059
rect 5014 51 5048 67
rect 5272 1043 5306 1059
rect 5272 51 5306 67
rect 5530 1043 5564 1059
rect 5530 51 5564 67
rect 5788 1043 5822 1059
rect 5788 51 5822 67
rect 6046 1043 6080 1059
rect 6046 51 6080 67
rect 6304 1043 6338 1059
rect 6304 51 6338 67
rect 6562 1043 6596 1059
rect 6562 51 6596 67
rect 6820 1043 6854 1059
rect 6820 51 6854 67
rect 7078 1043 7112 1059
rect 7078 51 7112 67
rect -7066 -17 -7050 17
rect -6882 -17 -6866 17
rect -6808 -17 -6792 17
rect -6624 -17 -6608 17
rect -6550 -17 -6534 17
rect -6366 -17 -6350 17
rect -6292 -17 -6276 17
rect -6108 -17 -6092 17
rect -6034 -17 -6018 17
rect -5850 -17 -5834 17
rect -5776 -17 -5760 17
rect -5592 -17 -5576 17
rect -5518 -17 -5502 17
rect -5334 -17 -5318 17
rect -5260 -17 -5244 17
rect -5076 -17 -5060 17
rect -5002 -17 -4986 17
rect -4818 -17 -4802 17
rect -4744 -17 -4728 17
rect -4560 -17 -4544 17
rect -4486 -17 -4470 17
rect -4302 -17 -4286 17
rect -4228 -17 -4212 17
rect -4044 -17 -4028 17
rect -3970 -17 -3954 17
rect -3786 -17 -3770 17
rect -3712 -17 -3696 17
rect -3528 -17 -3512 17
rect -3454 -17 -3438 17
rect -3270 -17 -3254 17
rect -3196 -17 -3180 17
rect -3012 -17 -2996 17
rect -2938 -17 -2922 17
rect -2754 -17 -2738 17
rect -2680 -17 -2664 17
rect -2496 -17 -2480 17
rect -2422 -17 -2406 17
rect -2238 -17 -2222 17
rect -2164 -17 -2148 17
rect -1980 -17 -1964 17
rect -1906 -17 -1890 17
rect -1722 -17 -1706 17
rect -1648 -17 -1632 17
rect -1464 -17 -1448 17
rect -1390 -17 -1374 17
rect -1206 -17 -1190 17
rect -1132 -17 -1116 17
rect -948 -17 -932 17
rect -874 -17 -858 17
rect -690 -17 -674 17
rect -616 -17 -600 17
rect -432 -17 -416 17
rect -358 -17 -342 17
rect -174 -17 -158 17
rect -100 -17 -84 17
rect 84 -17 100 17
rect 158 -17 174 17
rect 342 -17 358 17
rect 416 -17 432 17
rect 600 -17 616 17
rect 674 -17 690 17
rect 858 -17 874 17
rect 932 -17 948 17
rect 1116 -17 1132 17
rect 1190 -17 1206 17
rect 1374 -17 1390 17
rect 1448 -17 1464 17
rect 1632 -17 1648 17
rect 1706 -17 1722 17
rect 1890 -17 1906 17
rect 1964 -17 1980 17
rect 2148 -17 2164 17
rect 2222 -17 2238 17
rect 2406 -17 2422 17
rect 2480 -17 2496 17
rect 2664 -17 2680 17
rect 2738 -17 2754 17
rect 2922 -17 2938 17
rect 2996 -17 3012 17
rect 3180 -17 3196 17
rect 3254 -17 3270 17
rect 3438 -17 3454 17
rect 3512 -17 3528 17
rect 3696 -17 3712 17
rect 3770 -17 3786 17
rect 3954 -17 3970 17
rect 4028 -17 4044 17
rect 4212 -17 4228 17
rect 4286 -17 4302 17
rect 4470 -17 4486 17
rect 4544 -17 4560 17
rect 4728 -17 4744 17
rect 4802 -17 4818 17
rect 4986 -17 5002 17
rect 5060 -17 5076 17
rect 5244 -17 5260 17
rect 5318 -17 5334 17
rect 5502 -17 5518 17
rect 5576 -17 5592 17
rect 5760 -17 5776 17
rect 5834 -17 5850 17
rect 6018 -17 6034 17
rect 6092 -17 6108 17
rect 6276 -17 6292 17
rect 6350 -17 6366 17
rect 6534 -17 6550 17
rect 6608 -17 6624 17
rect 6792 -17 6808 17
rect 6866 -17 6882 17
rect 7050 -17 7066 17
rect -7112 -67 -7078 -51
rect -7112 -1059 -7078 -1043
rect -6854 -67 -6820 -51
rect -6854 -1059 -6820 -1043
rect -6596 -67 -6562 -51
rect -6596 -1059 -6562 -1043
rect -6338 -67 -6304 -51
rect -6338 -1059 -6304 -1043
rect -6080 -67 -6046 -51
rect -6080 -1059 -6046 -1043
rect -5822 -67 -5788 -51
rect -5822 -1059 -5788 -1043
rect -5564 -67 -5530 -51
rect -5564 -1059 -5530 -1043
rect -5306 -67 -5272 -51
rect -5306 -1059 -5272 -1043
rect -5048 -67 -5014 -51
rect -5048 -1059 -5014 -1043
rect -4790 -67 -4756 -51
rect -4790 -1059 -4756 -1043
rect -4532 -67 -4498 -51
rect -4532 -1059 -4498 -1043
rect -4274 -67 -4240 -51
rect -4274 -1059 -4240 -1043
rect -4016 -67 -3982 -51
rect -4016 -1059 -3982 -1043
rect -3758 -67 -3724 -51
rect -3758 -1059 -3724 -1043
rect -3500 -67 -3466 -51
rect -3500 -1059 -3466 -1043
rect -3242 -67 -3208 -51
rect -3242 -1059 -3208 -1043
rect -2984 -67 -2950 -51
rect -2984 -1059 -2950 -1043
rect -2726 -67 -2692 -51
rect -2726 -1059 -2692 -1043
rect -2468 -67 -2434 -51
rect -2468 -1059 -2434 -1043
rect -2210 -67 -2176 -51
rect -2210 -1059 -2176 -1043
rect -1952 -67 -1918 -51
rect -1952 -1059 -1918 -1043
rect -1694 -67 -1660 -51
rect -1694 -1059 -1660 -1043
rect -1436 -67 -1402 -51
rect -1436 -1059 -1402 -1043
rect -1178 -67 -1144 -51
rect -1178 -1059 -1144 -1043
rect -920 -67 -886 -51
rect -920 -1059 -886 -1043
rect -662 -67 -628 -51
rect -662 -1059 -628 -1043
rect -404 -67 -370 -51
rect -404 -1059 -370 -1043
rect -146 -67 -112 -51
rect -146 -1059 -112 -1043
rect 112 -67 146 -51
rect 112 -1059 146 -1043
rect 370 -67 404 -51
rect 370 -1059 404 -1043
rect 628 -67 662 -51
rect 628 -1059 662 -1043
rect 886 -67 920 -51
rect 886 -1059 920 -1043
rect 1144 -67 1178 -51
rect 1144 -1059 1178 -1043
rect 1402 -67 1436 -51
rect 1402 -1059 1436 -1043
rect 1660 -67 1694 -51
rect 1660 -1059 1694 -1043
rect 1918 -67 1952 -51
rect 1918 -1059 1952 -1043
rect 2176 -67 2210 -51
rect 2176 -1059 2210 -1043
rect 2434 -67 2468 -51
rect 2434 -1059 2468 -1043
rect 2692 -67 2726 -51
rect 2692 -1059 2726 -1043
rect 2950 -67 2984 -51
rect 2950 -1059 2984 -1043
rect 3208 -67 3242 -51
rect 3208 -1059 3242 -1043
rect 3466 -67 3500 -51
rect 3466 -1059 3500 -1043
rect 3724 -67 3758 -51
rect 3724 -1059 3758 -1043
rect 3982 -67 4016 -51
rect 3982 -1059 4016 -1043
rect 4240 -67 4274 -51
rect 4240 -1059 4274 -1043
rect 4498 -67 4532 -51
rect 4498 -1059 4532 -1043
rect 4756 -67 4790 -51
rect 4756 -1059 4790 -1043
rect 5014 -67 5048 -51
rect 5014 -1059 5048 -1043
rect 5272 -67 5306 -51
rect 5272 -1059 5306 -1043
rect 5530 -67 5564 -51
rect 5530 -1059 5564 -1043
rect 5788 -67 5822 -51
rect 5788 -1059 5822 -1043
rect 6046 -67 6080 -51
rect 6046 -1059 6080 -1043
rect 6304 -67 6338 -51
rect 6304 -1059 6338 -1043
rect 6562 -67 6596 -51
rect 6562 -1059 6596 -1043
rect 6820 -67 6854 -51
rect 6820 -1059 6854 -1043
rect 7078 -67 7112 -51
rect 7078 -1059 7112 -1043
rect -7066 -1127 -7050 -1093
rect -6882 -1127 -6866 -1093
rect -6808 -1127 -6792 -1093
rect -6624 -1127 -6608 -1093
rect -6550 -1127 -6534 -1093
rect -6366 -1127 -6350 -1093
rect -6292 -1127 -6276 -1093
rect -6108 -1127 -6092 -1093
rect -6034 -1127 -6018 -1093
rect -5850 -1127 -5834 -1093
rect -5776 -1127 -5760 -1093
rect -5592 -1127 -5576 -1093
rect -5518 -1127 -5502 -1093
rect -5334 -1127 -5318 -1093
rect -5260 -1127 -5244 -1093
rect -5076 -1127 -5060 -1093
rect -5002 -1127 -4986 -1093
rect -4818 -1127 -4802 -1093
rect -4744 -1127 -4728 -1093
rect -4560 -1127 -4544 -1093
rect -4486 -1127 -4470 -1093
rect -4302 -1127 -4286 -1093
rect -4228 -1127 -4212 -1093
rect -4044 -1127 -4028 -1093
rect -3970 -1127 -3954 -1093
rect -3786 -1127 -3770 -1093
rect -3712 -1127 -3696 -1093
rect -3528 -1127 -3512 -1093
rect -3454 -1127 -3438 -1093
rect -3270 -1127 -3254 -1093
rect -3196 -1127 -3180 -1093
rect -3012 -1127 -2996 -1093
rect -2938 -1127 -2922 -1093
rect -2754 -1127 -2738 -1093
rect -2680 -1127 -2664 -1093
rect -2496 -1127 -2480 -1093
rect -2422 -1127 -2406 -1093
rect -2238 -1127 -2222 -1093
rect -2164 -1127 -2148 -1093
rect -1980 -1127 -1964 -1093
rect -1906 -1127 -1890 -1093
rect -1722 -1127 -1706 -1093
rect -1648 -1127 -1632 -1093
rect -1464 -1127 -1448 -1093
rect -1390 -1127 -1374 -1093
rect -1206 -1127 -1190 -1093
rect -1132 -1127 -1116 -1093
rect -948 -1127 -932 -1093
rect -874 -1127 -858 -1093
rect -690 -1127 -674 -1093
rect -616 -1127 -600 -1093
rect -432 -1127 -416 -1093
rect -358 -1127 -342 -1093
rect -174 -1127 -158 -1093
rect -100 -1127 -84 -1093
rect 84 -1127 100 -1093
rect 158 -1127 174 -1093
rect 342 -1127 358 -1093
rect 416 -1127 432 -1093
rect 600 -1127 616 -1093
rect 674 -1127 690 -1093
rect 858 -1127 874 -1093
rect 932 -1127 948 -1093
rect 1116 -1127 1132 -1093
rect 1190 -1127 1206 -1093
rect 1374 -1127 1390 -1093
rect 1448 -1127 1464 -1093
rect 1632 -1127 1648 -1093
rect 1706 -1127 1722 -1093
rect 1890 -1127 1906 -1093
rect 1964 -1127 1980 -1093
rect 2148 -1127 2164 -1093
rect 2222 -1127 2238 -1093
rect 2406 -1127 2422 -1093
rect 2480 -1127 2496 -1093
rect 2664 -1127 2680 -1093
rect 2738 -1127 2754 -1093
rect 2922 -1127 2938 -1093
rect 2996 -1127 3012 -1093
rect 3180 -1127 3196 -1093
rect 3254 -1127 3270 -1093
rect 3438 -1127 3454 -1093
rect 3512 -1127 3528 -1093
rect 3696 -1127 3712 -1093
rect 3770 -1127 3786 -1093
rect 3954 -1127 3970 -1093
rect 4028 -1127 4044 -1093
rect 4212 -1127 4228 -1093
rect 4286 -1127 4302 -1093
rect 4470 -1127 4486 -1093
rect 4544 -1127 4560 -1093
rect 4728 -1127 4744 -1093
rect 4802 -1127 4818 -1093
rect 4986 -1127 5002 -1093
rect 5060 -1127 5076 -1093
rect 5244 -1127 5260 -1093
rect 5318 -1127 5334 -1093
rect 5502 -1127 5518 -1093
rect 5576 -1127 5592 -1093
rect 5760 -1127 5776 -1093
rect 5834 -1127 5850 -1093
rect 6018 -1127 6034 -1093
rect 6092 -1127 6108 -1093
rect 6276 -1127 6292 -1093
rect 6350 -1127 6366 -1093
rect 6534 -1127 6550 -1093
rect 6608 -1127 6624 -1093
rect 6792 -1127 6808 -1093
rect 6866 -1127 6882 -1093
rect 7050 -1127 7066 -1093
rect -7112 -1177 -7078 -1161
rect -7112 -2169 -7078 -2153
rect -6854 -1177 -6820 -1161
rect -6854 -2169 -6820 -2153
rect -6596 -1177 -6562 -1161
rect -6596 -2169 -6562 -2153
rect -6338 -1177 -6304 -1161
rect -6338 -2169 -6304 -2153
rect -6080 -1177 -6046 -1161
rect -6080 -2169 -6046 -2153
rect -5822 -1177 -5788 -1161
rect -5822 -2169 -5788 -2153
rect -5564 -1177 -5530 -1161
rect -5564 -2169 -5530 -2153
rect -5306 -1177 -5272 -1161
rect -5306 -2169 -5272 -2153
rect -5048 -1177 -5014 -1161
rect -5048 -2169 -5014 -2153
rect -4790 -1177 -4756 -1161
rect -4790 -2169 -4756 -2153
rect -4532 -1177 -4498 -1161
rect -4532 -2169 -4498 -2153
rect -4274 -1177 -4240 -1161
rect -4274 -2169 -4240 -2153
rect -4016 -1177 -3982 -1161
rect -4016 -2169 -3982 -2153
rect -3758 -1177 -3724 -1161
rect -3758 -2169 -3724 -2153
rect -3500 -1177 -3466 -1161
rect -3500 -2169 -3466 -2153
rect -3242 -1177 -3208 -1161
rect -3242 -2169 -3208 -2153
rect -2984 -1177 -2950 -1161
rect -2984 -2169 -2950 -2153
rect -2726 -1177 -2692 -1161
rect -2726 -2169 -2692 -2153
rect -2468 -1177 -2434 -1161
rect -2468 -2169 -2434 -2153
rect -2210 -1177 -2176 -1161
rect -2210 -2169 -2176 -2153
rect -1952 -1177 -1918 -1161
rect -1952 -2169 -1918 -2153
rect -1694 -1177 -1660 -1161
rect -1694 -2169 -1660 -2153
rect -1436 -1177 -1402 -1161
rect -1436 -2169 -1402 -2153
rect -1178 -1177 -1144 -1161
rect -1178 -2169 -1144 -2153
rect -920 -1177 -886 -1161
rect -920 -2169 -886 -2153
rect -662 -1177 -628 -1161
rect -662 -2169 -628 -2153
rect -404 -1177 -370 -1161
rect -404 -2169 -370 -2153
rect -146 -1177 -112 -1161
rect -146 -2169 -112 -2153
rect 112 -1177 146 -1161
rect 112 -2169 146 -2153
rect 370 -1177 404 -1161
rect 370 -2169 404 -2153
rect 628 -1177 662 -1161
rect 628 -2169 662 -2153
rect 886 -1177 920 -1161
rect 886 -2169 920 -2153
rect 1144 -1177 1178 -1161
rect 1144 -2169 1178 -2153
rect 1402 -1177 1436 -1161
rect 1402 -2169 1436 -2153
rect 1660 -1177 1694 -1161
rect 1660 -2169 1694 -2153
rect 1918 -1177 1952 -1161
rect 1918 -2169 1952 -2153
rect 2176 -1177 2210 -1161
rect 2176 -2169 2210 -2153
rect 2434 -1177 2468 -1161
rect 2434 -2169 2468 -2153
rect 2692 -1177 2726 -1161
rect 2692 -2169 2726 -2153
rect 2950 -1177 2984 -1161
rect 2950 -2169 2984 -2153
rect 3208 -1177 3242 -1161
rect 3208 -2169 3242 -2153
rect 3466 -1177 3500 -1161
rect 3466 -2169 3500 -2153
rect 3724 -1177 3758 -1161
rect 3724 -2169 3758 -2153
rect 3982 -1177 4016 -1161
rect 3982 -2169 4016 -2153
rect 4240 -1177 4274 -1161
rect 4240 -2169 4274 -2153
rect 4498 -1177 4532 -1161
rect 4498 -2169 4532 -2153
rect 4756 -1177 4790 -1161
rect 4756 -2169 4790 -2153
rect 5014 -1177 5048 -1161
rect 5014 -2169 5048 -2153
rect 5272 -1177 5306 -1161
rect 5272 -2169 5306 -2153
rect 5530 -1177 5564 -1161
rect 5530 -2169 5564 -2153
rect 5788 -1177 5822 -1161
rect 5788 -2169 5822 -2153
rect 6046 -1177 6080 -1161
rect 6046 -2169 6080 -2153
rect 6304 -1177 6338 -1161
rect 6304 -2169 6338 -2153
rect 6562 -1177 6596 -1161
rect 6562 -2169 6596 -2153
rect 6820 -1177 6854 -1161
rect 6820 -2169 6854 -2153
rect 7078 -1177 7112 -1161
rect 7078 -2169 7112 -2153
rect -7066 -2237 -7050 -2203
rect -6882 -2237 -6866 -2203
rect -6808 -2237 -6792 -2203
rect -6624 -2237 -6608 -2203
rect -6550 -2237 -6534 -2203
rect -6366 -2237 -6350 -2203
rect -6292 -2237 -6276 -2203
rect -6108 -2237 -6092 -2203
rect -6034 -2237 -6018 -2203
rect -5850 -2237 -5834 -2203
rect -5776 -2237 -5760 -2203
rect -5592 -2237 -5576 -2203
rect -5518 -2237 -5502 -2203
rect -5334 -2237 -5318 -2203
rect -5260 -2237 -5244 -2203
rect -5076 -2237 -5060 -2203
rect -5002 -2237 -4986 -2203
rect -4818 -2237 -4802 -2203
rect -4744 -2237 -4728 -2203
rect -4560 -2237 -4544 -2203
rect -4486 -2237 -4470 -2203
rect -4302 -2237 -4286 -2203
rect -4228 -2237 -4212 -2203
rect -4044 -2237 -4028 -2203
rect -3970 -2237 -3954 -2203
rect -3786 -2237 -3770 -2203
rect -3712 -2237 -3696 -2203
rect -3528 -2237 -3512 -2203
rect -3454 -2237 -3438 -2203
rect -3270 -2237 -3254 -2203
rect -3196 -2237 -3180 -2203
rect -3012 -2237 -2996 -2203
rect -2938 -2237 -2922 -2203
rect -2754 -2237 -2738 -2203
rect -2680 -2237 -2664 -2203
rect -2496 -2237 -2480 -2203
rect -2422 -2237 -2406 -2203
rect -2238 -2237 -2222 -2203
rect -2164 -2237 -2148 -2203
rect -1980 -2237 -1964 -2203
rect -1906 -2237 -1890 -2203
rect -1722 -2237 -1706 -2203
rect -1648 -2237 -1632 -2203
rect -1464 -2237 -1448 -2203
rect -1390 -2237 -1374 -2203
rect -1206 -2237 -1190 -2203
rect -1132 -2237 -1116 -2203
rect -948 -2237 -932 -2203
rect -874 -2237 -858 -2203
rect -690 -2237 -674 -2203
rect -616 -2237 -600 -2203
rect -432 -2237 -416 -2203
rect -358 -2237 -342 -2203
rect -174 -2237 -158 -2203
rect -100 -2237 -84 -2203
rect 84 -2237 100 -2203
rect 158 -2237 174 -2203
rect 342 -2237 358 -2203
rect 416 -2237 432 -2203
rect 600 -2237 616 -2203
rect 674 -2237 690 -2203
rect 858 -2237 874 -2203
rect 932 -2237 948 -2203
rect 1116 -2237 1132 -2203
rect 1190 -2237 1206 -2203
rect 1374 -2237 1390 -2203
rect 1448 -2237 1464 -2203
rect 1632 -2237 1648 -2203
rect 1706 -2237 1722 -2203
rect 1890 -2237 1906 -2203
rect 1964 -2237 1980 -2203
rect 2148 -2237 2164 -2203
rect 2222 -2237 2238 -2203
rect 2406 -2237 2422 -2203
rect 2480 -2237 2496 -2203
rect 2664 -2237 2680 -2203
rect 2738 -2237 2754 -2203
rect 2922 -2237 2938 -2203
rect 2996 -2237 3012 -2203
rect 3180 -2237 3196 -2203
rect 3254 -2237 3270 -2203
rect 3438 -2237 3454 -2203
rect 3512 -2237 3528 -2203
rect 3696 -2237 3712 -2203
rect 3770 -2237 3786 -2203
rect 3954 -2237 3970 -2203
rect 4028 -2237 4044 -2203
rect 4212 -2237 4228 -2203
rect 4286 -2237 4302 -2203
rect 4470 -2237 4486 -2203
rect 4544 -2237 4560 -2203
rect 4728 -2237 4744 -2203
rect 4802 -2237 4818 -2203
rect 4986 -2237 5002 -2203
rect 5060 -2237 5076 -2203
rect 5244 -2237 5260 -2203
rect 5318 -2237 5334 -2203
rect 5502 -2237 5518 -2203
rect 5576 -2237 5592 -2203
rect 5760 -2237 5776 -2203
rect 5834 -2237 5850 -2203
rect 6018 -2237 6034 -2203
rect 6092 -2237 6108 -2203
rect 6276 -2237 6292 -2203
rect 6350 -2237 6366 -2203
rect 6534 -2237 6550 -2203
rect 6608 -2237 6624 -2203
rect 6792 -2237 6808 -2203
rect 6866 -2237 6882 -2203
rect 7050 -2237 7066 -2203
rect -7246 -2341 -7212 -2279
rect 7212 -2341 7246 -2279
rect -7246 -2375 -7150 -2341
rect 7150 -2375 7246 -2341
<< viali >>
rect -7050 2203 -6882 2237
rect -6792 2203 -6624 2237
rect -6534 2203 -6366 2237
rect -6276 2203 -6108 2237
rect -6018 2203 -5850 2237
rect -5760 2203 -5592 2237
rect -5502 2203 -5334 2237
rect -5244 2203 -5076 2237
rect -4986 2203 -4818 2237
rect -4728 2203 -4560 2237
rect -4470 2203 -4302 2237
rect -4212 2203 -4044 2237
rect -3954 2203 -3786 2237
rect -3696 2203 -3528 2237
rect -3438 2203 -3270 2237
rect -3180 2203 -3012 2237
rect -2922 2203 -2754 2237
rect -2664 2203 -2496 2237
rect -2406 2203 -2238 2237
rect -2148 2203 -1980 2237
rect -1890 2203 -1722 2237
rect -1632 2203 -1464 2237
rect -1374 2203 -1206 2237
rect -1116 2203 -948 2237
rect -858 2203 -690 2237
rect -600 2203 -432 2237
rect -342 2203 -174 2237
rect -84 2203 84 2237
rect 174 2203 342 2237
rect 432 2203 600 2237
rect 690 2203 858 2237
rect 948 2203 1116 2237
rect 1206 2203 1374 2237
rect 1464 2203 1632 2237
rect 1722 2203 1890 2237
rect 1980 2203 2148 2237
rect 2238 2203 2406 2237
rect 2496 2203 2664 2237
rect 2754 2203 2922 2237
rect 3012 2203 3180 2237
rect 3270 2203 3438 2237
rect 3528 2203 3696 2237
rect 3786 2203 3954 2237
rect 4044 2203 4212 2237
rect 4302 2203 4470 2237
rect 4560 2203 4728 2237
rect 4818 2203 4986 2237
rect 5076 2203 5244 2237
rect 5334 2203 5502 2237
rect 5592 2203 5760 2237
rect 5850 2203 6018 2237
rect 6108 2203 6276 2237
rect 6366 2203 6534 2237
rect 6624 2203 6792 2237
rect 6882 2203 7050 2237
rect -7112 1177 -7078 2153
rect -6854 1177 -6820 2153
rect -6596 1177 -6562 2153
rect -6338 1177 -6304 2153
rect -6080 1177 -6046 2153
rect -5822 1177 -5788 2153
rect -5564 1177 -5530 2153
rect -5306 1177 -5272 2153
rect -5048 1177 -5014 2153
rect -4790 1177 -4756 2153
rect -4532 1177 -4498 2153
rect -4274 1177 -4240 2153
rect -4016 1177 -3982 2153
rect -3758 1177 -3724 2153
rect -3500 1177 -3466 2153
rect -3242 1177 -3208 2153
rect -2984 1177 -2950 2153
rect -2726 1177 -2692 2153
rect -2468 1177 -2434 2153
rect -2210 1177 -2176 2153
rect -1952 1177 -1918 2153
rect -1694 1177 -1660 2153
rect -1436 1177 -1402 2153
rect -1178 1177 -1144 2153
rect -920 1177 -886 2153
rect -662 1177 -628 2153
rect -404 1177 -370 2153
rect -146 1177 -112 2153
rect 112 1177 146 2153
rect 370 1177 404 2153
rect 628 1177 662 2153
rect 886 1177 920 2153
rect 1144 1177 1178 2153
rect 1402 1177 1436 2153
rect 1660 1177 1694 2153
rect 1918 1177 1952 2153
rect 2176 1177 2210 2153
rect 2434 1177 2468 2153
rect 2692 1177 2726 2153
rect 2950 1177 2984 2153
rect 3208 1177 3242 2153
rect 3466 1177 3500 2153
rect 3724 1177 3758 2153
rect 3982 1177 4016 2153
rect 4240 1177 4274 2153
rect 4498 1177 4532 2153
rect 4756 1177 4790 2153
rect 5014 1177 5048 2153
rect 5272 1177 5306 2153
rect 5530 1177 5564 2153
rect 5788 1177 5822 2153
rect 6046 1177 6080 2153
rect 6304 1177 6338 2153
rect 6562 1177 6596 2153
rect 6820 1177 6854 2153
rect 7078 1177 7112 2153
rect -7050 1093 -6882 1127
rect -6792 1093 -6624 1127
rect -6534 1093 -6366 1127
rect -6276 1093 -6108 1127
rect -6018 1093 -5850 1127
rect -5760 1093 -5592 1127
rect -5502 1093 -5334 1127
rect -5244 1093 -5076 1127
rect -4986 1093 -4818 1127
rect -4728 1093 -4560 1127
rect -4470 1093 -4302 1127
rect -4212 1093 -4044 1127
rect -3954 1093 -3786 1127
rect -3696 1093 -3528 1127
rect -3438 1093 -3270 1127
rect -3180 1093 -3012 1127
rect -2922 1093 -2754 1127
rect -2664 1093 -2496 1127
rect -2406 1093 -2238 1127
rect -2148 1093 -1980 1127
rect -1890 1093 -1722 1127
rect -1632 1093 -1464 1127
rect -1374 1093 -1206 1127
rect -1116 1093 -948 1127
rect -858 1093 -690 1127
rect -600 1093 -432 1127
rect -342 1093 -174 1127
rect -84 1093 84 1127
rect 174 1093 342 1127
rect 432 1093 600 1127
rect 690 1093 858 1127
rect 948 1093 1116 1127
rect 1206 1093 1374 1127
rect 1464 1093 1632 1127
rect 1722 1093 1890 1127
rect 1980 1093 2148 1127
rect 2238 1093 2406 1127
rect 2496 1093 2664 1127
rect 2754 1093 2922 1127
rect 3012 1093 3180 1127
rect 3270 1093 3438 1127
rect 3528 1093 3696 1127
rect 3786 1093 3954 1127
rect 4044 1093 4212 1127
rect 4302 1093 4470 1127
rect 4560 1093 4728 1127
rect 4818 1093 4986 1127
rect 5076 1093 5244 1127
rect 5334 1093 5502 1127
rect 5592 1093 5760 1127
rect 5850 1093 6018 1127
rect 6108 1093 6276 1127
rect 6366 1093 6534 1127
rect 6624 1093 6792 1127
rect 6882 1093 7050 1127
rect -7112 67 -7078 1043
rect -6854 67 -6820 1043
rect -6596 67 -6562 1043
rect -6338 67 -6304 1043
rect -6080 67 -6046 1043
rect -5822 67 -5788 1043
rect -5564 67 -5530 1043
rect -5306 67 -5272 1043
rect -5048 67 -5014 1043
rect -4790 67 -4756 1043
rect -4532 67 -4498 1043
rect -4274 67 -4240 1043
rect -4016 67 -3982 1043
rect -3758 67 -3724 1043
rect -3500 67 -3466 1043
rect -3242 67 -3208 1043
rect -2984 67 -2950 1043
rect -2726 67 -2692 1043
rect -2468 67 -2434 1043
rect -2210 67 -2176 1043
rect -1952 67 -1918 1043
rect -1694 67 -1660 1043
rect -1436 67 -1402 1043
rect -1178 67 -1144 1043
rect -920 67 -886 1043
rect -662 67 -628 1043
rect -404 67 -370 1043
rect -146 67 -112 1043
rect 112 67 146 1043
rect 370 67 404 1043
rect 628 67 662 1043
rect 886 67 920 1043
rect 1144 67 1178 1043
rect 1402 67 1436 1043
rect 1660 67 1694 1043
rect 1918 67 1952 1043
rect 2176 67 2210 1043
rect 2434 67 2468 1043
rect 2692 67 2726 1043
rect 2950 67 2984 1043
rect 3208 67 3242 1043
rect 3466 67 3500 1043
rect 3724 67 3758 1043
rect 3982 67 4016 1043
rect 4240 67 4274 1043
rect 4498 67 4532 1043
rect 4756 67 4790 1043
rect 5014 67 5048 1043
rect 5272 67 5306 1043
rect 5530 67 5564 1043
rect 5788 67 5822 1043
rect 6046 67 6080 1043
rect 6304 67 6338 1043
rect 6562 67 6596 1043
rect 6820 67 6854 1043
rect 7078 67 7112 1043
rect -7050 -17 -6882 17
rect -6792 -17 -6624 17
rect -6534 -17 -6366 17
rect -6276 -17 -6108 17
rect -6018 -17 -5850 17
rect -5760 -17 -5592 17
rect -5502 -17 -5334 17
rect -5244 -17 -5076 17
rect -4986 -17 -4818 17
rect -4728 -17 -4560 17
rect -4470 -17 -4302 17
rect -4212 -17 -4044 17
rect -3954 -17 -3786 17
rect -3696 -17 -3528 17
rect -3438 -17 -3270 17
rect -3180 -17 -3012 17
rect -2922 -17 -2754 17
rect -2664 -17 -2496 17
rect -2406 -17 -2238 17
rect -2148 -17 -1980 17
rect -1890 -17 -1722 17
rect -1632 -17 -1464 17
rect -1374 -17 -1206 17
rect -1116 -17 -948 17
rect -858 -17 -690 17
rect -600 -17 -432 17
rect -342 -17 -174 17
rect -84 -17 84 17
rect 174 -17 342 17
rect 432 -17 600 17
rect 690 -17 858 17
rect 948 -17 1116 17
rect 1206 -17 1374 17
rect 1464 -17 1632 17
rect 1722 -17 1890 17
rect 1980 -17 2148 17
rect 2238 -17 2406 17
rect 2496 -17 2664 17
rect 2754 -17 2922 17
rect 3012 -17 3180 17
rect 3270 -17 3438 17
rect 3528 -17 3696 17
rect 3786 -17 3954 17
rect 4044 -17 4212 17
rect 4302 -17 4470 17
rect 4560 -17 4728 17
rect 4818 -17 4986 17
rect 5076 -17 5244 17
rect 5334 -17 5502 17
rect 5592 -17 5760 17
rect 5850 -17 6018 17
rect 6108 -17 6276 17
rect 6366 -17 6534 17
rect 6624 -17 6792 17
rect 6882 -17 7050 17
rect -7112 -1043 -7078 -67
rect -6854 -1043 -6820 -67
rect -6596 -1043 -6562 -67
rect -6338 -1043 -6304 -67
rect -6080 -1043 -6046 -67
rect -5822 -1043 -5788 -67
rect -5564 -1043 -5530 -67
rect -5306 -1043 -5272 -67
rect -5048 -1043 -5014 -67
rect -4790 -1043 -4756 -67
rect -4532 -1043 -4498 -67
rect -4274 -1043 -4240 -67
rect -4016 -1043 -3982 -67
rect -3758 -1043 -3724 -67
rect -3500 -1043 -3466 -67
rect -3242 -1043 -3208 -67
rect -2984 -1043 -2950 -67
rect -2726 -1043 -2692 -67
rect -2468 -1043 -2434 -67
rect -2210 -1043 -2176 -67
rect -1952 -1043 -1918 -67
rect -1694 -1043 -1660 -67
rect -1436 -1043 -1402 -67
rect -1178 -1043 -1144 -67
rect -920 -1043 -886 -67
rect -662 -1043 -628 -67
rect -404 -1043 -370 -67
rect -146 -1043 -112 -67
rect 112 -1043 146 -67
rect 370 -1043 404 -67
rect 628 -1043 662 -67
rect 886 -1043 920 -67
rect 1144 -1043 1178 -67
rect 1402 -1043 1436 -67
rect 1660 -1043 1694 -67
rect 1918 -1043 1952 -67
rect 2176 -1043 2210 -67
rect 2434 -1043 2468 -67
rect 2692 -1043 2726 -67
rect 2950 -1043 2984 -67
rect 3208 -1043 3242 -67
rect 3466 -1043 3500 -67
rect 3724 -1043 3758 -67
rect 3982 -1043 4016 -67
rect 4240 -1043 4274 -67
rect 4498 -1043 4532 -67
rect 4756 -1043 4790 -67
rect 5014 -1043 5048 -67
rect 5272 -1043 5306 -67
rect 5530 -1043 5564 -67
rect 5788 -1043 5822 -67
rect 6046 -1043 6080 -67
rect 6304 -1043 6338 -67
rect 6562 -1043 6596 -67
rect 6820 -1043 6854 -67
rect 7078 -1043 7112 -67
rect -7050 -1127 -6882 -1093
rect -6792 -1127 -6624 -1093
rect -6534 -1127 -6366 -1093
rect -6276 -1127 -6108 -1093
rect -6018 -1127 -5850 -1093
rect -5760 -1127 -5592 -1093
rect -5502 -1127 -5334 -1093
rect -5244 -1127 -5076 -1093
rect -4986 -1127 -4818 -1093
rect -4728 -1127 -4560 -1093
rect -4470 -1127 -4302 -1093
rect -4212 -1127 -4044 -1093
rect -3954 -1127 -3786 -1093
rect -3696 -1127 -3528 -1093
rect -3438 -1127 -3270 -1093
rect -3180 -1127 -3012 -1093
rect -2922 -1127 -2754 -1093
rect -2664 -1127 -2496 -1093
rect -2406 -1127 -2238 -1093
rect -2148 -1127 -1980 -1093
rect -1890 -1127 -1722 -1093
rect -1632 -1127 -1464 -1093
rect -1374 -1127 -1206 -1093
rect -1116 -1127 -948 -1093
rect -858 -1127 -690 -1093
rect -600 -1127 -432 -1093
rect -342 -1127 -174 -1093
rect -84 -1127 84 -1093
rect 174 -1127 342 -1093
rect 432 -1127 600 -1093
rect 690 -1127 858 -1093
rect 948 -1127 1116 -1093
rect 1206 -1127 1374 -1093
rect 1464 -1127 1632 -1093
rect 1722 -1127 1890 -1093
rect 1980 -1127 2148 -1093
rect 2238 -1127 2406 -1093
rect 2496 -1127 2664 -1093
rect 2754 -1127 2922 -1093
rect 3012 -1127 3180 -1093
rect 3270 -1127 3438 -1093
rect 3528 -1127 3696 -1093
rect 3786 -1127 3954 -1093
rect 4044 -1127 4212 -1093
rect 4302 -1127 4470 -1093
rect 4560 -1127 4728 -1093
rect 4818 -1127 4986 -1093
rect 5076 -1127 5244 -1093
rect 5334 -1127 5502 -1093
rect 5592 -1127 5760 -1093
rect 5850 -1127 6018 -1093
rect 6108 -1127 6276 -1093
rect 6366 -1127 6534 -1093
rect 6624 -1127 6792 -1093
rect 6882 -1127 7050 -1093
rect -7112 -2153 -7078 -1177
rect -6854 -2153 -6820 -1177
rect -6596 -2153 -6562 -1177
rect -6338 -2153 -6304 -1177
rect -6080 -2153 -6046 -1177
rect -5822 -2153 -5788 -1177
rect -5564 -2153 -5530 -1177
rect -5306 -2153 -5272 -1177
rect -5048 -2153 -5014 -1177
rect -4790 -2153 -4756 -1177
rect -4532 -2153 -4498 -1177
rect -4274 -2153 -4240 -1177
rect -4016 -2153 -3982 -1177
rect -3758 -2153 -3724 -1177
rect -3500 -2153 -3466 -1177
rect -3242 -2153 -3208 -1177
rect -2984 -2153 -2950 -1177
rect -2726 -2153 -2692 -1177
rect -2468 -2153 -2434 -1177
rect -2210 -2153 -2176 -1177
rect -1952 -2153 -1918 -1177
rect -1694 -2153 -1660 -1177
rect -1436 -2153 -1402 -1177
rect -1178 -2153 -1144 -1177
rect -920 -2153 -886 -1177
rect -662 -2153 -628 -1177
rect -404 -2153 -370 -1177
rect -146 -2153 -112 -1177
rect 112 -2153 146 -1177
rect 370 -2153 404 -1177
rect 628 -2153 662 -1177
rect 886 -2153 920 -1177
rect 1144 -2153 1178 -1177
rect 1402 -2153 1436 -1177
rect 1660 -2153 1694 -1177
rect 1918 -2153 1952 -1177
rect 2176 -2153 2210 -1177
rect 2434 -2153 2468 -1177
rect 2692 -2153 2726 -1177
rect 2950 -2153 2984 -1177
rect 3208 -2153 3242 -1177
rect 3466 -2153 3500 -1177
rect 3724 -2153 3758 -1177
rect 3982 -2153 4016 -1177
rect 4240 -2153 4274 -1177
rect 4498 -2153 4532 -1177
rect 4756 -2153 4790 -1177
rect 5014 -2153 5048 -1177
rect 5272 -2153 5306 -1177
rect 5530 -2153 5564 -1177
rect 5788 -2153 5822 -1177
rect 6046 -2153 6080 -1177
rect 6304 -2153 6338 -1177
rect 6562 -2153 6596 -1177
rect 6820 -2153 6854 -1177
rect 7078 -2153 7112 -1177
rect -7050 -2237 -6882 -2203
rect -6792 -2237 -6624 -2203
rect -6534 -2237 -6366 -2203
rect -6276 -2237 -6108 -2203
rect -6018 -2237 -5850 -2203
rect -5760 -2237 -5592 -2203
rect -5502 -2237 -5334 -2203
rect -5244 -2237 -5076 -2203
rect -4986 -2237 -4818 -2203
rect -4728 -2237 -4560 -2203
rect -4470 -2237 -4302 -2203
rect -4212 -2237 -4044 -2203
rect -3954 -2237 -3786 -2203
rect -3696 -2237 -3528 -2203
rect -3438 -2237 -3270 -2203
rect -3180 -2237 -3012 -2203
rect -2922 -2237 -2754 -2203
rect -2664 -2237 -2496 -2203
rect -2406 -2237 -2238 -2203
rect -2148 -2237 -1980 -2203
rect -1890 -2237 -1722 -2203
rect -1632 -2237 -1464 -2203
rect -1374 -2237 -1206 -2203
rect -1116 -2237 -948 -2203
rect -858 -2237 -690 -2203
rect -600 -2237 -432 -2203
rect -342 -2237 -174 -2203
rect -84 -2237 84 -2203
rect 174 -2237 342 -2203
rect 432 -2237 600 -2203
rect 690 -2237 858 -2203
rect 948 -2237 1116 -2203
rect 1206 -2237 1374 -2203
rect 1464 -2237 1632 -2203
rect 1722 -2237 1890 -2203
rect 1980 -2237 2148 -2203
rect 2238 -2237 2406 -2203
rect 2496 -2237 2664 -2203
rect 2754 -2237 2922 -2203
rect 3012 -2237 3180 -2203
rect 3270 -2237 3438 -2203
rect 3528 -2237 3696 -2203
rect 3786 -2237 3954 -2203
rect 4044 -2237 4212 -2203
rect 4302 -2237 4470 -2203
rect 4560 -2237 4728 -2203
rect 4818 -2237 4986 -2203
rect 5076 -2237 5244 -2203
rect 5334 -2237 5502 -2203
rect 5592 -2237 5760 -2203
rect 5850 -2237 6018 -2203
rect 6108 -2237 6276 -2203
rect 6366 -2237 6534 -2203
rect 6624 -2237 6792 -2203
rect 6882 -2237 7050 -2203
<< metal1 >>
rect -7062 2237 -6870 2243
rect -7062 2203 -7050 2237
rect -6882 2203 -6870 2237
rect -7062 2197 -6870 2203
rect -6804 2237 -6612 2243
rect -6804 2203 -6792 2237
rect -6624 2203 -6612 2237
rect -6804 2197 -6612 2203
rect -6546 2237 -6354 2243
rect -6546 2203 -6534 2237
rect -6366 2203 -6354 2237
rect -6546 2197 -6354 2203
rect -6288 2237 -6096 2243
rect -6288 2203 -6276 2237
rect -6108 2203 -6096 2237
rect -6288 2197 -6096 2203
rect -6030 2237 -5838 2243
rect -6030 2203 -6018 2237
rect -5850 2203 -5838 2237
rect -6030 2197 -5838 2203
rect -5772 2237 -5580 2243
rect -5772 2203 -5760 2237
rect -5592 2203 -5580 2237
rect -5772 2197 -5580 2203
rect -5514 2237 -5322 2243
rect -5514 2203 -5502 2237
rect -5334 2203 -5322 2237
rect -5514 2197 -5322 2203
rect -5256 2237 -5064 2243
rect -5256 2203 -5244 2237
rect -5076 2203 -5064 2237
rect -5256 2197 -5064 2203
rect -4998 2237 -4806 2243
rect -4998 2203 -4986 2237
rect -4818 2203 -4806 2237
rect -4998 2197 -4806 2203
rect -4740 2237 -4548 2243
rect -4740 2203 -4728 2237
rect -4560 2203 -4548 2237
rect -4740 2197 -4548 2203
rect -4482 2237 -4290 2243
rect -4482 2203 -4470 2237
rect -4302 2203 -4290 2237
rect -4482 2197 -4290 2203
rect -4224 2237 -4032 2243
rect -4224 2203 -4212 2237
rect -4044 2203 -4032 2237
rect -4224 2197 -4032 2203
rect -3966 2237 -3774 2243
rect -3966 2203 -3954 2237
rect -3786 2203 -3774 2237
rect -3966 2197 -3774 2203
rect -3708 2237 -3516 2243
rect -3708 2203 -3696 2237
rect -3528 2203 -3516 2237
rect -3708 2197 -3516 2203
rect -3450 2237 -3258 2243
rect -3450 2203 -3438 2237
rect -3270 2203 -3258 2237
rect -3450 2197 -3258 2203
rect -3192 2237 -3000 2243
rect -3192 2203 -3180 2237
rect -3012 2203 -3000 2237
rect -3192 2197 -3000 2203
rect -2934 2237 -2742 2243
rect -2934 2203 -2922 2237
rect -2754 2203 -2742 2237
rect -2934 2197 -2742 2203
rect -2676 2237 -2484 2243
rect -2676 2203 -2664 2237
rect -2496 2203 -2484 2237
rect -2676 2197 -2484 2203
rect -2418 2237 -2226 2243
rect -2418 2203 -2406 2237
rect -2238 2203 -2226 2237
rect -2418 2197 -2226 2203
rect -2160 2237 -1968 2243
rect -2160 2203 -2148 2237
rect -1980 2203 -1968 2237
rect -2160 2197 -1968 2203
rect -1902 2237 -1710 2243
rect -1902 2203 -1890 2237
rect -1722 2203 -1710 2237
rect -1902 2197 -1710 2203
rect -1644 2237 -1452 2243
rect -1644 2203 -1632 2237
rect -1464 2203 -1452 2237
rect -1644 2197 -1452 2203
rect -1386 2237 -1194 2243
rect -1386 2203 -1374 2237
rect -1206 2203 -1194 2237
rect -1386 2197 -1194 2203
rect -1128 2237 -936 2243
rect -1128 2203 -1116 2237
rect -948 2203 -936 2237
rect -1128 2197 -936 2203
rect -870 2237 -678 2243
rect -870 2203 -858 2237
rect -690 2203 -678 2237
rect -870 2197 -678 2203
rect -612 2237 -420 2243
rect -612 2203 -600 2237
rect -432 2203 -420 2237
rect -612 2197 -420 2203
rect -354 2237 -162 2243
rect -354 2203 -342 2237
rect -174 2203 -162 2237
rect -354 2197 -162 2203
rect -96 2237 96 2243
rect -96 2203 -84 2237
rect 84 2203 96 2237
rect -96 2197 96 2203
rect 162 2237 354 2243
rect 162 2203 174 2237
rect 342 2203 354 2237
rect 162 2197 354 2203
rect 420 2237 612 2243
rect 420 2203 432 2237
rect 600 2203 612 2237
rect 420 2197 612 2203
rect 678 2237 870 2243
rect 678 2203 690 2237
rect 858 2203 870 2237
rect 678 2197 870 2203
rect 936 2237 1128 2243
rect 936 2203 948 2237
rect 1116 2203 1128 2237
rect 936 2197 1128 2203
rect 1194 2237 1386 2243
rect 1194 2203 1206 2237
rect 1374 2203 1386 2237
rect 1194 2197 1386 2203
rect 1452 2237 1644 2243
rect 1452 2203 1464 2237
rect 1632 2203 1644 2237
rect 1452 2197 1644 2203
rect 1710 2237 1902 2243
rect 1710 2203 1722 2237
rect 1890 2203 1902 2237
rect 1710 2197 1902 2203
rect 1968 2237 2160 2243
rect 1968 2203 1980 2237
rect 2148 2203 2160 2237
rect 1968 2197 2160 2203
rect 2226 2237 2418 2243
rect 2226 2203 2238 2237
rect 2406 2203 2418 2237
rect 2226 2197 2418 2203
rect 2484 2237 2676 2243
rect 2484 2203 2496 2237
rect 2664 2203 2676 2237
rect 2484 2197 2676 2203
rect 2742 2237 2934 2243
rect 2742 2203 2754 2237
rect 2922 2203 2934 2237
rect 2742 2197 2934 2203
rect 3000 2237 3192 2243
rect 3000 2203 3012 2237
rect 3180 2203 3192 2237
rect 3000 2197 3192 2203
rect 3258 2237 3450 2243
rect 3258 2203 3270 2237
rect 3438 2203 3450 2237
rect 3258 2197 3450 2203
rect 3516 2237 3708 2243
rect 3516 2203 3528 2237
rect 3696 2203 3708 2237
rect 3516 2197 3708 2203
rect 3774 2237 3966 2243
rect 3774 2203 3786 2237
rect 3954 2203 3966 2237
rect 3774 2197 3966 2203
rect 4032 2237 4224 2243
rect 4032 2203 4044 2237
rect 4212 2203 4224 2237
rect 4032 2197 4224 2203
rect 4290 2237 4482 2243
rect 4290 2203 4302 2237
rect 4470 2203 4482 2237
rect 4290 2197 4482 2203
rect 4548 2237 4740 2243
rect 4548 2203 4560 2237
rect 4728 2203 4740 2237
rect 4548 2197 4740 2203
rect 4806 2237 4998 2243
rect 4806 2203 4818 2237
rect 4986 2203 4998 2237
rect 4806 2197 4998 2203
rect 5064 2237 5256 2243
rect 5064 2203 5076 2237
rect 5244 2203 5256 2237
rect 5064 2197 5256 2203
rect 5322 2237 5514 2243
rect 5322 2203 5334 2237
rect 5502 2203 5514 2237
rect 5322 2197 5514 2203
rect 5580 2237 5772 2243
rect 5580 2203 5592 2237
rect 5760 2203 5772 2237
rect 5580 2197 5772 2203
rect 5838 2237 6030 2243
rect 5838 2203 5850 2237
rect 6018 2203 6030 2237
rect 5838 2197 6030 2203
rect 6096 2237 6288 2243
rect 6096 2203 6108 2237
rect 6276 2203 6288 2237
rect 6096 2197 6288 2203
rect 6354 2237 6546 2243
rect 6354 2203 6366 2237
rect 6534 2203 6546 2237
rect 6354 2197 6546 2203
rect 6612 2237 6804 2243
rect 6612 2203 6624 2237
rect 6792 2203 6804 2237
rect 6612 2197 6804 2203
rect 6870 2237 7062 2243
rect 6870 2203 6882 2237
rect 7050 2203 7062 2237
rect 6870 2197 7062 2203
rect -7118 2153 -7072 2165
rect -7118 1177 -7112 2153
rect -7078 1177 -7072 2153
rect -7118 1165 -7072 1177
rect -6860 2153 -6814 2165
rect -6860 1177 -6854 2153
rect -6820 1177 -6814 2153
rect -6860 1165 -6814 1177
rect -6602 2153 -6556 2165
rect -6602 1177 -6596 2153
rect -6562 1177 -6556 2153
rect -6602 1165 -6556 1177
rect -6344 2153 -6298 2165
rect -6344 1177 -6338 2153
rect -6304 1177 -6298 2153
rect -6344 1165 -6298 1177
rect -6086 2153 -6040 2165
rect -6086 1177 -6080 2153
rect -6046 1177 -6040 2153
rect -6086 1165 -6040 1177
rect -5828 2153 -5782 2165
rect -5828 1177 -5822 2153
rect -5788 1177 -5782 2153
rect -5828 1165 -5782 1177
rect -5570 2153 -5524 2165
rect -5570 1177 -5564 2153
rect -5530 1177 -5524 2153
rect -5570 1165 -5524 1177
rect -5312 2153 -5266 2165
rect -5312 1177 -5306 2153
rect -5272 1177 -5266 2153
rect -5312 1165 -5266 1177
rect -5054 2153 -5008 2165
rect -5054 1177 -5048 2153
rect -5014 1177 -5008 2153
rect -5054 1165 -5008 1177
rect -4796 2153 -4750 2165
rect -4796 1177 -4790 2153
rect -4756 1177 -4750 2153
rect -4796 1165 -4750 1177
rect -4538 2153 -4492 2165
rect -4538 1177 -4532 2153
rect -4498 1177 -4492 2153
rect -4538 1165 -4492 1177
rect -4280 2153 -4234 2165
rect -4280 1177 -4274 2153
rect -4240 1177 -4234 2153
rect -4280 1165 -4234 1177
rect -4022 2153 -3976 2165
rect -4022 1177 -4016 2153
rect -3982 1177 -3976 2153
rect -4022 1165 -3976 1177
rect -3764 2153 -3718 2165
rect -3764 1177 -3758 2153
rect -3724 1177 -3718 2153
rect -3764 1165 -3718 1177
rect -3506 2153 -3460 2165
rect -3506 1177 -3500 2153
rect -3466 1177 -3460 2153
rect -3506 1165 -3460 1177
rect -3248 2153 -3202 2165
rect -3248 1177 -3242 2153
rect -3208 1177 -3202 2153
rect -3248 1165 -3202 1177
rect -2990 2153 -2944 2165
rect -2990 1177 -2984 2153
rect -2950 1177 -2944 2153
rect -2990 1165 -2944 1177
rect -2732 2153 -2686 2165
rect -2732 1177 -2726 2153
rect -2692 1177 -2686 2153
rect -2732 1165 -2686 1177
rect -2474 2153 -2428 2165
rect -2474 1177 -2468 2153
rect -2434 1177 -2428 2153
rect -2474 1165 -2428 1177
rect -2216 2153 -2170 2165
rect -2216 1177 -2210 2153
rect -2176 1177 -2170 2153
rect -2216 1165 -2170 1177
rect -1958 2153 -1912 2165
rect -1958 1177 -1952 2153
rect -1918 1177 -1912 2153
rect -1958 1165 -1912 1177
rect -1700 2153 -1654 2165
rect -1700 1177 -1694 2153
rect -1660 1177 -1654 2153
rect -1700 1165 -1654 1177
rect -1442 2153 -1396 2165
rect -1442 1177 -1436 2153
rect -1402 1177 -1396 2153
rect -1442 1165 -1396 1177
rect -1184 2153 -1138 2165
rect -1184 1177 -1178 2153
rect -1144 1177 -1138 2153
rect -1184 1165 -1138 1177
rect -926 2153 -880 2165
rect -926 1177 -920 2153
rect -886 1177 -880 2153
rect -926 1165 -880 1177
rect -668 2153 -622 2165
rect -668 1177 -662 2153
rect -628 1177 -622 2153
rect -668 1165 -622 1177
rect -410 2153 -364 2165
rect -410 1177 -404 2153
rect -370 1177 -364 2153
rect -410 1165 -364 1177
rect -152 2153 -106 2165
rect -152 1177 -146 2153
rect -112 1177 -106 2153
rect -152 1165 -106 1177
rect 106 2153 152 2165
rect 106 1177 112 2153
rect 146 1177 152 2153
rect 106 1165 152 1177
rect 364 2153 410 2165
rect 364 1177 370 2153
rect 404 1177 410 2153
rect 364 1165 410 1177
rect 622 2153 668 2165
rect 622 1177 628 2153
rect 662 1177 668 2153
rect 622 1165 668 1177
rect 880 2153 926 2165
rect 880 1177 886 2153
rect 920 1177 926 2153
rect 880 1165 926 1177
rect 1138 2153 1184 2165
rect 1138 1177 1144 2153
rect 1178 1177 1184 2153
rect 1138 1165 1184 1177
rect 1396 2153 1442 2165
rect 1396 1177 1402 2153
rect 1436 1177 1442 2153
rect 1396 1165 1442 1177
rect 1654 2153 1700 2165
rect 1654 1177 1660 2153
rect 1694 1177 1700 2153
rect 1654 1165 1700 1177
rect 1912 2153 1958 2165
rect 1912 1177 1918 2153
rect 1952 1177 1958 2153
rect 1912 1165 1958 1177
rect 2170 2153 2216 2165
rect 2170 1177 2176 2153
rect 2210 1177 2216 2153
rect 2170 1165 2216 1177
rect 2428 2153 2474 2165
rect 2428 1177 2434 2153
rect 2468 1177 2474 2153
rect 2428 1165 2474 1177
rect 2686 2153 2732 2165
rect 2686 1177 2692 2153
rect 2726 1177 2732 2153
rect 2686 1165 2732 1177
rect 2944 2153 2990 2165
rect 2944 1177 2950 2153
rect 2984 1177 2990 2153
rect 2944 1165 2990 1177
rect 3202 2153 3248 2165
rect 3202 1177 3208 2153
rect 3242 1177 3248 2153
rect 3202 1165 3248 1177
rect 3460 2153 3506 2165
rect 3460 1177 3466 2153
rect 3500 1177 3506 2153
rect 3460 1165 3506 1177
rect 3718 2153 3764 2165
rect 3718 1177 3724 2153
rect 3758 1177 3764 2153
rect 3718 1165 3764 1177
rect 3976 2153 4022 2165
rect 3976 1177 3982 2153
rect 4016 1177 4022 2153
rect 3976 1165 4022 1177
rect 4234 2153 4280 2165
rect 4234 1177 4240 2153
rect 4274 1177 4280 2153
rect 4234 1165 4280 1177
rect 4492 2153 4538 2165
rect 4492 1177 4498 2153
rect 4532 1177 4538 2153
rect 4492 1165 4538 1177
rect 4750 2153 4796 2165
rect 4750 1177 4756 2153
rect 4790 1177 4796 2153
rect 4750 1165 4796 1177
rect 5008 2153 5054 2165
rect 5008 1177 5014 2153
rect 5048 1177 5054 2153
rect 5008 1165 5054 1177
rect 5266 2153 5312 2165
rect 5266 1177 5272 2153
rect 5306 1177 5312 2153
rect 5266 1165 5312 1177
rect 5524 2153 5570 2165
rect 5524 1177 5530 2153
rect 5564 1177 5570 2153
rect 5524 1165 5570 1177
rect 5782 2153 5828 2165
rect 5782 1177 5788 2153
rect 5822 1177 5828 2153
rect 5782 1165 5828 1177
rect 6040 2153 6086 2165
rect 6040 1177 6046 2153
rect 6080 1177 6086 2153
rect 6040 1165 6086 1177
rect 6298 2153 6344 2165
rect 6298 1177 6304 2153
rect 6338 1177 6344 2153
rect 6298 1165 6344 1177
rect 6556 2153 6602 2165
rect 6556 1177 6562 2153
rect 6596 1177 6602 2153
rect 6556 1165 6602 1177
rect 6814 2153 6860 2165
rect 6814 1177 6820 2153
rect 6854 1177 6860 2153
rect 6814 1165 6860 1177
rect 7072 2153 7118 2165
rect 7072 1177 7078 2153
rect 7112 1177 7118 2153
rect 7072 1165 7118 1177
rect -7062 1127 -6870 1133
rect -7062 1093 -7050 1127
rect -6882 1093 -6870 1127
rect -7062 1087 -6870 1093
rect -6804 1127 -6612 1133
rect -6804 1093 -6792 1127
rect -6624 1093 -6612 1127
rect -6804 1087 -6612 1093
rect -6546 1127 -6354 1133
rect -6546 1093 -6534 1127
rect -6366 1093 -6354 1127
rect -6546 1087 -6354 1093
rect -6288 1127 -6096 1133
rect -6288 1093 -6276 1127
rect -6108 1093 -6096 1127
rect -6288 1087 -6096 1093
rect -6030 1127 -5838 1133
rect -6030 1093 -6018 1127
rect -5850 1093 -5838 1127
rect -6030 1087 -5838 1093
rect -5772 1127 -5580 1133
rect -5772 1093 -5760 1127
rect -5592 1093 -5580 1127
rect -5772 1087 -5580 1093
rect -5514 1127 -5322 1133
rect -5514 1093 -5502 1127
rect -5334 1093 -5322 1127
rect -5514 1087 -5322 1093
rect -5256 1127 -5064 1133
rect -5256 1093 -5244 1127
rect -5076 1093 -5064 1127
rect -5256 1087 -5064 1093
rect -4998 1127 -4806 1133
rect -4998 1093 -4986 1127
rect -4818 1093 -4806 1127
rect -4998 1087 -4806 1093
rect -4740 1127 -4548 1133
rect -4740 1093 -4728 1127
rect -4560 1093 -4548 1127
rect -4740 1087 -4548 1093
rect -4482 1127 -4290 1133
rect -4482 1093 -4470 1127
rect -4302 1093 -4290 1127
rect -4482 1087 -4290 1093
rect -4224 1127 -4032 1133
rect -4224 1093 -4212 1127
rect -4044 1093 -4032 1127
rect -4224 1087 -4032 1093
rect -3966 1127 -3774 1133
rect -3966 1093 -3954 1127
rect -3786 1093 -3774 1127
rect -3966 1087 -3774 1093
rect -3708 1127 -3516 1133
rect -3708 1093 -3696 1127
rect -3528 1093 -3516 1127
rect -3708 1087 -3516 1093
rect -3450 1127 -3258 1133
rect -3450 1093 -3438 1127
rect -3270 1093 -3258 1127
rect -3450 1087 -3258 1093
rect -3192 1127 -3000 1133
rect -3192 1093 -3180 1127
rect -3012 1093 -3000 1127
rect -3192 1087 -3000 1093
rect -2934 1127 -2742 1133
rect -2934 1093 -2922 1127
rect -2754 1093 -2742 1127
rect -2934 1087 -2742 1093
rect -2676 1127 -2484 1133
rect -2676 1093 -2664 1127
rect -2496 1093 -2484 1127
rect -2676 1087 -2484 1093
rect -2418 1127 -2226 1133
rect -2418 1093 -2406 1127
rect -2238 1093 -2226 1127
rect -2418 1087 -2226 1093
rect -2160 1127 -1968 1133
rect -2160 1093 -2148 1127
rect -1980 1093 -1968 1127
rect -2160 1087 -1968 1093
rect -1902 1127 -1710 1133
rect -1902 1093 -1890 1127
rect -1722 1093 -1710 1127
rect -1902 1087 -1710 1093
rect -1644 1127 -1452 1133
rect -1644 1093 -1632 1127
rect -1464 1093 -1452 1127
rect -1644 1087 -1452 1093
rect -1386 1127 -1194 1133
rect -1386 1093 -1374 1127
rect -1206 1093 -1194 1127
rect -1386 1087 -1194 1093
rect -1128 1127 -936 1133
rect -1128 1093 -1116 1127
rect -948 1093 -936 1127
rect -1128 1087 -936 1093
rect -870 1127 -678 1133
rect -870 1093 -858 1127
rect -690 1093 -678 1127
rect -870 1087 -678 1093
rect -612 1127 -420 1133
rect -612 1093 -600 1127
rect -432 1093 -420 1127
rect -612 1087 -420 1093
rect -354 1127 -162 1133
rect -354 1093 -342 1127
rect -174 1093 -162 1127
rect -354 1087 -162 1093
rect -96 1127 96 1133
rect -96 1093 -84 1127
rect 84 1093 96 1127
rect -96 1087 96 1093
rect 162 1127 354 1133
rect 162 1093 174 1127
rect 342 1093 354 1127
rect 162 1087 354 1093
rect 420 1127 612 1133
rect 420 1093 432 1127
rect 600 1093 612 1127
rect 420 1087 612 1093
rect 678 1127 870 1133
rect 678 1093 690 1127
rect 858 1093 870 1127
rect 678 1087 870 1093
rect 936 1127 1128 1133
rect 936 1093 948 1127
rect 1116 1093 1128 1127
rect 936 1087 1128 1093
rect 1194 1127 1386 1133
rect 1194 1093 1206 1127
rect 1374 1093 1386 1127
rect 1194 1087 1386 1093
rect 1452 1127 1644 1133
rect 1452 1093 1464 1127
rect 1632 1093 1644 1127
rect 1452 1087 1644 1093
rect 1710 1127 1902 1133
rect 1710 1093 1722 1127
rect 1890 1093 1902 1127
rect 1710 1087 1902 1093
rect 1968 1127 2160 1133
rect 1968 1093 1980 1127
rect 2148 1093 2160 1127
rect 1968 1087 2160 1093
rect 2226 1127 2418 1133
rect 2226 1093 2238 1127
rect 2406 1093 2418 1127
rect 2226 1087 2418 1093
rect 2484 1127 2676 1133
rect 2484 1093 2496 1127
rect 2664 1093 2676 1127
rect 2484 1087 2676 1093
rect 2742 1127 2934 1133
rect 2742 1093 2754 1127
rect 2922 1093 2934 1127
rect 2742 1087 2934 1093
rect 3000 1127 3192 1133
rect 3000 1093 3012 1127
rect 3180 1093 3192 1127
rect 3000 1087 3192 1093
rect 3258 1127 3450 1133
rect 3258 1093 3270 1127
rect 3438 1093 3450 1127
rect 3258 1087 3450 1093
rect 3516 1127 3708 1133
rect 3516 1093 3528 1127
rect 3696 1093 3708 1127
rect 3516 1087 3708 1093
rect 3774 1127 3966 1133
rect 3774 1093 3786 1127
rect 3954 1093 3966 1127
rect 3774 1087 3966 1093
rect 4032 1127 4224 1133
rect 4032 1093 4044 1127
rect 4212 1093 4224 1127
rect 4032 1087 4224 1093
rect 4290 1127 4482 1133
rect 4290 1093 4302 1127
rect 4470 1093 4482 1127
rect 4290 1087 4482 1093
rect 4548 1127 4740 1133
rect 4548 1093 4560 1127
rect 4728 1093 4740 1127
rect 4548 1087 4740 1093
rect 4806 1127 4998 1133
rect 4806 1093 4818 1127
rect 4986 1093 4998 1127
rect 4806 1087 4998 1093
rect 5064 1127 5256 1133
rect 5064 1093 5076 1127
rect 5244 1093 5256 1127
rect 5064 1087 5256 1093
rect 5322 1127 5514 1133
rect 5322 1093 5334 1127
rect 5502 1093 5514 1127
rect 5322 1087 5514 1093
rect 5580 1127 5772 1133
rect 5580 1093 5592 1127
rect 5760 1093 5772 1127
rect 5580 1087 5772 1093
rect 5838 1127 6030 1133
rect 5838 1093 5850 1127
rect 6018 1093 6030 1127
rect 5838 1087 6030 1093
rect 6096 1127 6288 1133
rect 6096 1093 6108 1127
rect 6276 1093 6288 1127
rect 6096 1087 6288 1093
rect 6354 1127 6546 1133
rect 6354 1093 6366 1127
rect 6534 1093 6546 1127
rect 6354 1087 6546 1093
rect 6612 1127 6804 1133
rect 6612 1093 6624 1127
rect 6792 1093 6804 1127
rect 6612 1087 6804 1093
rect 6870 1127 7062 1133
rect 6870 1093 6882 1127
rect 7050 1093 7062 1127
rect 6870 1087 7062 1093
rect -7118 1043 -7072 1055
rect -7118 67 -7112 1043
rect -7078 67 -7072 1043
rect -7118 55 -7072 67
rect -6860 1043 -6814 1055
rect -6860 67 -6854 1043
rect -6820 67 -6814 1043
rect -6860 55 -6814 67
rect -6602 1043 -6556 1055
rect -6602 67 -6596 1043
rect -6562 67 -6556 1043
rect -6602 55 -6556 67
rect -6344 1043 -6298 1055
rect -6344 67 -6338 1043
rect -6304 67 -6298 1043
rect -6344 55 -6298 67
rect -6086 1043 -6040 1055
rect -6086 67 -6080 1043
rect -6046 67 -6040 1043
rect -6086 55 -6040 67
rect -5828 1043 -5782 1055
rect -5828 67 -5822 1043
rect -5788 67 -5782 1043
rect -5828 55 -5782 67
rect -5570 1043 -5524 1055
rect -5570 67 -5564 1043
rect -5530 67 -5524 1043
rect -5570 55 -5524 67
rect -5312 1043 -5266 1055
rect -5312 67 -5306 1043
rect -5272 67 -5266 1043
rect -5312 55 -5266 67
rect -5054 1043 -5008 1055
rect -5054 67 -5048 1043
rect -5014 67 -5008 1043
rect -5054 55 -5008 67
rect -4796 1043 -4750 1055
rect -4796 67 -4790 1043
rect -4756 67 -4750 1043
rect -4796 55 -4750 67
rect -4538 1043 -4492 1055
rect -4538 67 -4532 1043
rect -4498 67 -4492 1043
rect -4538 55 -4492 67
rect -4280 1043 -4234 1055
rect -4280 67 -4274 1043
rect -4240 67 -4234 1043
rect -4280 55 -4234 67
rect -4022 1043 -3976 1055
rect -4022 67 -4016 1043
rect -3982 67 -3976 1043
rect -4022 55 -3976 67
rect -3764 1043 -3718 1055
rect -3764 67 -3758 1043
rect -3724 67 -3718 1043
rect -3764 55 -3718 67
rect -3506 1043 -3460 1055
rect -3506 67 -3500 1043
rect -3466 67 -3460 1043
rect -3506 55 -3460 67
rect -3248 1043 -3202 1055
rect -3248 67 -3242 1043
rect -3208 67 -3202 1043
rect -3248 55 -3202 67
rect -2990 1043 -2944 1055
rect -2990 67 -2984 1043
rect -2950 67 -2944 1043
rect -2990 55 -2944 67
rect -2732 1043 -2686 1055
rect -2732 67 -2726 1043
rect -2692 67 -2686 1043
rect -2732 55 -2686 67
rect -2474 1043 -2428 1055
rect -2474 67 -2468 1043
rect -2434 67 -2428 1043
rect -2474 55 -2428 67
rect -2216 1043 -2170 1055
rect -2216 67 -2210 1043
rect -2176 67 -2170 1043
rect -2216 55 -2170 67
rect -1958 1043 -1912 1055
rect -1958 67 -1952 1043
rect -1918 67 -1912 1043
rect -1958 55 -1912 67
rect -1700 1043 -1654 1055
rect -1700 67 -1694 1043
rect -1660 67 -1654 1043
rect -1700 55 -1654 67
rect -1442 1043 -1396 1055
rect -1442 67 -1436 1043
rect -1402 67 -1396 1043
rect -1442 55 -1396 67
rect -1184 1043 -1138 1055
rect -1184 67 -1178 1043
rect -1144 67 -1138 1043
rect -1184 55 -1138 67
rect -926 1043 -880 1055
rect -926 67 -920 1043
rect -886 67 -880 1043
rect -926 55 -880 67
rect -668 1043 -622 1055
rect -668 67 -662 1043
rect -628 67 -622 1043
rect -668 55 -622 67
rect -410 1043 -364 1055
rect -410 67 -404 1043
rect -370 67 -364 1043
rect -410 55 -364 67
rect -152 1043 -106 1055
rect -152 67 -146 1043
rect -112 67 -106 1043
rect -152 55 -106 67
rect 106 1043 152 1055
rect 106 67 112 1043
rect 146 67 152 1043
rect 106 55 152 67
rect 364 1043 410 1055
rect 364 67 370 1043
rect 404 67 410 1043
rect 364 55 410 67
rect 622 1043 668 1055
rect 622 67 628 1043
rect 662 67 668 1043
rect 622 55 668 67
rect 880 1043 926 1055
rect 880 67 886 1043
rect 920 67 926 1043
rect 880 55 926 67
rect 1138 1043 1184 1055
rect 1138 67 1144 1043
rect 1178 67 1184 1043
rect 1138 55 1184 67
rect 1396 1043 1442 1055
rect 1396 67 1402 1043
rect 1436 67 1442 1043
rect 1396 55 1442 67
rect 1654 1043 1700 1055
rect 1654 67 1660 1043
rect 1694 67 1700 1043
rect 1654 55 1700 67
rect 1912 1043 1958 1055
rect 1912 67 1918 1043
rect 1952 67 1958 1043
rect 1912 55 1958 67
rect 2170 1043 2216 1055
rect 2170 67 2176 1043
rect 2210 67 2216 1043
rect 2170 55 2216 67
rect 2428 1043 2474 1055
rect 2428 67 2434 1043
rect 2468 67 2474 1043
rect 2428 55 2474 67
rect 2686 1043 2732 1055
rect 2686 67 2692 1043
rect 2726 67 2732 1043
rect 2686 55 2732 67
rect 2944 1043 2990 1055
rect 2944 67 2950 1043
rect 2984 67 2990 1043
rect 2944 55 2990 67
rect 3202 1043 3248 1055
rect 3202 67 3208 1043
rect 3242 67 3248 1043
rect 3202 55 3248 67
rect 3460 1043 3506 1055
rect 3460 67 3466 1043
rect 3500 67 3506 1043
rect 3460 55 3506 67
rect 3718 1043 3764 1055
rect 3718 67 3724 1043
rect 3758 67 3764 1043
rect 3718 55 3764 67
rect 3976 1043 4022 1055
rect 3976 67 3982 1043
rect 4016 67 4022 1043
rect 3976 55 4022 67
rect 4234 1043 4280 1055
rect 4234 67 4240 1043
rect 4274 67 4280 1043
rect 4234 55 4280 67
rect 4492 1043 4538 1055
rect 4492 67 4498 1043
rect 4532 67 4538 1043
rect 4492 55 4538 67
rect 4750 1043 4796 1055
rect 4750 67 4756 1043
rect 4790 67 4796 1043
rect 4750 55 4796 67
rect 5008 1043 5054 1055
rect 5008 67 5014 1043
rect 5048 67 5054 1043
rect 5008 55 5054 67
rect 5266 1043 5312 1055
rect 5266 67 5272 1043
rect 5306 67 5312 1043
rect 5266 55 5312 67
rect 5524 1043 5570 1055
rect 5524 67 5530 1043
rect 5564 67 5570 1043
rect 5524 55 5570 67
rect 5782 1043 5828 1055
rect 5782 67 5788 1043
rect 5822 67 5828 1043
rect 5782 55 5828 67
rect 6040 1043 6086 1055
rect 6040 67 6046 1043
rect 6080 67 6086 1043
rect 6040 55 6086 67
rect 6298 1043 6344 1055
rect 6298 67 6304 1043
rect 6338 67 6344 1043
rect 6298 55 6344 67
rect 6556 1043 6602 1055
rect 6556 67 6562 1043
rect 6596 67 6602 1043
rect 6556 55 6602 67
rect 6814 1043 6860 1055
rect 6814 67 6820 1043
rect 6854 67 6860 1043
rect 6814 55 6860 67
rect 7072 1043 7118 1055
rect 7072 67 7078 1043
rect 7112 67 7118 1043
rect 7072 55 7118 67
rect -7062 17 -6870 23
rect -7062 -17 -7050 17
rect -6882 -17 -6870 17
rect -7062 -23 -6870 -17
rect -6804 17 -6612 23
rect -6804 -17 -6792 17
rect -6624 -17 -6612 17
rect -6804 -23 -6612 -17
rect -6546 17 -6354 23
rect -6546 -17 -6534 17
rect -6366 -17 -6354 17
rect -6546 -23 -6354 -17
rect -6288 17 -6096 23
rect -6288 -17 -6276 17
rect -6108 -17 -6096 17
rect -6288 -23 -6096 -17
rect -6030 17 -5838 23
rect -6030 -17 -6018 17
rect -5850 -17 -5838 17
rect -6030 -23 -5838 -17
rect -5772 17 -5580 23
rect -5772 -17 -5760 17
rect -5592 -17 -5580 17
rect -5772 -23 -5580 -17
rect -5514 17 -5322 23
rect -5514 -17 -5502 17
rect -5334 -17 -5322 17
rect -5514 -23 -5322 -17
rect -5256 17 -5064 23
rect -5256 -17 -5244 17
rect -5076 -17 -5064 17
rect -5256 -23 -5064 -17
rect -4998 17 -4806 23
rect -4998 -17 -4986 17
rect -4818 -17 -4806 17
rect -4998 -23 -4806 -17
rect -4740 17 -4548 23
rect -4740 -17 -4728 17
rect -4560 -17 -4548 17
rect -4740 -23 -4548 -17
rect -4482 17 -4290 23
rect -4482 -17 -4470 17
rect -4302 -17 -4290 17
rect -4482 -23 -4290 -17
rect -4224 17 -4032 23
rect -4224 -17 -4212 17
rect -4044 -17 -4032 17
rect -4224 -23 -4032 -17
rect -3966 17 -3774 23
rect -3966 -17 -3954 17
rect -3786 -17 -3774 17
rect -3966 -23 -3774 -17
rect -3708 17 -3516 23
rect -3708 -17 -3696 17
rect -3528 -17 -3516 17
rect -3708 -23 -3516 -17
rect -3450 17 -3258 23
rect -3450 -17 -3438 17
rect -3270 -17 -3258 17
rect -3450 -23 -3258 -17
rect -3192 17 -3000 23
rect -3192 -17 -3180 17
rect -3012 -17 -3000 17
rect -3192 -23 -3000 -17
rect -2934 17 -2742 23
rect -2934 -17 -2922 17
rect -2754 -17 -2742 17
rect -2934 -23 -2742 -17
rect -2676 17 -2484 23
rect -2676 -17 -2664 17
rect -2496 -17 -2484 17
rect -2676 -23 -2484 -17
rect -2418 17 -2226 23
rect -2418 -17 -2406 17
rect -2238 -17 -2226 17
rect -2418 -23 -2226 -17
rect -2160 17 -1968 23
rect -2160 -17 -2148 17
rect -1980 -17 -1968 17
rect -2160 -23 -1968 -17
rect -1902 17 -1710 23
rect -1902 -17 -1890 17
rect -1722 -17 -1710 17
rect -1902 -23 -1710 -17
rect -1644 17 -1452 23
rect -1644 -17 -1632 17
rect -1464 -17 -1452 17
rect -1644 -23 -1452 -17
rect -1386 17 -1194 23
rect -1386 -17 -1374 17
rect -1206 -17 -1194 17
rect -1386 -23 -1194 -17
rect -1128 17 -936 23
rect -1128 -17 -1116 17
rect -948 -17 -936 17
rect -1128 -23 -936 -17
rect -870 17 -678 23
rect -870 -17 -858 17
rect -690 -17 -678 17
rect -870 -23 -678 -17
rect -612 17 -420 23
rect -612 -17 -600 17
rect -432 -17 -420 17
rect -612 -23 -420 -17
rect -354 17 -162 23
rect -354 -17 -342 17
rect -174 -17 -162 17
rect -354 -23 -162 -17
rect -96 17 96 23
rect -96 -17 -84 17
rect 84 -17 96 17
rect -96 -23 96 -17
rect 162 17 354 23
rect 162 -17 174 17
rect 342 -17 354 17
rect 162 -23 354 -17
rect 420 17 612 23
rect 420 -17 432 17
rect 600 -17 612 17
rect 420 -23 612 -17
rect 678 17 870 23
rect 678 -17 690 17
rect 858 -17 870 17
rect 678 -23 870 -17
rect 936 17 1128 23
rect 936 -17 948 17
rect 1116 -17 1128 17
rect 936 -23 1128 -17
rect 1194 17 1386 23
rect 1194 -17 1206 17
rect 1374 -17 1386 17
rect 1194 -23 1386 -17
rect 1452 17 1644 23
rect 1452 -17 1464 17
rect 1632 -17 1644 17
rect 1452 -23 1644 -17
rect 1710 17 1902 23
rect 1710 -17 1722 17
rect 1890 -17 1902 17
rect 1710 -23 1902 -17
rect 1968 17 2160 23
rect 1968 -17 1980 17
rect 2148 -17 2160 17
rect 1968 -23 2160 -17
rect 2226 17 2418 23
rect 2226 -17 2238 17
rect 2406 -17 2418 17
rect 2226 -23 2418 -17
rect 2484 17 2676 23
rect 2484 -17 2496 17
rect 2664 -17 2676 17
rect 2484 -23 2676 -17
rect 2742 17 2934 23
rect 2742 -17 2754 17
rect 2922 -17 2934 17
rect 2742 -23 2934 -17
rect 3000 17 3192 23
rect 3000 -17 3012 17
rect 3180 -17 3192 17
rect 3000 -23 3192 -17
rect 3258 17 3450 23
rect 3258 -17 3270 17
rect 3438 -17 3450 17
rect 3258 -23 3450 -17
rect 3516 17 3708 23
rect 3516 -17 3528 17
rect 3696 -17 3708 17
rect 3516 -23 3708 -17
rect 3774 17 3966 23
rect 3774 -17 3786 17
rect 3954 -17 3966 17
rect 3774 -23 3966 -17
rect 4032 17 4224 23
rect 4032 -17 4044 17
rect 4212 -17 4224 17
rect 4032 -23 4224 -17
rect 4290 17 4482 23
rect 4290 -17 4302 17
rect 4470 -17 4482 17
rect 4290 -23 4482 -17
rect 4548 17 4740 23
rect 4548 -17 4560 17
rect 4728 -17 4740 17
rect 4548 -23 4740 -17
rect 4806 17 4998 23
rect 4806 -17 4818 17
rect 4986 -17 4998 17
rect 4806 -23 4998 -17
rect 5064 17 5256 23
rect 5064 -17 5076 17
rect 5244 -17 5256 17
rect 5064 -23 5256 -17
rect 5322 17 5514 23
rect 5322 -17 5334 17
rect 5502 -17 5514 17
rect 5322 -23 5514 -17
rect 5580 17 5772 23
rect 5580 -17 5592 17
rect 5760 -17 5772 17
rect 5580 -23 5772 -17
rect 5838 17 6030 23
rect 5838 -17 5850 17
rect 6018 -17 6030 17
rect 5838 -23 6030 -17
rect 6096 17 6288 23
rect 6096 -17 6108 17
rect 6276 -17 6288 17
rect 6096 -23 6288 -17
rect 6354 17 6546 23
rect 6354 -17 6366 17
rect 6534 -17 6546 17
rect 6354 -23 6546 -17
rect 6612 17 6804 23
rect 6612 -17 6624 17
rect 6792 -17 6804 17
rect 6612 -23 6804 -17
rect 6870 17 7062 23
rect 6870 -17 6882 17
rect 7050 -17 7062 17
rect 6870 -23 7062 -17
rect -7118 -67 -7072 -55
rect -7118 -1043 -7112 -67
rect -7078 -1043 -7072 -67
rect -7118 -1055 -7072 -1043
rect -6860 -67 -6814 -55
rect -6860 -1043 -6854 -67
rect -6820 -1043 -6814 -67
rect -6860 -1055 -6814 -1043
rect -6602 -67 -6556 -55
rect -6602 -1043 -6596 -67
rect -6562 -1043 -6556 -67
rect -6602 -1055 -6556 -1043
rect -6344 -67 -6298 -55
rect -6344 -1043 -6338 -67
rect -6304 -1043 -6298 -67
rect -6344 -1055 -6298 -1043
rect -6086 -67 -6040 -55
rect -6086 -1043 -6080 -67
rect -6046 -1043 -6040 -67
rect -6086 -1055 -6040 -1043
rect -5828 -67 -5782 -55
rect -5828 -1043 -5822 -67
rect -5788 -1043 -5782 -67
rect -5828 -1055 -5782 -1043
rect -5570 -67 -5524 -55
rect -5570 -1043 -5564 -67
rect -5530 -1043 -5524 -67
rect -5570 -1055 -5524 -1043
rect -5312 -67 -5266 -55
rect -5312 -1043 -5306 -67
rect -5272 -1043 -5266 -67
rect -5312 -1055 -5266 -1043
rect -5054 -67 -5008 -55
rect -5054 -1043 -5048 -67
rect -5014 -1043 -5008 -67
rect -5054 -1055 -5008 -1043
rect -4796 -67 -4750 -55
rect -4796 -1043 -4790 -67
rect -4756 -1043 -4750 -67
rect -4796 -1055 -4750 -1043
rect -4538 -67 -4492 -55
rect -4538 -1043 -4532 -67
rect -4498 -1043 -4492 -67
rect -4538 -1055 -4492 -1043
rect -4280 -67 -4234 -55
rect -4280 -1043 -4274 -67
rect -4240 -1043 -4234 -67
rect -4280 -1055 -4234 -1043
rect -4022 -67 -3976 -55
rect -4022 -1043 -4016 -67
rect -3982 -1043 -3976 -67
rect -4022 -1055 -3976 -1043
rect -3764 -67 -3718 -55
rect -3764 -1043 -3758 -67
rect -3724 -1043 -3718 -67
rect -3764 -1055 -3718 -1043
rect -3506 -67 -3460 -55
rect -3506 -1043 -3500 -67
rect -3466 -1043 -3460 -67
rect -3506 -1055 -3460 -1043
rect -3248 -67 -3202 -55
rect -3248 -1043 -3242 -67
rect -3208 -1043 -3202 -67
rect -3248 -1055 -3202 -1043
rect -2990 -67 -2944 -55
rect -2990 -1043 -2984 -67
rect -2950 -1043 -2944 -67
rect -2990 -1055 -2944 -1043
rect -2732 -67 -2686 -55
rect -2732 -1043 -2726 -67
rect -2692 -1043 -2686 -67
rect -2732 -1055 -2686 -1043
rect -2474 -67 -2428 -55
rect -2474 -1043 -2468 -67
rect -2434 -1043 -2428 -67
rect -2474 -1055 -2428 -1043
rect -2216 -67 -2170 -55
rect -2216 -1043 -2210 -67
rect -2176 -1043 -2170 -67
rect -2216 -1055 -2170 -1043
rect -1958 -67 -1912 -55
rect -1958 -1043 -1952 -67
rect -1918 -1043 -1912 -67
rect -1958 -1055 -1912 -1043
rect -1700 -67 -1654 -55
rect -1700 -1043 -1694 -67
rect -1660 -1043 -1654 -67
rect -1700 -1055 -1654 -1043
rect -1442 -67 -1396 -55
rect -1442 -1043 -1436 -67
rect -1402 -1043 -1396 -67
rect -1442 -1055 -1396 -1043
rect -1184 -67 -1138 -55
rect -1184 -1043 -1178 -67
rect -1144 -1043 -1138 -67
rect -1184 -1055 -1138 -1043
rect -926 -67 -880 -55
rect -926 -1043 -920 -67
rect -886 -1043 -880 -67
rect -926 -1055 -880 -1043
rect -668 -67 -622 -55
rect -668 -1043 -662 -67
rect -628 -1043 -622 -67
rect -668 -1055 -622 -1043
rect -410 -67 -364 -55
rect -410 -1043 -404 -67
rect -370 -1043 -364 -67
rect -410 -1055 -364 -1043
rect -152 -67 -106 -55
rect -152 -1043 -146 -67
rect -112 -1043 -106 -67
rect -152 -1055 -106 -1043
rect 106 -67 152 -55
rect 106 -1043 112 -67
rect 146 -1043 152 -67
rect 106 -1055 152 -1043
rect 364 -67 410 -55
rect 364 -1043 370 -67
rect 404 -1043 410 -67
rect 364 -1055 410 -1043
rect 622 -67 668 -55
rect 622 -1043 628 -67
rect 662 -1043 668 -67
rect 622 -1055 668 -1043
rect 880 -67 926 -55
rect 880 -1043 886 -67
rect 920 -1043 926 -67
rect 880 -1055 926 -1043
rect 1138 -67 1184 -55
rect 1138 -1043 1144 -67
rect 1178 -1043 1184 -67
rect 1138 -1055 1184 -1043
rect 1396 -67 1442 -55
rect 1396 -1043 1402 -67
rect 1436 -1043 1442 -67
rect 1396 -1055 1442 -1043
rect 1654 -67 1700 -55
rect 1654 -1043 1660 -67
rect 1694 -1043 1700 -67
rect 1654 -1055 1700 -1043
rect 1912 -67 1958 -55
rect 1912 -1043 1918 -67
rect 1952 -1043 1958 -67
rect 1912 -1055 1958 -1043
rect 2170 -67 2216 -55
rect 2170 -1043 2176 -67
rect 2210 -1043 2216 -67
rect 2170 -1055 2216 -1043
rect 2428 -67 2474 -55
rect 2428 -1043 2434 -67
rect 2468 -1043 2474 -67
rect 2428 -1055 2474 -1043
rect 2686 -67 2732 -55
rect 2686 -1043 2692 -67
rect 2726 -1043 2732 -67
rect 2686 -1055 2732 -1043
rect 2944 -67 2990 -55
rect 2944 -1043 2950 -67
rect 2984 -1043 2990 -67
rect 2944 -1055 2990 -1043
rect 3202 -67 3248 -55
rect 3202 -1043 3208 -67
rect 3242 -1043 3248 -67
rect 3202 -1055 3248 -1043
rect 3460 -67 3506 -55
rect 3460 -1043 3466 -67
rect 3500 -1043 3506 -67
rect 3460 -1055 3506 -1043
rect 3718 -67 3764 -55
rect 3718 -1043 3724 -67
rect 3758 -1043 3764 -67
rect 3718 -1055 3764 -1043
rect 3976 -67 4022 -55
rect 3976 -1043 3982 -67
rect 4016 -1043 4022 -67
rect 3976 -1055 4022 -1043
rect 4234 -67 4280 -55
rect 4234 -1043 4240 -67
rect 4274 -1043 4280 -67
rect 4234 -1055 4280 -1043
rect 4492 -67 4538 -55
rect 4492 -1043 4498 -67
rect 4532 -1043 4538 -67
rect 4492 -1055 4538 -1043
rect 4750 -67 4796 -55
rect 4750 -1043 4756 -67
rect 4790 -1043 4796 -67
rect 4750 -1055 4796 -1043
rect 5008 -67 5054 -55
rect 5008 -1043 5014 -67
rect 5048 -1043 5054 -67
rect 5008 -1055 5054 -1043
rect 5266 -67 5312 -55
rect 5266 -1043 5272 -67
rect 5306 -1043 5312 -67
rect 5266 -1055 5312 -1043
rect 5524 -67 5570 -55
rect 5524 -1043 5530 -67
rect 5564 -1043 5570 -67
rect 5524 -1055 5570 -1043
rect 5782 -67 5828 -55
rect 5782 -1043 5788 -67
rect 5822 -1043 5828 -67
rect 5782 -1055 5828 -1043
rect 6040 -67 6086 -55
rect 6040 -1043 6046 -67
rect 6080 -1043 6086 -67
rect 6040 -1055 6086 -1043
rect 6298 -67 6344 -55
rect 6298 -1043 6304 -67
rect 6338 -1043 6344 -67
rect 6298 -1055 6344 -1043
rect 6556 -67 6602 -55
rect 6556 -1043 6562 -67
rect 6596 -1043 6602 -67
rect 6556 -1055 6602 -1043
rect 6814 -67 6860 -55
rect 6814 -1043 6820 -67
rect 6854 -1043 6860 -67
rect 6814 -1055 6860 -1043
rect 7072 -67 7118 -55
rect 7072 -1043 7078 -67
rect 7112 -1043 7118 -67
rect 7072 -1055 7118 -1043
rect -7062 -1093 -6870 -1087
rect -7062 -1127 -7050 -1093
rect -6882 -1127 -6870 -1093
rect -7062 -1133 -6870 -1127
rect -6804 -1093 -6612 -1087
rect -6804 -1127 -6792 -1093
rect -6624 -1127 -6612 -1093
rect -6804 -1133 -6612 -1127
rect -6546 -1093 -6354 -1087
rect -6546 -1127 -6534 -1093
rect -6366 -1127 -6354 -1093
rect -6546 -1133 -6354 -1127
rect -6288 -1093 -6096 -1087
rect -6288 -1127 -6276 -1093
rect -6108 -1127 -6096 -1093
rect -6288 -1133 -6096 -1127
rect -6030 -1093 -5838 -1087
rect -6030 -1127 -6018 -1093
rect -5850 -1127 -5838 -1093
rect -6030 -1133 -5838 -1127
rect -5772 -1093 -5580 -1087
rect -5772 -1127 -5760 -1093
rect -5592 -1127 -5580 -1093
rect -5772 -1133 -5580 -1127
rect -5514 -1093 -5322 -1087
rect -5514 -1127 -5502 -1093
rect -5334 -1127 -5322 -1093
rect -5514 -1133 -5322 -1127
rect -5256 -1093 -5064 -1087
rect -5256 -1127 -5244 -1093
rect -5076 -1127 -5064 -1093
rect -5256 -1133 -5064 -1127
rect -4998 -1093 -4806 -1087
rect -4998 -1127 -4986 -1093
rect -4818 -1127 -4806 -1093
rect -4998 -1133 -4806 -1127
rect -4740 -1093 -4548 -1087
rect -4740 -1127 -4728 -1093
rect -4560 -1127 -4548 -1093
rect -4740 -1133 -4548 -1127
rect -4482 -1093 -4290 -1087
rect -4482 -1127 -4470 -1093
rect -4302 -1127 -4290 -1093
rect -4482 -1133 -4290 -1127
rect -4224 -1093 -4032 -1087
rect -4224 -1127 -4212 -1093
rect -4044 -1127 -4032 -1093
rect -4224 -1133 -4032 -1127
rect -3966 -1093 -3774 -1087
rect -3966 -1127 -3954 -1093
rect -3786 -1127 -3774 -1093
rect -3966 -1133 -3774 -1127
rect -3708 -1093 -3516 -1087
rect -3708 -1127 -3696 -1093
rect -3528 -1127 -3516 -1093
rect -3708 -1133 -3516 -1127
rect -3450 -1093 -3258 -1087
rect -3450 -1127 -3438 -1093
rect -3270 -1127 -3258 -1093
rect -3450 -1133 -3258 -1127
rect -3192 -1093 -3000 -1087
rect -3192 -1127 -3180 -1093
rect -3012 -1127 -3000 -1093
rect -3192 -1133 -3000 -1127
rect -2934 -1093 -2742 -1087
rect -2934 -1127 -2922 -1093
rect -2754 -1127 -2742 -1093
rect -2934 -1133 -2742 -1127
rect -2676 -1093 -2484 -1087
rect -2676 -1127 -2664 -1093
rect -2496 -1127 -2484 -1093
rect -2676 -1133 -2484 -1127
rect -2418 -1093 -2226 -1087
rect -2418 -1127 -2406 -1093
rect -2238 -1127 -2226 -1093
rect -2418 -1133 -2226 -1127
rect -2160 -1093 -1968 -1087
rect -2160 -1127 -2148 -1093
rect -1980 -1127 -1968 -1093
rect -2160 -1133 -1968 -1127
rect -1902 -1093 -1710 -1087
rect -1902 -1127 -1890 -1093
rect -1722 -1127 -1710 -1093
rect -1902 -1133 -1710 -1127
rect -1644 -1093 -1452 -1087
rect -1644 -1127 -1632 -1093
rect -1464 -1127 -1452 -1093
rect -1644 -1133 -1452 -1127
rect -1386 -1093 -1194 -1087
rect -1386 -1127 -1374 -1093
rect -1206 -1127 -1194 -1093
rect -1386 -1133 -1194 -1127
rect -1128 -1093 -936 -1087
rect -1128 -1127 -1116 -1093
rect -948 -1127 -936 -1093
rect -1128 -1133 -936 -1127
rect -870 -1093 -678 -1087
rect -870 -1127 -858 -1093
rect -690 -1127 -678 -1093
rect -870 -1133 -678 -1127
rect -612 -1093 -420 -1087
rect -612 -1127 -600 -1093
rect -432 -1127 -420 -1093
rect -612 -1133 -420 -1127
rect -354 -1093 -162 -1087
rect -354 -1127 -342 -1093
rect -174 -1127 -162 -1093
rect -354 -1133 -162 -1127
rect -96 -1093 96 -1087
rect -96 -1127 -84 -1093
rect 84 -1127 96 -1093
rect -96 -1133 96 -1127
rect 162 -1093 354 -1087
rect 162 -1127 174 -1093
rect 342 -1127 354 -1093
rect 162 -1133 354 -1127
rect 420 -1093 612 -1087
rect 420 -1127 432 -1093
rect 600 -1127 612 -1093
rect 420 -1133 612 -1127
rect 678 -1093 870 -1087
rect 678 -1127 690 -1093
rect 858 -1127 870 -1093
rect 678 -1133 870 -1127
rect 936 -1093 1128 -1087
rect 936 -1127 948 -1093
rect 1116 -1127 1128 -1093
rect 936 -1133 1128 -1127
rect 1194 -1093 1386 -1087
rect 1194 -1127 1206 -1093
rect 1374 -1127 1386 -1093
rect 1194 -1133 1386 -1127
rect 1452 -1093 1644 -1087
rect 1452 -1127 1464 -1093
rect 1632 -1127 1644 -1093
rect 1452 -1133 1644 -1127
rect 1710 -1093 1902 -1087
rect 1710 -1127 1722 -1093
rect 1890 -1127 1902 -1093
rect 1710 -1133 1902 -1127
rect 1968 -1093 2160 -1087
rect 1968 -1127 1980 -1093
rect 2148 -1127 2160 -1093
rect 1968 -1133 2160 -1127
rect 2226 -1093 2418 -1087
rect 2226 -1127 2238 -1093
rect 2406 -1127 2418 -1093
rect 2226 -1133 2418 -1127
rect 2484 -1093 2676 -1087
rect 2484 -1127 2496 -1093
rect 2664 -1127 2676 -1093
rect 2484 -1133 2676 -1127
rect 2742 -1093 2934 -1087
rect 2742 -1127 2754 -1093
rect 2922 -1127 2934 -1093
rect 2742 -1133 2934 -1127
rect 3000 -1093 3192 -1087
rect 3000 -1127 3012 -1093
rect 3180 -1127 3192 -1093
rect 3000 -1133 3192 -1127
rect 3258 -1093 3450 -1087
rect 3258 -1127 3270 -1093
rect 3438 -1127 3450 -1093
rect 3258 -1133 3450 -1127
rect 3516 -1093 3708 -1087
rect 3516 -1127 3528 -1093
rect 3696 -1127 3708 -1093
rect 3516 -1133 3708 -1127
rect 3774 -1093 3966 -1087
rect 3774 -1127 3786 -1093
rect 3954 -1127 3966 -1093
rect 3774 -1133 3966 -1127
rect 4032 -1093 4224 -1087
rect 4032 -1127 4044 -1093
rect 4212 -1127 4224 -1093
rect 4032 -1133 4224 -1127
rect 4290 -1093 4482 -1087
rect 4290 -1127 4302 -1093
rect 4470 -1127 4482 -1093
rect 4290 -1133 4482 -1127
rect 4548 -1093 4740 -1087
rect 4548 -1127 4560 -1093
rect 4728 -1127 4740 -1093
rect 4548 -1133 4740 -1127
rect 4806 -1093 4998 -1087
rect 4806 -1127 4818 -1093
rect 4986 -1127 4998 -1093
rect 4806 -1133 4998 -1127
rect 5064 -1093 5256 -1087
rect 5064 -1127 5076 -1093
rect 5244 -1127 5256 -1093
rect 5064 -1133 5256 -1127
rect 5322 -1093 5514 -1087
rect 5322 -1127 5334 -1093
rect 5502 -1127 5514 -1093
rect 5322 -1133 5514 -1127
rect 5580 -1093 5772 -1087
rect 5580 -1127 5592 -1093
rect 5760 -1127 5772 -1093
rect 5580 -1133 5772 -1127
rect 5838 -1093 6030 -1087
rect 5838 -1127 5850 -1093
rect 6018 -1127 6030 -1093
rect 5838 -1133 6030 -1127
rect 6096 -1093 6288 -1087
rect 6096 -1127 6108 -1093
rect 6276 -1127 6288 -1093
rect 6096 -1133 6288 -1127
rect 6354 -1093 6546 -1087
rect 6354 -1127 6366 -1093
rect 6534 -1127 6546 -1093
rect 6354 -1133 6546 -1127
rect 6612 -1093 6804 -1087
rect 6612 -1127 6624 -1093
rect 6792 -1127 6804 -1093
rect 6612 -1133 6804 -1127
rect 6870 -1093 7062 -1087
rect 6870 -1127 6882 -1093
rect 7050 -1127 7062 -1093
rect 6870 -1133 7062 -1127
rect -7118 -1177 -7072 -1165
rect -7118 -2153 -7112 -1177
rect -7078 -2153 -7072 -1177
rect -7118 -2165 -7072 -2153
rect -6860 -1177 -6814 -1165
rect -6860 -2153 -6854 -1177
rect -6820 -2153 -6814 -1177
rect -6860 -2165 -6814 -2153
rect -6602 -1177 -6556 -1165
rect -6602 -2153 -6596 -1177
rect -6562 -2153 -6556 -1177
rect -6602 -2165 -6556 -2153
rect -6344 -1177 -6298 -1165
rect -6344 -2153 -6338 -1177
rect -6304 -2153 -6298 -1177
rect -6344 -2165 -6298 -2153
rect -6086 -1177 -6040 -1165
rect -6086 -2153 -6080 -1177
rect -6046 -2153 -6040 -1177
rect -6086 -2165 -6040 -2153
rect -5828 -1177 -5782 -1165
rect -5828 -2153 -5822 -1177
rect -5788 -2153 -5782 -1177
rect -5828 -2165 -5782 -2153
rect -5570 -1177 -5524 -1165
rect -5570 -2153 -5564 -1177
rect -5530 -2153 -5524 -1177
rect -5570 -2165 -5524 -2153
rect -5312 -1177 -5266 -1165
rect -5312 -2153 -5306 -1177
rect -5272 -2153 -5266 -1177
rect -5312 -2165 -5266 -2153
rect -5054 -1177 -5008 -1165
rect -5054 -2153 -5048 -1177
rect -5014 -2153 -5008 -1177
rect -5054 -2165 -5008 -2153
rect -4796 -1177 -4750 -1165
rect -4796 -2153 -4790 -1177
rect -4756 -2153 -4750 -1177
rect -4796 -2165 -4750 -2153
rect -4538 -1177 -4492 -1165
rect -4538 -2153 -4532 -1177
rect -4498 -2153 -4492 -1177
rect -4538 -2165 -4492 -2153
rect -4280 -1177 -4234 -1165
rect -4280 -2153 -4274 -1177
rect -4240 -2153 -4234 -1177
rect -4280 -2165 -4234 -2153
rect -4022 -1177 -3976 -1165
rect -4022 -2153 -4016 -1177
rect -3982 -2153 -3976 -1177
rect -4022 -2165 -3976 -2153
rect -3764 -1177 -3718 -1165
rect -3764 -2153 -3758 -1177
rect -3724 -2153 -3718 -1177
rect -3764 -2165 -3718 -2153
rect -3506 -1177 -3460 -1165
rect -3506 -2153 -3500 -1177
rect -3466 -2153 -3460 -1177
rect -3506 -2165 -3460 -2153
rect -3248 -1177 -3202 -1165
rect -3248 -2153 -3242 -1177
rect -3208 -2153 -3202 -1177
rect -3248 -2165 -3202 -2153
rect -2990 -1177 -2944 -1165
rect -2990 -2153 -2984 -1177
rect -2950 -2153 -2944 -1177
rect -2990 -2165 -2944 -2153
rect -2732 -1177 -2686 -1165
rect -2732 -2153 -2726 -1177
rect -2692 -2153 -2686 -1177
rect -2732 -2165 -2686 -2153
rect -2474 -1177 -2428 -1165
rect -2474 -2153 -2468 -1177
rect -2434 -2153 -2428 -1177
rect -2474 -2165 -2428 -2153
rect -2216 -1177 -2170 -1165
rect -2216 -2153 -2210 -1177
rect -2176 -2153 -2170 -1177
rect -2216 -2165 -2170 -2153
rect -1958 -1177 -1912 -1165
rect -1958 -2153 -1952 -1177
rect -1918 -2153 -1912 -1177
rect -1958 -2165 -1912 -2153
rect -1700 -1177 -1654 -1165
rect -1700 -2153 -1694 -1177
rect -1660 -2153 -1654 -1177
rect -1700 -2165 -1654 -2153
rect -1442 -1177 -1396 -1165
rect -1442 -2153 -1436 -1177
rect -1402 -2153 -1396 -1177
rect -1442 -2165 -1396 -2153
rect -1184 -1177 -1138 -1165
rect -1184 -2153 -1178 -1177
rect -1144 -2153 -1138 -1177
rect -1184 -2165 -1138 -2153
rect -926 -1177 -880 -1165
rect -926 -2153 -920 -1177
rect -886 -2153 -880 -1177
rect -926 -2165 -880 -2153
rect -668 -1177 -622 -1165
rect -668 -2153 -662 -1177
rect -628 -2153 -622 -1177
rect -668 -2165 -622 -2153
rect -410 -1177 -364 -1165
rect -410 -2153 -404 -1177
rect -370 -2153 -364 -1177
rect -410 -2165 -364 -2153
rect -152 -1177 -106 -1165
rect -152 -2153 -146 -1177
rect -112 -2153 -106 -1177
rect -152 -2165 -106 -2153
rect 106 -1177 152 -1165
rect 106 -2153 112 -1177
rect 146 -2153 152 -1177
rect 106 -2165 152 -2153
rect 364 -1177 410 -1165
rect 364 -2153 370 -1177
rect 404 -2153 410 -1177
rect 364 -2165 410 -2153
rect 622 -1177 668 -1165
rect 622 -2153 628 -1177
rect 662 -2153 668 -1177
rect 622 -2165 668 -2153
rect 880 -1177 926 -1165
rect 880 -2153 886 -1177
rect 920 -2153 926 -1177
rect 880 -2165 926 -2153
rect 1138 -1177 1184 -1165
rect 1138 -2153 1144 -1177
rect 1178 -2153 1184 -1177
rect 1138 -2165 1184 -2153
rect 1396 -1177 1442 -1165
rect 1396 -2153 1402 -1177
rect 1436 -2153 1442 -1177
rect 1396 -2165 1442 -2153
rect 1654 -1177 1700 -1165
rect 1654 -2153 1660 -1177
rect 1694 -2153 1700 -1177
rect 1654 -2165 1700 -2153
rect 1912 -1177 1958 -1165
rect 1912 -2153 1918 -1177
rect 1952 -2153 1958 -1177
rect 1912 -2165 1958 -2153
rect 2170 -1177 2216 -1165
rect 2170 -2153 2176 -1177
rect 2210 -2153 2216 -1177
rect 2170 -2165 2216 -2153
rect 2428 -1177 2474 -1165
rect 2428 -2153 2434 -1177
rect 2468 -2153 2474 -1177
rect 2428 -2165 2474 -2153
rect 2686 -1177 2732 -1165
rect 2686 -2153 2692 -1177
rect 2726 -2153 2732 -1177
rect 2686 -2165 2732 -2153
rect 2944 -1177 2990 -1165
rect 2944 -2153 2950 -1177
rect 2984 -2153 2990 -1177
rect 2944 -2165 2990 -2153
rect 3202 -1177 3248 -1165
rect 3202 -2153 3208 -1177
rect 3242 -2153 3248 -1177
rect 3202 -2165 3248 -2153
rect 3460 -1177 3506 -1165
rect 3460 -2153 3466 -1177
rect 3500 -2153 3506 -1177
rect 3460 -2165 3506 -2153
rect 3718 -1177 3764 -1165
rect 3718 -2153 3724 -1177
rect 3758 -2153 3764 -1177
rect 3718 -2165 3764 -2153
rect 3976 -1177 4022 -1165
rect 3976 -2153 3982 -1177
rect 4016 -2153 4022 -1177
rect 3976 -2165 4022 -2153
rect 4234 -1177 4280 -1165
rect 4234 -2153 4240 -1177
rect 4274 -2153 4280 -1177
rect 4234 -2165 4280 -2153
rect 4492 -1177 4538 -1165
rect 4492 -2153 4498 -1177
rect 4532 -2153 4538 -1177
rect 4492 -2165 4538 -2153
rect 4750 -1177 4796 -1165
rect 4750 -2153 4756 -1177
rect 4790 -2153 4796 -1177
rect 4750 -2165 4796 -2153
rect 5008 -1177 5054 -1165
rect 5008 -2153 5014 -1177
rect 5048 -2153 5054 -1177
rect 5008 -2165 5054 -2153
rect 5266 -1177 5312 -1165
rect 5266 -2153 5272 -1177
rect 5306 -2153 5312 -1177
rect 5266 -2165 5312 -2153
rect 5524 -1177 5570 -1165
rect 5524 -2153 5530 -1177
rect 5564 -2153 5570 -1177
rect 5524 -2165 5570 -2153
rect 5782 -1177 5828 -1165
rect 5782 -2153 5788 -1177
rect 5822 -2153 5828 -1177
rect 5782 -2165 5828 -2153
rect 6040 -1177 6086 -1165
rect 6040 -2153 6046 -1177
rect 6080 -2153 6086 -1177
rect 6040 -2165 6086 -2153
rect 6298 -1177 6344 -1165
rect 6298 -2153 6304 -1177
rect 6338 -2153 6344 -1177
rect 6298 -2165 6344 -2153
rect 6556 -1177 6602 -1165
rect 6556 -2153 6562 -1177
rect 6596 -2153 6602 -1177
rect 6556 -2165 6602 -2153
rect 6814 -1177 6860 -1165
rect 6814 -2153 6820 -1177
rect 6854 -2153 6860 -1177
rect 6814 -2165 6860 -2153
rect 7072 -1177 7118 -1165
rect 7072 -2153 7078 -1177
rect 7112 -2153 7118 -1177
rect 7072 -2165 7118 -2153
rect -7062 -2203 -6870 -2197
rect -7062 -2237 -7050 -2203
rect -6882 -2237 -6870 -2203
rect -7062 -2243 -6870 -2237
rect -6804 -2203 -6612 -2197
rect -6804 -2237 -6792 -2203
rect -6624 -2237 -6612 -2203
rect -6804 -2243 -6612 -2237
rect -6546 -2203 -6354 -2197
rect -6546 -2237 -6534 -2203
rect -6366 -2237 -6354 -2203
rect -6546 -2243 -6354 -2237
rect -6288 -2203 -6096 -2197
rect -6288 -2237 -6276 -2203
rect -6108 -2237 -6096 -2203
rect -6288 -2243 -6096 -2237
rect -6030 -2203 -5838 -2197
rect -6030 -2237 -6018 -2203
rect -5850 -2237 -5838 -2203
rect -6030 -2243 -5838 -2237
rect -5772 -2203 -5580 -2197
rect -5772 -2237 -5760 -2203
rect -5592 -2237 -5580 -2203
rect -5772 -2243 -5580 -2237
rect -5514 -2203 -5322 -2197
rect -5514 -2237 -5502 -2203
rect -5334 -2237 -5322 -2203
rect -5514 -2243 -5322 -2237
rect -5256 -2203 -5064 -2197
rect -5256 -2237 -5244 -2203
rect -5076 -2237 -5064 -2203
rect -5256 -2243 -5064 -2237
rect -4998 -2203 -4806 -2197
rect -4998 -2237 -4986 -2203
rect -4818 -2237 -4806 -2203
rect -4998 -2243 -4806 -2237
rect -4740 -2203 -4548 -2197
rect -4740 -2237 -4728 -2203
rect -4560 -2237 -4548 -2203
rect -4740 -2243 -4548 -2237
rect -4482 -2203 -4290 -2197
rect -4482 -2237 -4470 -2203
rect -4302 -2237 -4290 -2203
rect -4482 -2243 -4290 -2237
rect -4224 -2203 -4032 -2197
rect -4224 -2237 -4212 -2203
rect -4044 -2237 -4032 -2203
rect -4224 -2243 -4032 -2237
rect -3966 -2203 -3774 -2197
rect -3966 -2237 -3954 -2203
rect -3786 -2237 -3774 -2203
rect -3966 -2243 -3774 -2237
rect -3708 -2203 -3516 -2197
rect -3708 -2237 -3696 -2203
rect -3528 -2237 -3516 -2203
rect -3708 -2243 -3516 -2237
rect -3450 -2203 -3258 -2197
rect -3450 -2237 -3438 -2203
rect -3270 -2237 -3258 -2203
rect -3450 -2243 -3258 -2237
rect -3192 -2203 -3000 -2197
rect -3192 -2237 -3180 -2203
rect -3012 -2237 -3000 -2203
rect -3192 -2243 -3000 -2237
rect -2934 -2203 -2742 -2197
rect -2934 -2237 -2922 -2203
rect -2754 -2237 -2742 -2203
rect -2934 -2243 -2742 -2237
rect -2676 -2203 -2484 -2197
rect -2676 -2237 -2664 -2203
rect -2496 -2237 -2484 -2203
rect -2676 -2243 -2484 -2237
rect -2418 -2203 -2226 -2197
rect -2418 -2237 -2406 -2203
rect -2238 -2237 -2226 -2203
rect -2418 -2243 -2226 -2237
rect -2160 -2203 -1968 -2197
rect -2160 -2237 -2148 -2203
rect -1980 -2237 -1968 -2203
rect -2160 -2243 -1968 -2237
rect -1902 -2203 -1710 -2197
rect -1902 -2237 -1890 -2203
rect -1722 -2237 -1710 -2203
rect -1902 -2243 -1710 -2237
rect -1644 -2203 -1452 -2197
rect -1644 -2237 -1632 -2203
rect -1464 -2237 -1452 -2203
rect -1644 -2243 -1452 -2237
rect -1386 -2203 -1194 -2197
rect -1386 -2237 -1374 -2203
rect -1206 -2237 -1194 -2203
rect -1386 -2243 -1194 -2237
rect -1128 -2203 -936 -2197
rect -1128 -2237 -1116 -2203
rect -948 -2237 -936 -2203
rect -1128 -2243 -936 -2237
rect -870 -2203 -678 -2197
rect -870 -2237 -858 -2203
rect -690 -2237 -678 -2203
rect -870 -2243 -678 -2237
rect -612 -2203 -420 -2197
rect -612 -2237 -600 -2203
rect -432 -2237 -420 -2203
rect -612 -2243 -420 -2237
rect -354 -2203 -162 -2197
rect -354 -2237 -342 -2203
rect -174 -2237 -162 -2203
rect -354 -2243 -162 -2237
rect -96 -2203 96 -2197
rect -96 -2237 -84 -2203
rect 84 -2237 96 -2203
rect -96 -2243 96 -2237
rect 162 -2203 354 -2197
rect 162 -2237 174 -2203
rect 342 -2237 354 -2203
rect 162 -2243 354 -2237
rect 420 -2203 612 -2197
rect 420 -2237 432 -2203
rect 600 -2237 612 -2203
rect 420 -2243 612 -2237
rect 678 -2203 870 -2197
rect 678 -2237 690 -2203
rect 858 -2237 870 -2203
rect 678 -2243 870 -2237
rect 936 -2203 1128 -2197
rect 936 -2237 948 -2203
rect 1116 -2237 1128 -2203
rect 936 -2243 1128 -2237
rect 1194 -2203 1386 -2197
rect 1194 -2237 1206 -2203
rect 1374 -2237 1386 -2203
rect 1194 -2243 1386 -2237
rect 1452 -2203 1644 -2197
rect 1452 -2237 1464 -2203
rect 1632 -2237 1644 -2203
rect 1452 -2243 1644 -2237
rect 1710 -2203 1902 -2197
rect 1710 -2237 1722 -2203
rect 1890 -2237 1902 -2203
rect 1710 -2243 1902 -2237
rect 1968 -2203 2160 -2197
rect 1968 -2237 1980 -2203
rect 2148 -2237 2160 -2203
rect 1968 -2243 2160 -2237
rect 2226 -2203 2418 -2197
rect 2226 -2237 2238 -2203
rect 2406 -2237 2418 -2203
rect 2226 -2243 2418 -2237
rect 2484 -2203 2676 -2197
rect 2484 -2237 2496 -2203
rect 2664 -2237 2676 -2203
rect 2484 -2243 2676 -2237
rect 2742 -2203 2934 -2197
rect 2742 -2237 2754 -2203
rect 2922 -2237 2934 -2203
rect 2742 -2243 2934 -2237
rect 3000 -2203 3192 -2197
rect 3000 -2237 3012 -2203
rect 3180 -2237 3192 -2203
rect 3000 -2243 3192 -2237
rect 3258 -2203 3450 -2197
rect 3258 -2237 3270 -2203
rect 3438 -2237 3450 -2203
rect 3258 -2243 3450 -2237
rect 3516 -2203 3708 -2197
rect 3516 -2237 3528 -2203
rect 3696 -2237 3708 -2203
rect 3516 -2243 3708 -2237
rect 3774 -2203 3966 -2197
rect 3774 -2237 3786 -2203
rect 3954 -2237 3966 -2203
rect 3774 -2243 3966 -2237
rect 4032 -2203 4224 -2197
rect 4032 -2237 4044 -2203
rect 4212 -2237 4224 -2203
rect 4032 -2243 4224 -2237
rect 4290 -2203 4482 -2197
rect 4290 -2237 4302 -2203
rect 4470 -2237 4482 -2203
rect 4290 -2243 4482 -2237
rect 4548 -2203 4740 -2197
rect 4548 -2237 4560 -2203
rect 4728 -2237 4740 -2203
rect 4548 -2243 4740 -2237
rect 4806 -2203 4998 -2197
rect 4806 -2237 4818 -2203
rect 4986 -2237 4998 -2203
rect 4806 -2243 4998 -2237
rect 5064 -2203 5256 -2197
rect 5064 -2237 5076 -2203
rect 5244 -2237 5256 -2203
rect 5064 -2243 5256 -2237
rect 5322 -2203 5514 -2197
rect 5322 -2237 5334 -2203
rect 5502 -2237 5514 -2203
rect 5322 -2243 5514 -2237
rect 5580 -2203 5772 -2197
rect 5580 -2237 5592 -2203
rect 5760 -2237 5772 -2203
rect 5580 -2243 5772 -2237
rect 5838 -2203 6030 -2197
rect 5838 -2237 5850 -2203
rect 6018 -2237 6030 -2203
rect 5838 -2243 6030 -2237
rect 6096 -2203 6288 -2197
rect 6096 -2237 6108 -2203
rect 6276 -2237 6288 -2203
rect 6096 -2243 6288 -2237
rect 6354 -2203 6546 -2197
rect 6354 -2237 6366 -2203
rect 6534 -2237 6546 -2203
rect 6354 -2243 6546 -2237
rect 6612 -2203 6804 -2197
rect 6612 -2237 6624 -2203
rect 6792 -2237 6804 -2203
rect 6612 -2243 6804 -2237
rect 6870 -2203 7062 -2197
rect 6870 -2237 6882 -2203
rect 7050 -2237 7062 -2203
rect 6870 -2243 7062 -2237
<< properties >>
string FIXED_BBOX -7229 -2358 7229 2358
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 1.0 m 4 nf 55 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
