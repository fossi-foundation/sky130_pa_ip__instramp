magic
tech sky130A
timestamp 1729620069
<< pwell >>
rect -1487 -379 1487 379
<< mvnmos >>
rect -1373 -250 -1273 250
rect -1184 -250 -1084 250
rect -995 -250 -895 250
rect -806 -250 -706 250
rect -617 -250 -517 250
rect -428 -250 -328 250
rect -239 -250 -139 250
rect -50 -250 50 250
rect 139 -250 239 250
rect 328 -250 428 250
rect 517 -250 617 250
rect 706 -250 806 250
rect 895 -250 995 250
rect 1084 -250 1184 250
rect 1273 -250 1373 250
<< mvndiff >>
rect -1402 244 -1373 250
rect -1402 -244 -1396 244
rect -1379 -244 -1373 244
rect -1402 -250 -1373 -244
rect -1273 244 -1244 250
rect -1273 -244 -1267 244
rect -1250 -244 -1244 244
rect -1273 -250 -1244 -244
rect -1213 244 -1184 250
rect -1213 -244 -1207 244
rect -1190 -244 -1184 244
rect -1213 -250 -1184 -244
rect -1084 244 -1055 250
rect -1084 -244 -1078 244
rect -1061 -244 -1055 244
rect -1084 -250 -1055 -244
rect -1024 244 -995 250
rect -1024 -244 -1018 244
rect -1001 -244 -995 244
rect -1024 -250 -995 -244
rect -895 244 -866 250
rect -895 -244 -889 244
rect -872 -244 -866 244
rect -895 -250 -866 -244
rect -835 244 -806 250
rect -835 -244 -829 244
rect -812 -244 -806 244
rect -835 -250 -806 -244
rect -706 244 -677 250
rect -706 -244 -700 244
rect -683 -244 -677 244
rect -706 -250 -677 -244
rect -646 244 -617 250
rect -646 -244 -640 244
rect -623 -244 -617 244
rect -646 -250 -617 -244
rect -517 244 -488 250
rect -517 -244 -511 244
rect -494 -244 -488 244
rect -517 -250 -488 -244
rect -457 244 -428 250
rect -457 -244 -451 244
rect -434 -244 -428 244
rect -457 -250 -428 -244
rect -328 244 -299 250
rect -328 -244 -322 244
rect -305 -244 -299 244
rect -328 -250 -299 -244
rect -268 244 -239 250
rect -268 -244 -262 244
rect -245 -244 -239 244
rect -268 -250 -239 -244
rect -139 244 -110 250
rect -139 -244 -133 244
rect -116 -244 -110 244
rect -139 -250 -110 -244
rect -79 244 -50 250
rect -79 -244 -73 244
rect -56 -244 -50 244
rect -79 -250 -50 -244
rect 50 244 79 250
rect 50 -244 56 244
rect 73 -244 79 244
rect 50 -250 79 -244
rect 110 244 139 250
rect 110 -244 116 244
rect 133 -244 139 244
rect 110 -250 139 -244
rect 239 244 268 250
rect 239 -244 245 244
rect 262 -244 268 244
rect 239 -250 268 -244
rect 299 244 328 250
rect 299 -244 305 244
rect 322 -244 328 244
rect 299 -250 328 -244
rect 428 244 457 250
rect 428 -244 434 244
rect 451 -244 457 244
rect 428 -250 457 -244
rect 488 244 517 250
rect 488 -244 494 244
rect 511 -244 517 244
rect 488 -250 517 -244
rect 617 244 646 250
rect 617 -244 623 244
rect 640 -244 646 244
rect 617 -250 646 -244
rect 677 244 706 250
rect 677 -244 683 244
rect 700 -244 706 244
rect 677 -250 706 -244
rect 806 244 835 250
rect 806 -244 812 244
rect 829 -244 835 244
rect 806 -250 835 -244
rect 866 244 895 250
rect 866 -244 872 244
rect 889 -244 895 244
rect 866 -250 895 -244
rect 995 244 1024 250
rect 995 -244 1001 244
rect 1018 -244 1024 244
rect 995 -250 1024 -244
rect 1055 244 1084 250
rect 1055 -244 1061 244
rect 1078 -244 1084 244
rect 1055 -250 1084 -244
rect 1184 244 1213 250
rect 1184 -244 1190 244
rect 1207 -244 1213 244
rect 1184 -250 1213 -244
rect 1244 244 1273 250
rect 1244 -244 1250 244
rect 1267 -244 1273 244
rect 1244 -250 1273 -244
rect 1373 244 1402 250
rect 1373 -244 1379 244
rect 1396 -244 1402 244
rect 1373 -250 1402 -244
<< mvndiffc >>
rect -1396 -244 -1379 244
rect -1267 -244 -1250 244
rect -1207 -244 -1190 244
rect -1078 -244 -1061 244
rect -1018 -244 -1001 244
rect -889 -244 -872 244
rect -829 -244 -812 244
rect -700 -244 -683 244
rect -640 -244 -623 244
rect -511 -244 -494 244
rect -451 -244 -434 244
rect -322 -244 -305 244
rect -262 -244 -245 244
rect -133 -244 -116 244
rect -73 -244 -56 244
rect 56 -244 73 244
rect 116 -244 133 244
rect 245 -244 262 244
rect 305 -244 322 244
rect 434 -244 451 244
rect 494 -244 511 244
rect 623 -244 640 244
rect 683 -244 700 244
rect 812 -244 829 244
rect 872 -244 889 244
rect 1001 -244 1018 244
rect 1061 -244 1078 244
rect 1190 -244 1207 244
rect 1250 -244 1267 244
rect 1379 -244 1396 244
<< mvpsubdiff >>
rect -1469 355 1469 361
rect -1469 338 -1415 355
rect 1415 338 1469 355
rect -1469 332 1469 338
rect -1469 307 -1440 332
rect -1469 -307 -1463 307
rect -1446 -307 -1440 307
rect 1440 307 1469 332
rect -1469 -332 -1440 -307
rect 1440 -307 1446 307
rect 1463 -307 1469 307
rect 1440 -332 1469 -307
rect -1469 -338 1469 -332
rect -1469 -355 -1415 -338
rect 1415 -355 1469 -338
rect -1469 -361 1469 -355
<< mvpsubdiffcont >>
rect -1415 338 1415 355
rect -1463 -307 -1446 307
rect 1446 -307 1463 307
rect -1415 -355 1415 -338
<< poly >>
rect -1373 286 -1273 294
rect -1373 269 -1365 286
rect -1281 269 -1273 286
rect -1373 250 -1273 269
rect -1184 286 -1084 294
rect -1184 269 -1176 286
rect -1092 269 -1084 286
rect -1184 250 -1084 269
rect -995 286 -895 294
rect -995 269 -987 286
rect -903 269 -895 286
rect -995 250 -895 269
rect -806 286 -706 294
rect -806 269 -798 286
rect -714 269 -706 286
rect -806 250 -706 269
rect -617 286 -517 294
rect -617 269 -609 286
rect -525 269 -517 286
rect -617 250 -517 269
rect -428 286 -328 294
rect -428 269 -420 286
rect -336 269 -328 286
rect -428 250 -328 269
rect -239 286 -139 294
rect -239 269 -231 286
rect -147 269 -139 286
rect -239 250 -139 269
rect -50 286 50 294
rect -50 269 -42 286
rect 42 269 50 286
rect -50 250 50 269
rect 139 286 239 294
rect 139 269 147 286
rect 231 269 239 286
rect 139 250 239 269
rect 328 286 428 294
rect 328 269 336 286
rect 420 269 428 286
rect 328 250 428 269
rect 517 286 617 294
rect 517 269 525 286
rect 609 269 617 286
rect 517 250 617 269
rect 706 286 806 294
rect 706 269 714 286
rect 798 269 806 286
rect 706 250 806 269
rect 895 286 995 294
rect 895 269 903 286
rect 987 269 995 286
rect 895 250 995 269
rect 1084 286 1184 294
rect 1084 269 1092 286
rect 1176 269 1184 286
rect 1084 250 1184 269
rect 1273 286 1373 294
rect 1273 269 1281 286
rect 1365 269 1373 286
rect 1273 250 1373 269
rect -1373 -269 -1273 -250
rect -1373 -286 -1365 -269
rect -1281 -286 -1273 -269
rect -1373 -294 -1273 -286
rect -1184 -269 -1084 -250
rect -1184 -286 -1176 -269
rect -1092 -286 -1084 -269
rect -1184 -294 -1084 -286
rect -995 -269 -895 -250
rect -995 -286 -987 -269
rect -903 -286 -895 -269
rect -995 -294 -895 -286
rect -806 -269 -706 -250
rect -806 -286 -798 -269
rect -714 -286 -706 -269
rect -806 -294 -706 -286
rect -617 -269 -517 -250
rect -617 -286 -609 -269
rect -525 -286 -517 -269
rect -617 -294 -517 -286
rect -428 -269 -328 -250
rect -428 -286 -420 -269
rect -336 -286 -328 -269
rect -428 -294 -328 -286
rect -239 -269 -139 -250
rect -239 -286 -231 -269
rect -147 -286 -139 -269
rect -239 -294 -139 -286
rect -50 -269 50 -250
rect -50 -286 -42 -269
rect 42 -286 50 -269
rect -50 -294 50 -286
rect 139 -269 239 -250
rect 139 -286 147 -269
rect 231 -286 239 -269
rect 139 -294 239 -286
rect 328 -269 428 -250
rect 328 -286 336 -269
rect 420 -286 428 -269
rect 328 -294 428 -286
rect 517 -269 617 -250
rect 517 -286 525 -269
rect 609 -286 617 -269
rect 517 -294 617 -286
rect 706 -269 806 -250
rect 706 -286 714 -269
rect 798 -286 806 -269
rect 706 -294 806 -286
rect 895 -269 995 -250
rect 895 -286 903 -269
rect 987 -286 995 -269
rect 895 -294 995 -286
rect 1084 -269 1184 -250
rect 1084 -286 1092 -269
rect 1176 -286 1184 -269
rect 1084 -294 1184 -286
rect 1273 -269 1373 -250
rect 1273 -286 1281 -269
rect 1365 -286 1373 -269
rect 1273 -294 1373 -286
<< polycont >>
rect -1365 269 -1281 286
rect -1176 269 -1092 286
rect -987 269 -903 286
rect -798 269 -714 286
rect -609 269 -525 286
rect -420 269 -336 286
rect -231 269 -147 286
rect -42 269 42 286
rect 147 269 231 286
rect 336 269 420 286
rect 525 269 609 286
rect 714 269 798 286
rect 903 269 987 286
rect 1092 269 1176 286
rect 1281 269 1365 286
rect -1365 -286 -1281 -269
rect -1176 -286 -1092 -269
rect -987 -286 -903 -269
rect -798 -286 -714 -269
rect -609 -286 -525 -269
rect -420 -286 -336 -269
rect -231 -286 -147 -269
rect -42 -286 42 -269
rect 147 -286 231 -269
rect 336 -286 420 -269
rect 525 -286 609 -269
rect 714 -286 798 -269
rect 903 -286 987 -269
rect 1092 -286 1176 -269
rect 1281 -286 1365 -269
<< locali >>
rect -1463 338 -1415 355
rect 1415 338 1463 355
rect -1463 307 -1446 338
rect 1446 307 1463 338
rect -1373 269 -1365 286
rect -1281 269 -1273 286
rect -1184 269 -1176 286
rect -1092 269 -1084 286
rect -995 269 -987 286
rect -903 269 -895 286
rect -806 269 -798 286
rect -714 269 -706 286
rect -617 269 -609 286
rect -525 269 -517 286
rect -428 269 -420 286
rect -336 269 -328 286
rect -239 269 -231 286
rect -147 269 -139 286
rect -50 269 -42 286
rect 42 269 50 286
rect 139 269 147 286
rect 231 269 239 286
rect 328 269 336 286
rect 420 269 428 286
rect 517 269 525 286
rect 609 269 617 286
rect 706 269 714 286
rect 798 269 806 286
rect 895 269 903 286
rect 987 269 995 286
rect 1084 269 1092 286
rect 1176 269 1184 286
rect 1273 269 1281 286
rect 1365 269 1373 286
rect -1396 244 -1379 252
rect -1396 -252 -1379 -244
rect -1267 244 -1250 252
rect -1267 -252 -1250 -244
rect -1207 244 -1190 252
rect -1207 -252 -1190 -244
rect -1078 244 -1061 252
rect -1078 -252 -1061 -244
rect -1018 244 -1001 252
rect -1018 -252 -1001 -244
rect -889 244 -872 252
rect -889 -252 -872 -244
rect -829 244 -812 252
rect -829 -252 -812 -244
rect -700 244 -683 252
rect -700 -252 -683 -244
rect -640 244 -623 252
rect -640 -252 -623 -244
rect -511 244 -494 252
rect -511 -252 -494 -244
rect -451 244 -434 252
rect -451 -252 -434 -244
rect -322 244 -305 252
rect -322 -252 -305 -244
rect -262 244 -245 252
rect -262 -252 -245 -244
rect -133 244 -116 252
rect -133 -252 -116 -244
rect -73 244 -56 252
rect -73 -252 -56 -244
rect 56 244 73 252
rect 56 -252 73 -244
rect 116 244 133 252
rect 116 -252 133 -244
rect 245 244 262 252
rect 245 -252 262 -244
rect 305 244 322 252
rect 305 -252 322 -244
rect 434 244 451 252
rect 434 -252 451 -244
rect 494 244 511 252
rect 494 -252 511 -244
rect 623 244 640 252
rect 623 -252 640 -244
rect 683 244 700 252
rect 683 -252 700 -244
rect 812 244 829 252
rect 812 -252 829 -244
rect 872 244 889 252
rect 872 -252 889 -244
rect 1001 244 1018 252
rect 1001 -252 1018 -244
rect 1061 244 1078 252
rect 1061 -252 1078 -244
rect 1190 244 1207 252
rect 1190 -252 1207 -244
rect 1250 244 1267 252
rect 1250 -252 1267 -244
rect 1379 244 1396 252
rect 1379 -252 1396 -244
rect -1373 -286 -1365 -269
rect -1281 -286 -1273 -269
rect -1184 -286 -1176 -269
rect -1092 -286 -1084 -269
rect -995 -286 -987 -269
rect -903 -286 -895 -269
rect -806 -286 -798 -269
rect -714 -286 -706 -269
rect -617 -286 -609 -269
rect -525 -286 -517 -269
rect -428 -286 -420 -269
rect -336 -286 -328 -269
rect -239 -286 -231 -269
rect -147 -286 -139 -269
rect -50 -286 -42 -269
rect 42 -286 50 -269
rect 139 -286 147 -269
rect 231 -286 239 -269
rect 328 -286 336 -269
rect 420 -286 428 -269
rect 517 -286 525 -269
rect 609 -286 617 -269
rect 706 -286 714 -269
rect 798 -286 806 -269
rect 895 -286 903 -269
rect 987 -286 995 -269
rect 1084 -286 1092 -269
rect 1176 -286 1184 -269
rect 1273 -286 1281 -269
rect 1365 -286 1373 -269
rect -1463 -338 -1446 -307
rect 1446 -338 1463 -307
rect -1463 -355 -1415 -338
rect 1415 -355 1463 -338
<< viali >>
rect -1365 269 -1281 286
rect -1176 269 -1092 286
rect -987 269 -903 286
rect -798 269 -714 286
rect -609 269 -525 286
rect -420 269 -336 286
rect -231 269 -147 286
rect -42 269 42 286
rect 147 269 231 286
rect 336 269 420 286
rect 525 269 609 286
rect 714 269 798 286
rect 903 269 987 286
rect 1092 269 1176 286
rect 1281 269 1365 286
rect -1396 -244 -1379 244
rect -1267 -244 -1250 244
rect -1207 -244 -1190 244
rect -1078 -244 -1061 244
rect -1018 -244 -1001 244
rect -889 -244 -872 244
rect -829 -244 -812 244
rect -700 -244 -683 244
rect -640 -244 -623 244
rect -511 -244 -494 244
rect -451 -244 -434 244
rect -322 -244 -305 244
rect -262 -244 -245 244
rect -133 -244 -116 244
rect -73 -244 -56 244
rect 56 -244 73 244
rect 116 -244 133 244
rect 245 -244 262 244
rect 305 -244 322 244
rect 434 -244 451 244
rect 494 -244 511 244
rect 623 -244 640 244
rect 683 -244 700 244
rect 812 -244 829 244
rect 872 -244 889 244
rect 1001 -244 1018 244
rect 1061 -244 1078 244
rect 1190 -244 1207 244
rect 1250 -244 1267 244
rect 1379 -244 1396 244
rect -1365 -286 -1281 -269
rect -1176 -286 -1092 -269
rect -987 -286 -903 -269
rect -798 -286 -714 -269
rect -609 -286 -525 -269
rect -420 -286 -336 -269
rect -231 -286 -147 -269
rect -42 -286 42 -269
rect 147 -286 231 -269
rect 336 -286 420 -269
rect 525 -286 609 -269
rect 714 -286 798 -269
rect 903 -286 987 -269
rect 1092 -286 1176 -269
rect 1281 -286 1365 -269
<< metal1 >>
rect -1371 286 -1275 289
rect -1371 269 -1365 286
rect -1281 269 -1275 286
rect -1371 266 -1275 269
rect -1182 286 -1086 289
rect -1182 269 -1176 286
rect -1092 269 -1086 286
rect -1182 266 -1086 269
rect -993 286 -897 289
rect -993 269 -987 286
rect -903 269 -897 286
rect -993 266 -897 269
rect -804 286 -708 289
rect -804 269 -798 286
rect -714 269 -708 286
rect -804 266 -708 269
rect -615 286 -519 289
rect -615 269 -609 286
rect -525 269 -519 286
rect -615 266 -519 269
rect -426 286 -330 289
rect -426 269 -420 286
rect -336 269 -330 286
rect -426 266 -330 269
rect -237 286 -141 289
rect -237 269 -231 286
rect -147 269 -141 286
rect -237 266 -141 269
rect -48 286 48 289
rect -48 269 -42 286
rect 42 269 48 286
rect -48 266 48 269
rect 141 286 237 289
rect 141 269 147 286
rect 231 269 237 286
rect 141 266 237 269
rect 330 286 426 289
rect 330 269 336 286
rect 420 269 426 286
rect 330 266 426 269
rect 519 286 615 289
rect 519 269 525 286
rect 609 269 615 286
rect 519 266 615 269
rect 708 286 804 289
rect 708 269 714 286
rect 798 269 804 286
rect 708 266 804 269
rect 897 286 993 289
rect 897 269 903 286
rect 987 269 993 286
rect 897 266 993 269
rect 1086 286 1182 289
rect 1086 269 1092 286
rect 1176 269 1182 286
rect 1086 266 1182 269
rect 1275 286 1371 289
rect 1275 269 1281 286
rect 1365 269 1371 286
rect 1275 266 1371 269
rect -1399 244 -1376 250
rect -1399 -244 -1396 244
rect -1379 -244 -1376 244
rect -1399 -250 -1376 -244
rect -1270 244 -1247 250
rect -1270 -244 -1267 244
rect -1250 -244 -1247 244
rect -1270 -250 -1247 -244
rect -1210 244 -1187 250
rect -1210 -244 -1207 244
rect -1190 -244 -1187 244
rect -1210 -250 -1187 -244
rect -1081 244 -1058 250
rect -1081 -244 -1078 244
rect -1061 -244 -1058 244
rect -1081 -250 -1058 -244
rect -1021 244 -998 250
rect -1021 -244 -1018 244
rect -1001 -244 -998 244
rect -1021 -250 -998 -244
rect -892 244 -869 250
rect -892 -244 -889 244
rect -872 -244 -869 244
rect -892 -250 -869 -244
rect -832 244 -809 250
rect -832 -244 -829 244
rect -812 -244 -809 244
rect -832 -250 -809 -244
rect -703 244 -680 250
rect -703 -244 -700 244
rect -683 -244 -680 244
rect -703 -250 -680 -244
rect -643 244 -620 250
rect -643 -244 -640 244
rect -623 -244 -620 244
rect -643 -250 -620 -244
rect -514 244 -491 250
rect -514 -244 -511 244
rect -494 -244 -491 244
rect -514 -250 -491 -244
rect -454 244 -431 250
rect -454 -244 -451 244
rect -434 -244 -431 244
rect -454 -250 -431 -244
rect -325 244 -302 250
rect -325 -244 -322 244
rect -305 -244 -302 244
rect -325 -250 -302 -244
rect -265 244 -242 250
rect -265 -244 -262 244
rect -245 -244 -242 244
rect -265 -250 -242 -244
rect -136 244 -113 250
rect -136 -244 -133 244
rect -116 -244 -113 244
rect -136 -250 -113 -244
rect -76 244 -53 250
rect -76 -244 -73 244
rect -56 -244 -53 244
rect -76 -250 -53 -244
rect 53 244 76 250
rect 53 -244 56 244
rect 73 -244 76 244
rect 53 -250 76 -244
rect 113 244 136 250
rect 113 -244 116 244
rect 133 -244 136 244
rect 113 -250 136 -244
rect 242 244 265 250
rect 242 -244 245 244
rect 262 -244 265 244
rect 242 -250 265 -244
rect 302 244 325 250
rect 302 -244 305 244
rect 322 -244 325 244
rect 302 -250 325 -244
rect 431 244 454 250
rect 431 -244 434 244
rect 451 -244 454 244
rect 431 -250 454 -244
rect 491 244 514 250
rect 491 -244 494 244
rect 511 -244 514 244
rect 491 -250 514 -244
rect 620 244 643 250
rect 620 -244 623 244
rect 640 -244 643 244
rect 620 -250 643 -244
rect 680 244 703 250
rect 680 -244 683 244
rect 700 -244 703 244
rect 680 -250 703 -244
rect 809 244 832 250
rect 809 -244 812 244
rect 829 -244 832 244
rect 809 -250 832 -244
rect 869 244 892 250
rect 869 -244 872 244
rect 889 -244 892 244
rect 869 -250 892 -244
rect 998 244 1021 250
rect 998 -244 1001 244
rect 1018 -244 1021 244
rect 998 -250 1021 -244
rect 1058 244 1081 250
rect 1058 -244 1061 244
rect 1078 -244 1081 244
rect 1058 -250 1081 -244
rect 1187 244 1210 250
rect 1187 -244 1190 244
rect 1207 -244 1210 244
rect 1187 -250 1210 -244
rect 1247 244 1270 250
rect 1247 -244 1250 244
rect 1267 -244 1270 244
rect 1247 -250 1270 -244
rect 1376 244 1399 250
rect 1376 -244 1379 244
rect 1396 -244 1399 244
rect 1376 -250 1399 -244
rect -1371 -269 -1275 -266
rect -1371 -286 -1365 -269
rect -1281 -286 -1275 -269
rect -1371 -289 -1275 -286
rect -1182 -269 -1086 -266
rect -1182 -286 -1176 -269
rect -1092 -286 -1086 -269
rect -1182 -289 -1086 -286
rect -993 -269 -897 -266
rect -993 -286 -987 -269
rect -903 -286 -897 -269
rect -993 -289 -897 -286
rect -804 -269 -708 -266
rect -804 -286 -798 -269
rect -714 -286 -708 -269
rect -804 -289 -708 -286
rect -615 -269 -519 -266
rect -615 -286 -609 -269
rect -525 -286 -519 -269
rect -615 -289 -519 -286
rect -426 -269 -330 -266
rect -426 -286 -420 -269
rect -336 -286 -330 -269
rect -426 -289 -330 -286
rect -237 -269 -141 -266
rect -237 -286 -231 -269
rect -147 -286 -141 -269
rect -237 -289 -141 -286
rect -48 -269 48 -266
rect -48 -286 -42 -269
rect 42 -286 48 -269
rect -48 -289 48 -286
rect 141 -269 237 -266
rect 141 -286 147 -269
rect 231 -286 237 -269
rect 141 -289 237 -286
rect 330 -269 426 -266
rect 330 -286 336 -269
rect 420 -286 426 -269
rect 330 -289 426 -286
rect 519 -269 615 -266
rect 519 -286 525 -269
rect 609 -286 615 -269
rect 519 -289 615 -286
rect 708 -269 804 -266
rect 708 -286 714 -269
rect 798 -286 804 -269
rect 708 -289 804 -286
rect 897 -269 993 -266
rect 897 -286 903 -269
rect 987 -286 993 -269
rect 897 -289 993 -286
rect 1086 -269 1182 -266
rect 1086 -286 1092 -269
rect 1176 -286 1182 -269
rect 1086 -289 1182 -286
rect 1275 -269 1371 -266
rect 1275 -286 1281 -269
rect 1365 -286 1371 -269
rect 1275 -289 1371 -286
<< properties >>
string FIXED_BBOX -1454 -346 1454 346
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 1.0 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
