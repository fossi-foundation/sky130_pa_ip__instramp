magic
tech sky130A
magscale 1 2
timestamp 1731187918
<< error_s >>
rect 27004 22792 27006 23146
rect 27004 21886 27006 22446
rect 480 -9354 486 -9348
rect 534 -9354 540 -9348
rect 474 -9360 480 -9354
rect 540 -9360 546 -9354
rect 29224 -9360 29230 -9354
rect 29272 -9360 29278 -9354
rect 29218 -9366 29224 -9360
rect 29278 -9366 29284 -9360
rect 474 -10500 480 -10494
rect 540 -10500 546 -10494
rect 29218 -10498 29224 -10492
rect 29278 -10498 29284 -10492
rect 480 -10506 486 -10500
rect 534 -10506 540 -10500
rect 29224 -10504 29230 -10498
rect 29272 -10504 29278 -10498
<< dnwell >>
rect 364 22792 27006 25984
rect 364 21886 27004 22792
rect 364 21846 27006 21886
rect 364 11850 14926 21846
rect 364 6612 15240 11850
rect 364 -7116 14942 6612
rect 364 -11292 29434 -7116
<< locali >>
rect 9813 21480 11041 21499
rect 9813 18386 9826 21480
rect 9874 21429 11041 21480
rect 9874 18424 9883 21429
rect 10971 20744 11041 21429
rect 10971 18424 10980 20744
rect 9874 18418 10980 18424
rect 9874 18386 9936 18418
rect 9813 18360 9936 18386
rect 10926 18378 10980 18418
rect 11032 18424 11041 20744
rect 11314 21425 12525 21495
rect 11314 20758 11384 21425
rect 11032 18378 11042 18424
rect 11314 18423 11324 20758
rect 10926 18360 11042 18378
rect 9813 18354 11042 18360
rect 11313 18392 11324 18423
rect 11376 18423 11384 20758
rect 12455 20600 12525 21425
rect 12455 18423 12470 20600
rect 11376 18422 12470 18423
rect 11376 18392 11428 18422
rect 11313 18364 11428 18392
rect 12418 18378 12470 18422
rect 12520 18378 12525 20600
rect 12418 18364 12525 18378
rect 11313 18353 12525 18364
rect 12782 21442 14009 21491
rect 12782 21421 13954 21442
rect 12782 21342 12852 21421
rect 12782 18378 12786 21342
rect 12842 18417 12852 21342
rect 13939 18417 13954 21421
rect 12842 18412 13954 18417
rect 12842 18378 12904 18412
rect 12782 18354 12904 18378
rect 13894 18390 13954 18412
rect 14006 18390 14009 21442
rect 13894 18354 14009 18390
rect 12782 18350 14009 18354
rect 12785 18347 14009 18350
rect 9696 11800 15209 11817
rect 9696 11796 9802 11800
rect 9696 6706 9708 11796
rect 9746 11764 9802 11796
rect 15110 11796 15209 11800
rect 15110 11764 15154 11796
rect 9746 11751 15154 11764
rect 9746 6746 9762 11751
rect 15143 6746 15154 11751
rect 9746 6730 15154 6746
rect 9746 6706 10038 6730
rect 9696 6694 10038 6706
rect 14892 6700 15154 6730
rect 15198 6700 15209 11796
rect 14892 6694 15209 6700
rect 9696 6681 15209 6694
rect 9696 6680 15208 6681
rect 466 -7158 29290 -7142
rect 466 -7206 594 -7158
rect 14694 -7198 14944 -7158
rect 29200 -7198 29290 -7158
rect 14694 -7206 29290 -7198
rect 466 -7218 29290 -7206
rect 466 -7340 542 -7218
rect 29214 -7278 29290 -7218
rect 466 -11166 494 -7340
rect 466 -11218 542 -11166
rect 29214 -11182 29238 -7278
rect 29274 -11182 29290 -7278
rect 29214 -11218 29290 -11182
rect 466 -11228 29290 -11218
rect 466 -11276 594 -11228
rect 29198 -11276 29290 -11228
rect 466 -11294 29290 -11276
<< viali >>
rect 9826 18386 9874 21480
rect 9936 18360 10926 18418
rect 10980 18378 11032 20744
rect 11324 18392 11376 20758
rect 11428 18364 12418 18422
rect 12470 18378 12520 20600
rect 12786 18378 12842 21342
rect 12904 18354 13894 18412
rect 13954 18390 14006 21442
rect 9708 6706 9746 11796
rect 9802 11764 15110 11800
rect 10038 6694 14892 6730
rect 15154 6700 15198 11796
rect 594 -7206 14694 -7158
rect 14944 -7198 29200 -7158
rect 494 -11166 548 -7340
rect 29238 -11182 29274 -7278
rect 594 -11276 29198 -11228
<< metal1 >>
rect 26808 28030 27008 28230
rect 26786 27603 26986 27746
rect 2867 27546 26986 27603
rect 573 27506 2854 27518
rect 573 27283 590 27506
rect 1060 27283 2854 27506
rect 573 27268 2854 27283
rect 368 26054 384 26198
rect 598 26187 2890 26198
rect 598 26065 2551 26187
rect 2797 26065 2890 26187
rect 598 26054 2890 26065
rect 13328 22280 13532 22300
rect 3000 22116 3074 22206
rect 2886 22102 3322 22116
rect 2886 22010 2902 22102
rect 3306 22010 3322 22102
rect 3385 22096 3459 22196
rect 5440 22096 5514 22196
rect 3385 22022 5514 22096
rect 5785 22096 5859 22196
rect 7840 22096 7914 22196
rect 5785 22022 7914 22096
rect 8185 22096 8259 22196
rect 10240 22096 10314 22196
rect 8185 22022 10314 22096
rect 10585 22096 10659 22196
rect 12640 22096 12714 22196
rect 10585 22022 12714 22096
rect 2886 21996 3322 22010
rect 2816 21760 3016 21960
rect 12985 21950 13059 22196
rect 13328 22124 13350 22280
rect 13510 22124 13532 22280
rect 13328 22104 13532 22124
rect 14300 22288 14436 22300
rect 14300 22116 14312 22288
rect 14420 22116 14436 22288
rect 14928 22189 14929 22218
rect 14928 22156 15128 22189
rect 9694 21916 9892 21940
rect 9694 21664 9716 21916
rect 9872 21664 9892 21916
rect 9694 21640 9892 21664
rect 9814 21504 9892 21640
rect 9812 21480 9892 21504
rect 9812 18430 9826 21480
rect 9338 18386 9826 18430
rect 9874 18434 9892 21480
rect 9974 21873 13059 21950
rect 9974 20898 10050 21873
rect 13342 21867 13418 22104
rect 14234 21912 14436 22116
rect 15385 22096 15459 22196
rect 17440 22096 17514 22196
rect 15385 22022 17514 22096
rect 17785 22096 17859 22196
rect 19840 22096 19914 22196
rect 17785 22022 19914 22096
rect 20185 22096 20259 22196
rect 22240 22096 22314 22196
rect 20185 22022 22314 22096
rect 22585 22096 22659 22223
rect 24640 22096 24714 22204
rect 22585 22022 24714 22096
rect 24958 22114 25158 22196
rect 24958 22104 25260 22114
rect 24958 22012 24968 22104
rect 25246 22012 25260 22104
rect 24958 22004 25260 22012
rect 14214 21867 14234 21912
rect 13342 21832 14234 21867
rect 10476 21788 14234 21832
rect 14434 21788 15066 21912
rect 10476 21756 13418 21788
rect 10146 20906 10382 21338
rect 10476 20902 10552 21756
rect 12978 21710 13182 21720
rect 12978 21604 12992 21710
rect 13172 21604 13182 21710
rect 12978 21594 13182 21604
rect 10642 21552 11024 21562
rect 10642 21466 10654 21552
rect 11010 21466 11024 21552
rect 10642 21456 11024 21466
rect 10642 20906 10718 21456
rect 12290 21444 13010 21514
rect 11002 21392 11332 21408
rect 11002 21338 11018 21392
rect 10810 21278 11018 21338
rect 11314 21338 11332 21392
rect 11314 21278 11530 21338
rect 10810 20904 11530 21278
rect 11626 20906 11862 21338
rect 11958 20906 12196 21338
rect 12124 20812 12196 20906
rect 12290 20904 12360 21444
rect 12764 21342 12864 21382
rect 10970 20744 11050 20786
rect 9982 18508 10220 18940
rect 10314 18508 10552 18940
rect 10646 18508 10884 18940
rect 10970 18434 10980 20744
rect 9874 18418 10980 18434
rect 9874 18386 9936 18418
rect 9338 18360 9936 18386
rect 10926 18378 10980 18418
rect 11032 18430 11050 20744
rect 11306 20758 11386 20792
rect 11306 18430 11324 20758
rect 11032 18392 11324 18430
rect 11376 18432 11386 20758
rect 12124 20704 12684 20812
rect 12450 20600 12534 20634
rect 11458 18506 11696 18938
rect 11790 18506 12028 18938
rect 12122 18506 12360 18938
rect 12450 18432 12470 20600
rect 11376 18422 12470 18432
rect 11376 18392 11428 18422
rect 11032 18378 11428 18392
rect 10926 18364 11428 18378
rect 12418 18378 12470 18422
rect 12520 18432 12534 20600
rect 12520 18378 12536 18432
rect 12418 18364 12536 18378
rect 10926 18360 12536 18364
rect 9338 18340 12536 18360
rect 12628 18284 12684 20704
rect 12764 18378 12786 21342
rect 12842 18432 12864 21342
rect 12940 20906 13010 21444
rect 13106 20906 13176 21594
rect 13270 20906 13348 21756
rect 13770 21610 14728 21728
rect 14908 21610 14933 21728
rect 13438 20902 13676 21340
rect 13770 20906 13844 21610
rect 14278 21530 14620 21546
rect 13932 21442 14034 21498
rect 12940 18506 13178 18938
rect 13272 18506 13510 18938
rect 13604 18506 13842 18938
rect 13932 18432 13954 21442
rect 12842 18412 13954 18432
rect 12842 18378 12904 18412
rect 12764 18354 12904 18378
rect 13894 18390 13954 18412
rect 14006 18390 14034 21442
rect 14278 21440 14298 21530
rect 14604 21440 14620 21530
rect 14278 21430 14620 21440
rect 13894 18354 14034 18390
rect 12764 18338 14034 18354
rect 12628 18228 13720 18284
rect 13664 15206 13720 18228
rect 13934 17780 14034 18338
rect 13934 17604 14034 17614
rect 14506 15290 14600 21430
rect 14980 21075 15066 21788
rect 14819 20989 15066 21075
rect 14820 15738 14906 20989
rect 14820 15643 14946 15738
rect 14505 15216 14826 15290
rect 10452 15150 13720 15206
rect 2950 12199 3016 12639
rect 7040 12496 7240 12568
rect 7040 12402 7240 12410
rect 14752 12020 14826 15216
rect 14870 12310 14946 15643
rect 14870 12302 15368 12310
rect 14870 12204 14878 12302
rect 15354 12204 15368 12302
rect 14870 12194 15368 12204
rect 15528 12302 15888 12312
rect 15528 12200 15540 12302
rect 15876 12200 15888 12302
rect 15528 12192 15888 12200
rect 14752 11943 15332 12020
rect 9694 11800 15210 11818
rect 9694 11796 9802 11800
rect 9694 6706 9708 11796
rect 9746 11764 9802 11796
rect 15110 11796 15210 11800
rect 15110 11764 15154 11796
rect 9746 11750 15154 11764
rect 9746 6706 9762 11750
rect 9836 11224 10072 11656
rect 10168 11224 10404 11656
rect 10500 11224 10736 11656
rect 10832 11224 11068 11656
rect 11164 11224 11400 11656
rect 11496 11224 11732 11656
rect 11828 11224 12064 11656
rect 12160 11224 12396 11656
rect 12492 11224 12728 11656
rect 12824 11224 13060 11656
rect 13156 11224 13392 11656
rect 13488 11224 13724 11656
rect 13820 11224 14056 11656
rect 14152 11224 14388 11656
rect 14484 11224 14720 11656
rect 14816 11224 15052 11656
rect 9694 6680 9762 6706
rect 9830 6656 9912 7260
rect 10002 6824 10238 7256
rect 10334 6824 10570 7256
rect 10666 6824 10902 7256
rect 10998 6824 11234 7256
rect 11330 6824 11566 7256
rect 11662 6824 11898 7256
rect 11994 6824 12230 7256
rect 12326 6824 12562 7256
rect 12658 6824 12894 7256
rect 12990 6824 13226 7256
rect 13322 6824 13558 7256
rect 13654 6824 13890 7256
rect 13986 6824 14222 7256
rect 14318 6824 14554 7256
rect 14650 6824 14886 7256
rect 10012 6730 14912 6748
rect 10012 6694 10038 6730
rect 14892 6694 14912 6730
rect 10012 6680 14912 6694
rect 9820 6646 9948 6656
rect 9820 6310 9832 6646
rect 9938 6310 9948 6646
rect 14980 6439 15052 7256
rect 15142 6700 15154 11750
rect 15198 6700 15210 11796
rect 15142 6682 15210 6700
rect 15254 6439 15332 11943
rect 14561 6361 15332 6439
rect 9820 6298 9948 6310
rect 14562 5486 14618 6361
rect 15542 6091 15634 12192
rect 10382 5430 14618 5486
rect 14976 6021 15634 6091
rect 2948 2437 3014 3119
rect 7038 2762 7238 2848
rect 7038 2684 7238 2694
rect 14976 2598 15042 6021
rect 14880 2590 15192 2598
rect 14880 2522 14894 2590
rect 15184 2522 15192 2590
rect 14880 2514 15192 2522
rect 7036 -6976 7236 -6900
rect 2536 -7000 2802 -6990
rect 2536 -7152 2550 -7000
rect 466 -7158 2550 -7152
rect 2792 -7152 2802 -7000
rect 7036 -7042 7046 -6976
rect 7328 -7042 7338 -6976
rect 7600 -7070 7800 -6862
rect 14978 -6886 15042 2514
rect 11578 -6950 15042 -6886
rect 7926 -7042 7942 -6976
rect 8264 -6978 8280 -6976
rect 11578 -6978 11642 -6950
rect 8264 -7042 11642 -6978
rect 13850 -7006 14468 -6994
rect 13850 -7042 13868 -7006
rect 11688 -7070 13868 -7042
rect 7600 -7110 13868 -7070
rect 14454 -7026 14468 -7006
rect 14454 -7110 14856 -7026
rect 7600 -7124 11768 -7110
rect 2792 -7158 14710 -7152
rect 466 -7206 594 -7158
rect 14694 -7206 14710 -7158
rect 466 -7208 2550 -7206
rect 2792 -7208 14710 -7206
rect 466 -7218 14710 -7208
rect 466 -7340 566 -7218
rect 466 -9354 494 -7340
rect 466 -10500 480 -9354
rect 466 -11166 494 -10500
rect 548 -11166 566 -7340
rect 662 -7346 732 -7298
rect 14772 -7302 14856 -7110
rect 14916 -7158 29290 -7142
rect 14916 -7198 14944 -7158
rect 29200 -7198 29290 -7158
rect 14916 -7218 29290 -7198
rect 29214 -7278 29290 -7218
rect 662 -7734 732 -7720
rect 828 -7734 1064 -7302
rect 1160 -7734 1396 -7302
rect 1492 -7734 1728 -7302
rect 1824 -7734 2060 -7302
rect 2156 -7734 2392 -7302
rect 2488 -7734 2724 -7302
rect 2820 -7734 3056 -7302
rect 3152 -7734 3388 -7302
rect 3484 -7734 3720 -7302
rect 3816 -7734 4052 -7302
rect 4148 -7734 4384 -7302
rect 4480 -7734 4716 -7302
rect 4812 -7734 5048 -7302
rect 5144 -7734 5380 -7302
rect 5476 -7734 5712 -7302
rect 5808 -7734 6044 -7302
rect 6140 -7734 6376 -7302
rect 6472 -7734 6708 -7302
rect 6804 -7734 7040 -7302
rect 7136 -7734 7372 -7302
rect 7468 -7734 7704 -7302
rect 7800 -7734 8036 -7302
rect 8132 -7734 8368 -7302
rect 8464 -7734 8700 -7302
rect 8796 -7734 9032 -7302
rect 9128 -7734 9364 -7302
rect 9460 -7734 9696 -7302
rect 9792 -7734 10028 -7302
rect 10124 -7734 10360 -7302
rect 10456 -7734 10692 -7302
rect 10788 -7734 11024 -7302
rect 11120 -7734 11356 -7302
rect 11452 -7734 11688 -7302
rect 11784 -7734 12020 -7302
rect 12116 -7734 12352 -7302
rect 12448 -7734 12684 -7302
rect 12780 -7734 13016 -7302
rect 13112 -7734 13348 -7302
rect 13444 -7734 13680 -7302
rect 13776 -7734 14012 -7302
rect 14108 -7734 14344 -7302
rect 14440 -7734 14676 -7302
rect 14772 -7734 15008 -7302
rect 15104 -7734 15340 -7302
rect 15436 -7734 15672 -7302
rect 15768 -7734 16004 -7302
rect 16100 -7734 16336 -7302
rect 16432 -7734 16668 -7302
rect 16764 -7734 17000 -7302
rect 17096 -7734 17332 -7302
rect 17428 -7734 17664 -7302
rect 17760 -7734 17996 -7302
rect 18092 -7734 18328 -7302
rect 18424 -7734 18660 -7302
rect 18756 -7734 18992 -7302
rect 19088 -7734 19324 -7302
rect 19420 -7734 19656 -7302
rect 19752 -7734 19988 -7302
rect 20084 -7734 20320 -7302
rect 20416 -7734 20652 -7302
rect 20748 -7734 20984 -7302
rect 21080 -7734 21316 -7302
rect 21412 -7734 21648 -7302
rect 21744 -7734 21980 -7302
rect 22076 -7734 22312 -7302
rect 22408 -7734 22644 -7302
rect 22740 -7734 22976 -7302
rect 23072 -7734 23308 -7302
rect 23404 -7734 23640 -7302
rect 23736 -7734 23972 -7302
rect 24068 -7734 24304 -7302
rect 24400 -7734 24636 -7302
rect 24732 -7734 24968 -7302
rect 25064 -7734 25300 -7302
rect 25396 -7734 25632 -7302
rect 25728 -7734 25964 -7302
rect 26060 -7734 26296 -7302
rect 26392 -7734 26628 -7302
rect 26724 -7734 26960 -7302
rect 27056 -7734 27292 -7302
rect 27388 -7734 27624 -7302
rect 27720 -7734 27956 -7302
rect 28052 -7734 28288 -7302
rect 28384 -7734 28620 -7302
rect 28716 -7734 28952 -7302
rect 29048 -7350 29118 -7302
rect 29048 -7734 29118 -7720
rect 29214 -9360 29238 -7278
rect 29274 -9360 29290 -7278
rect 29214 -10498 29224 -9360
rect 29278 -10498 29290 -9360
rect 662 -11110 898 -10678
rect 994 -11110 1230 -10678
rect 1326 -11110 1562 -10678
rect 1658 -11110 1894 -10678
rect 1990 -11110 2226 -10678
rect 2322 -11110 2558 -10678
rect 2654 -11110 2890 -10678
rect 2986 -11110 3222 -10678
rect 3318 -11110 3554 -10678
rect 3650 -11110 3886 -10678
rect 3982 -11110 4218 -10678
rect 4314 -11110 4550 -10678
rect 4646 -11110 4882 -10678
rect 4978 -11110 5214 -10678
rect 5310 -11110 5546 -10678
rect 5642 -11110 5878 -10678
rect 5974 -11110 6210 -10678
rect 6306 -11110 6542 -10678
rect 6638 -11110 6874 -10678
rect 6970 -11110 7206 -10678
rect 7302 -11110 7538 -10678
rect 7634 -11110 7870 -10678
rect 7966 -11110 8202 -10678
rect 8298 -11110 8534 -10678
rect 8630 -11110 8866 -10678
rect 8962 -11110 9198 -10678
rect 9294 -11110 9530 -10678
rect 9626 -11110 9862 -10678
rect 9958 -11110 10194 -10678
rect 10290 -11110 10526 -10678
rect 10622 -11110 10858 -10678
rect 10954 -11110 11190 -10678
rect 11286 -11110 11522 -10678
rect 11618 -11110 11854 -10678
rect 11950 -11110 12186 -10678
rect 12282 -11110 12518 -10678
rect 12614 -11110 12850 -10678
rect 12946 -11110 13182 -10678
rect 13278 -11110 13514 -10678
rect 13610 -11110 13846 -10678
rect 13942 -11110 14178 -10678
rect 14274 -11110 14510 -10678
rect 14606 -11110 14842 -10678
rect 14938 -11110 15174 -10678
rect 15270 -11110 15506 -10678
rect 15602 -11110 15838 -10678
rect 15934 -11110 16170 -10678
rect 16266 -11110 16502 -10678
rect 16598 -11110 16834 -10678
rect 16930 -11110 17166 -10678
rect 17262 -11110 17498 -10678
rect 17594 -11110 17830 -10678
rect 17926 -11110 18162 -10678
rect 18258 -11110 18494 -10678
rect 18590 -11110 18826 -10678
rect 18922 -11110 19158 -10678
rect 19254 -11110 19490 -10678
rect 19586 -11110 19822 -10678
rect 19918 -11110 20154 -10678
rect 20250 -11110 20486 -10678
rect 20582 -11110 20818 -10678
rect 20914 -11110 21150 -10678
rect 21246 -11110 21482 -10678
rect 21578 -11110 21814 -10678
rect 21910 -11110 22146 -10678
rect 22242 -11110 22478 -10678
rect 22574 -11110 22810 -10678
rect 22906 -11110 23142 -10678
rect 23238 -11110 23474 -10678
rect 23570 -11110 23806 -10678
rect 23902 -11110 24138 -10678
rect 24234 -11110 24470 -10678
rect 24566 -11110 24802 -10678
rect 24898 -11110 25134 -10678
rect 25230 -11110 25466 -10678
rect 25562 -11110 25798 -10678
rect 25894 -11110 26130 -10678
rect 26226 -11110 26462 -10678
rect 26558 -11110 26794 -10678
rect 26890 -11110 27126 -10678
rect 27222 -11110 27458 -10678
rect 27554 -11110 27790 -10678
rect 27886 -11110 28122 -10678
rect 28218 -11110 28454 -10678
rect 28550 -11110 28786 -10678
rect 28882 -11110 29118 -10678
rect 466 -11206 566 -11166
rect 29214 -11182 29238 -10498
rect 29274 -11182 29290 -10498
rect 29214 -11206 29290 -11182
rect 466 -11228 29290 -11206
rect 466 -11276 594 -11228
rect 29198 -11276 29290 -11228
rect 466 -11294 29290 -11276
<< via1 >>
rect 590 27283 1060 27506
rect 384 26054 598 26198
rect 2551 26065 2797 26187
rect 2902 22010 3306 22102
rect 13350 22124 13510 22280
rect 14312 22116 14420 22288
rect 14929 22189 15128 22388
rect 9716 21664 9872 21916
rect 24968 22012 25246 22104
rect 14234 21788 14434 21912
rect 12992 21604 13172 21710
rect 10654 21466 11010 21552
rect 11018 21278 11314 21392
rect 14728 21610 14908 21728
rect 14298 21440 14604 21530
rect 13934 17614 14034 17780
rect 7040 12410 7240 12496
rect 14878 12204 15354 12302
rect 15540 12200 15876 12302
rect 9832 6310 9938 6646
rect 7038 2694 7238 2762
rect 14894 2522 15184 2590
rect 2550 -7158 2792 -7000
rect 7046 -7042 7328 -6976
rect 7942 -7042 8264 -6976
rect 13868 -7110 14454 -7006
rect 2550 -7206 2792 -7158
rect 2550 -7208 2792 -7206
rect 480 -10500 494 -9354
rect 494 -10500 540 -9354
rect 662 -7720 732 -7346
rect 29048 -7720 29118 -7350
rect 29224 -10498 29238 -9360
rect 29238 -10498 29274 -9360
rect 29274 -10498 29278 -9360
<< metal2 >>
rect 3188 28058 3388 28258
rect 5588 28058 5788 28258
rect 7988 28058 8188 28258
rect 10388 28058 10588 28258
rect 12788 28058 12988 28258
rect 15188 28058 15388 28258
rect 17588 28058 17788 28258
rect 19988 28058 20188 28258
rect 22388 28058 22588 28258
rect 24788 28058 24988 28258
rect 576 27506 1074 27520
rect 576 27283 590 27506
rect 1060 27283 1074 27506
rect 576 27267 1074 27283
rect 384 26198 598 26216
rect 2538 26187 2810 26200
rect 2538 26065 2551 26187
rect 2797 26065 2810 26187
rect 2538 26055 2810 26065
rect 384 21234 598 26054
rect 4878 22546 5082 22568
rect 4878 22390 4900 22546
rect 5062 22390 5082 22546
rect 4878 22372 5082 22390
rect 7278 22546 7482 22568
rect 7278 22390 7300 22546
rect 7462 22390 7482 22546
rect 7278 22372 7482 22390
rect 9678 22546 9882 22568
rect 9678 22390 9700 22546
rect 9862 22390 9882 22546
rect 9678 22372 9882 22390
rect 12078 22546 12282 22568
rect 12078 22390 12100 22546
rect 12262 22390 12282 22546
rect 12078 22372 12282 22390
rect 14478 22546 14682 22568
rect 14478 22390 14500 22546
rect 14662 22390 14682 22546
rect 14478 22372 14682 22390
rect 16878 22546 17082 22568
rect 16878 22390 16900 22546
rect 17062 22390 17082 22546
rect 14764 22388 15142 22389
rect 4632 22280 4836 22300
rect 4632 22124 4654 22280
rect 4814 22124 4836 22280
rect 2888 22102 3322 22116
rect 4632 22104 4836 22124
rect 7032 22280 7236 22300
rect 7032 22124 7054 22280
rect 7214 22124 7236 22280
rect 7032 22104 7236 22124
rect 9432 22280 9636 22300
rect 9432 22124 9454 22280
rect 9614 22124 9636 22280
rect 9432 22104 9636 22124
rect 11832 22280 12036 22300
rect 11832 22124 11854 22280
rect 12014 22124 12036 22280
rect 11832 22104 12036 22124
rect 13328 22280 13532 22300
rect 13328 22124 13350 22280
rect 13510 22124 13532 22280
rect 13328 22104 13532 22124
rect 14232 22288 14436 22300
rect 14232 22280 14312 22288
rect 14232 22124 14254 22280
rect 14232 22116 14312 22124
rect 14420 22116 14436 22288
rect 14764 22223 14929 22388
rect 14232 22104 14436 22116
rect 14763 22189 14929 22223
rect 15128 22189 15142 22388
rect 16878 22372 17082 22390
rect 19278 22546 19482 22568
rect 19278 22390 19300 22546
rect 19462 22390 19482 22546
rect 19278 22372 19482 22390
rect 21678 22546 21882 22568
rect 21678 22390 21700 22546
rect 21862 22390 21882 22546
rect 21678 22372 21882 22390
rect 24078 22546 24282 22568
rect 24078 22390 24100 22546
rect 24262 22390 24282 22546
rect 24078 22372 24282 22390
rect 26478 22546 26682 22568
rect 26478 22390 26500 22546
rect 26662 22390 26682 22546
rect 26478 22372 26682 22390
rect 16632 22280 16836 22300
rect 2888 22010 2902 22102
rect 3306 22010 3322 22102
rect 2888 21996 3322 22010
rect 9308 21916 12870 21940
rect 9308 21664 9716 21916
rect 9872 21664 12870 21916
rect 14234 21912 14434 22104
rect 14763 22013 14891 22189
rect 16632 22122 16654 22280
rect 16814 22178 16836 22280
rect 19032 22280 19236 22300
rect 16814 22122 16834 22178
rect 16632 22104 16834 22122
rect 19032 22124 19054 22280
rect 19214 22124 19236 22280
rect 19032 22104 19236 22124
rect 21432 22280 21636 22300
rect 21432 22124 21454 22280
rect 21614 22124 21636 22280
rect 21432 22104 21636 22124
rect 23832 22280 24036 22300
rect 23832 22124 23854 22280
rect 24014 22124 24036 22280
rect 23832 22104 24036 22124
rect 26232 22280 26436 22300
rect 26232 22124 26254 22280
rect 26414 22124 26436 22280
rect 24958 22104 25260 22114
rect 26232 22104 26436 22124
rect 24958 22072 24968 22104
rect 14234 21774 14434 21788
rect 14529 22005 14891 22013
rect 14529 21836 14671 22005
rect 14859 21836 14891 22005
rect 14529 21824 14891 21836
rect 15026 22012 24968 22072
rect 25246 22012 25260 22104
rect 15026 21996 25260 22012
rect 14529 21727 14645 21824
rect 15026 21728 15115 21996
rect 14712 21727 14728 21728
rect 9308 21638 12870 21664
rect 12978 21710 14645 21727
rect 12978 21604 12992 21710
rect 13172 21611 14645 21710
rect 13172 21604 13182 21611
rect 14711 21610 14728 21727
rect 14908 21610 15115 21728
rect 14711 21609 15115 21610
rect 12978 21594 13182 21604
rect 14728 21598 14908 21609
rect 15026 21608 15115 21609
rect 10642 21552 11024 21562
rect 10642 21466 10654 21552
rect 11010 21542 11024 21552
rect 14278 21542 14620 21546
rect 11010 21530 14620 21542
rect 11010 21466 14298 21530
rect 10642 21456 14298 21466
rect 14278 21440 14298 21456
rect 14604 21440 14620 21530
rect 14278 21430 14620 21440
rect 11002 21392 11332 21408
rect 11002 21278 11018 21392
rect 11314 21346 11332 21392
rect 14894 21346 15094 21466
rect 11314 21278 15094 21346
rect 11002 21266 15094 21278
rect 14978 21058 15094 21266
rect 9320 17614 13934 17780
rect 14034 17614 14049 17780
rect 7027 12410 7040 12496
rect 7240 12410 14684 12496
rect 364 12370 490 12380
rect 364 12270 376 12370
rect 480 12354 490 12370
rect 480 12346 14392 12354
rect 480 12274 14194 12346
rect 480 12270 490 12274
rect 364 12256 490 12270
rect 14178 12154 14194 12274
rect 14382 12154 14392 12346
rect 14590 12300 14684 12410
rect 14870 12304 15368 12310
rect 15528 12304 15888 12312
rect 14870 12302 15888 12304
rect 14870 12300 14878 12302
rect 14590 12212 14878 12300
rect 14870 12204 14878 12212
rect 15354 12204 15540 12302
rect 14870 12194 15368 12204
rect 15528 12200 15540 12204
rect 15876 12200 15888 12302
rect 15528 12192 15888 12200
rect 14178 12142 14392 12154
rect 14646 12130 14870 12138
rect 9306 11748 14474 12062
rect 14646 11884 14656 12130
rect 14858 11884 14870 12130
rect 14646 11876 14870 11884
rect 7018 2694 7038 2762
rect 7238 2694 14498 2762
rect 14430 2598 14498 2694
rect 14430 2590 15192 2598
rect 14430 2530 14894 2590
rect 14880 2522 14894 2530
rect 15184 2522 15192 2590
rect 14880 2514 15192 2522
rect 2536 -7000 2802 -6990
rect 2536 -7244 2550 -7000
rect 2792 -7244 2802 -7000
rect 7036 -7042 7046 -6976
rect 7328 -7042 7942 -6976
rect 8264 -7042 8280 -6976
rect 13850 -7006 14474 -6994
rect 13850 -7110 13868 -7006
rect 14454 -7110 14474 -7006
rect 13850 -7124 14474 -7110
rect 14644 -7128 14662 -7016
rect 14860 -7042 14870 -7016
rect 14860 -7128 15206 -7042
rect 2536 -7254 2802 -7244
rect 15094 -7278 15206 -7128
rect 384 -7342 736 -7334
rect 384 -7756 394 -7342
rect 468 -7346 736 -7342
rect 468 -7720 662 -7346
rect 732 -7720 736 -7346
rect 15094 -7350 29138 -7278
rect 15094 -7390 29048 -7350
rect 468 -7756 736 -7720
rect 384 -7770 736 -7756
rect 29036 -7720 29048 -7390
rect 29118 -7720 29138 -7350
rect 29036 -7770 29138 -7720
<< via2 >>
rect 590 27283 1060 27506
rect 2551 26065 2797 26187
rect 4900 22390 5062 22546
rect 7300 22390 7462 22546
rect 9700 22390 9862 22546
rect 12100 22390 12262 22546
rect 14500 22390 14662 22546
rect 16900 22390 17062 22546
rect 4654 22124 4814 22280
rect 7054 22124 7214 22280
rect 9454 22124 9614 22280
rect 11854 22124 12014 22280
rect 13350 22124 13510 22280
rect 14254 22124 14312 22280
rect 14312 22124 14414 22280
rect 19300 22390 19462 22546
rect 21700 22390 21862 22546
rect 24100 22390 24262 22546
rect 26500 22390 26662 22546
rect 2902 22010 3306 22102
rect 16654 22122 16814 22280
rect 19054 22124 19214 22280
rect 21454 22124 21614 22280
rect 23854 22124 24014 22280
rect 26254 22124 26414 22280
rect 14671 21836 14859 22005
rect 376 12270 480 12370
rect 14194 12154 14382 12346
rect 14656 11884 14858 12130
rect 2550 -7208 2792 -7000
rect 2550 -7244 2792 -7208
rect 13868 -7110 14454 -7006
rect 14662 -7128 14860 -7016
rect 394 -7756 468 -7342
<< metal3 >>
rect 576 27506 1076 28242
rect 576 27283 590 27506
rect 1060 27283 1076 27506
rect 576 21933 1076 27283
rect 2538 26187 2808 28242
rect 2538 26065 2551 26187
rect 2797 26065 2808 26187
rect 2538 21939 2808 26065
rect 4878 22546 5082 22568
rect 4878 22508 4900 22546
rect 2934 22396 4900 22508
rect 4878 22390 4900 22396
rect 5062 22508 5082 22546
rect 7278 22546 7482 22568
rect 7278 22508 7300 22546
rect 5062 22396 7300 22508
rect 5062 22390 5082 22396
rect 4878 22372 5082 22390
rect 7278 22390 7300 22396
rect 7462 22508 7482 22546
rect 9678 22546 9882 22568
rect 9678 22508 9700 22546
rect 7462 22396 9700 22508
rect 7462 22390 7482 22396
rect 7278 22372 7482 22390
rect 9678 22390 9700 22396
rect 9862 22508 9882 22546
rect 12078 22546 12282 22568
rect 12078 22508 12100 22546
rect 9862 22396 12100 22508
rect 9862 22390 9882 22396
rect 9678 22372 9882 22390
rect 12078 22390 12100 22396
rect 12262 22508 12282 22546
rect 14478 22546 14682 22568
rect 14478 22508 14500 22546
rect 12262 22396 14500 22508
rect 12262 22390 12282 22396
rect 12078 22372 12282 22390
rect 14478 22390 14500 22396
rect 14662 22508 14682 22546
rect 15002 22554 15572 22574
rect 15002 22508 15030 22554
rect 14662 22412 15030 22508
rect 15548 22508 15572 22554
rect 16878 22546 17082 22568
rect 16878 22508 16900 22546
rect 15548 22412 16900 22508
rect 14662 22396 16900 22412
rect 14662 22390 14682 22396
rect 14478 22372 14682 22390
rect 16878 22390 16900 22396
rect 17062 22508 17082 22546
rect 19278 22546 19482 22568
rect 19278 22508 19300 22546
rect 17062 22396 19300 22508
rect 17062 22390 17082 22396
rect 16878 22372 17082 22390
rect 19278 22390 19300 22396
rect 19462 22508 19482 22546
rect 21678 22546 21882 22568
rect 21678 22508 21700 22546
rect 19462 22396 21700 22508
rect 19462 22390 19482 22396
rect 19278 22372 19482 22390
rect 21678 22390 21700 22396
rect 21862 22508 21882 22546
rect 24078 22546 24282 22568
rect 24078 22508 24100 22546
rect 21862 22396 24100 22508
rect 21862 22390 21882 22396
rect 21678 22372 21882 22390
rect 24078 22390 24100 22396
rect 24262 22508 24282 22546
rect 26478 22546 26682 22568
rect 26478 22508 26500 22546
rect 24262 22396 26500 22508
rect 24262 22390 24282 22396
rect 24078 22372 24282 22390
rect 26478 22390 26500 22396
rect 26662 22508 26682 22546
rect 26662 22396 26824 22508
rect 26662 22390 26682 22396
rect 26478 22372 26682 22390
rect 4632 22290 4836 22300
rect 7032 22290 7236 22300
rect 9432 22290 9636 22300
rect 11832 22290 12036 22300
rect 13328 22290 13532 22300
rect 14232 22290 14436 22300
rect 16632 22290 16836 22300
rect 19032 22290 19236 22300
rect 21432 22290 21636 22300
rect 23832 22290 24036 22300
rect 26232 22290 26436 22300
rect 2934 22280 26934 22290
rect 2934 22178 4654 22280
rect 4632 22124 4654 22178
rect 4814 22178 7054 22280
rect 4814 22124 4836 22178
rect 2886 22102 3322 22116
rect 4632 22104 4836 22124
rect 7032 22124 7054 22178
rect 7214 22178 9454 22280
rect 7214 22124 7236 22178
rect 7032 22104 7236 22124
rect 9432 22124 9454 22178
rect 9614 22178 11854 22280
rect 9614 22124 9636 22178
rect 9432 22104 9636 22124
rect 11832 22124 11854 22178
rect 12014 22178 13350 22280
rect 12014 22124 12036 22178
rect 11832 22104 12036 22124
rect 13328 22124 13350 22178
rect 13510 22178 14254 22280
rect 13510 22124 13532 22178
rect 13328 22104 13532 22124
rect 14232 22124 14254 22178
rect 14414 22178 16654 22280
rect 14414 22124 14436 22178
rect 14232 22104 14436 22124
rect 16632 22122 16654 22178
rect 16814 22178 19054 22280
rect 16814 22122 16836 22178
rect 16632 22104 16836 22122
rect 19032 22124 19054 22178
rect 19214 22178 21454 22280
rect 19214 22124 19236 22178
rect 19032 22104 19236 22124
rect 21432 22124 21454 22178
rect 21614 22178 23854 22280
rect 21614 22124 21636 22178
rect 21432 22104 21636 22124
rect 23832 22124 23854 22178
rect 24014 22178 26254 22280
rect 24014 22124 24036 22178
rect 23832 22104 24036 22124
rect 26232 22124 26254 22178
rect 26414 22178 26934 22280
rect 26414 22124 26436 22178
rect 26232 22104 26436 22124
rect 2886 22010 2902 22102
rect 3306 22010 3322 22102
rect 26734 22090 26934 22178
rect 2886 21996 3322 22010
rect 14658 22005 14869 22038
rect 726 21686 926 21886
rect 14658 21836 14671 22005
rect 14859 21889 14869 22005
rect 14859 21836 14870 21889
rect 14658 21092 14870 21836
rect 2578 20814 2778 21014
rect 364 12370 490 12380
rect 364 12270 376 12370
rect 480 12270 490 12370
rect 364 12256 490 12270
rect 386 -7342 474 12256
rect 574 12216 1074 12564
rect 2538 12222 2808 13782
rect 14658 12490 14870 14044
rect 14180 12346 14870 12490
rect 14180 12154 14194 12346
rect 14382 12278 14870 12346
rect 14382 12154 14392 12278
rect 14180 12142 14392 12154
rect 14646 12130 14870 12138
rect 14646 11884 14656 12130
rect 14858 11884 14870 12130
rect 14646 11876 14870 11884
rect 14656 11378 14868 11876
rect 572 2454 1072 2850
rect 2536 2472 2806 4058
rect 386 -7756 394 -7342
rect 468 -7756 474 -7342
rect 386 -7770 474 -7756
rect 572 -11250 1072 -6892
rect 2534 -7000 2804 -5680
rect 2534 -7244 2550 -7000
rect 2792 -7244 2804 -7000
rect 13850 -7006 14474 -6994
rect 13850 -7110 13868 -7006
rect 14454 -7110 14474 -7006
rect 13850 -7124 14474 -7110
rect 14654 -7016 14866 -5412
rect 2534 -11244 2804 -7244
rect 14654 -7128 14662 -7016
rect 14860 -7128 14866 -7016
rect 14654 -11384 14866 -7128
<< via3 >>
rect 15030 22412 15548 22554
rect 2902 22010 3306 22102
rect 14660 11886 14856 12124
rect 13868 -7110 14454 -7006
<< metal4 >>
rect 15002 22554 15572 22574
rect 15002 22412 15030 22554
rect 15548 22412 15572 22554
rect 15002 22396 15572 22412
rect 2886 22102 3322 22116
rect 2886 22010 2902 22102
rect 3306 22096 3322 22102
rect 3306 22014 14900 22096
rect 3306 22010 3322 22014
rect 2886 21996 3322 22010
rect 14784 12504 14900 22014
rect 14646 12280 14900 12504
rect 14646 12124 14870 12280
rect 14646 11886 14660 12124
rect 14856 11886 14870 12124
rect 14646 11876 14870 11886
rect 15002 -6994 15122 22396
rect 13850 -7006 15122 -6994
rect 13850 -7110 13868 -7006
rect 14454 -7110 15122 -7006
rect 13850 -7124 15122 -7110
<< comment >>
rect 14868 -10456 14928 -7948
use sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP  sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP_0 paramcells
timestamp 1730992408
transform 1 0 13390 0 1 19922
box -616 -1582 616 1582
use sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP  sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP_1
timestamp 1730992408
transform 1 0 10430 0 1 19922
box -616 -1582 616 1582
use sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP  sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP_2
timestamp 1730992408
transform 1 0 11910 0 1 19922
box -616 -1582 616 1582
use sky130_fd_pr__res_xhigh_po_0p35_S4N9LQ  sky130_fd_pr__res_xhigh_po_0p35_S4N9LQ_0 paramcells
timestamp 1730992408
transform 1 0 12444 0 1 9240
box -2774 -2582 2774 2582
use sky130_fd_pr__res_xhigh_po_0p35_V6AMGK  sky130_fd_pr__res_xhigh_po_0p35_V6AMGK_0 paramcells
timestamp 1730992408
transform 1 0 14890 0 1 -9206
box -14394 -2070 14394 2070
use Universal_R_2R_Block2  x1
timestamp 1730992657
transform 0 1 24706 -1 0 29868
box 1610 -2760 7768 -198
use Universal_R_2R_Block2  x2
timestamp 1730992657
transform 0 1 17506 -1 0 29868
box 1610 -2760 7768 -198
use Universal_R_2R_Block2  x3
timestamp 1730992657
transform 0 1 10306 -1 0 29868
box 1610 -2760 7768 -198
use Universal_R_2R_Block2  x4
timestamp 1730992657
transform 0 1 5506 -1 0 29868
box 1610 -2760 7768 -198
use Universal_R_2R_Block2  x5
timestamp 1730992657
transform 0 1 19906 -1 0 29868
box 1610 -2760 7768 -198
use x1_x32_OA  x6
timestamp 1730992408
transform -1 0 15498 0 1 13652
box 628 -1152 15010 8321
use Output_OA  x7
timestamp 1730992408
transform -1 0 15494 0 1 -5816
box 628 -1154 15010 8321
use x1_x32_OA  x8
timestamp 1730992408
transform -1 0 15496 0 1 3932
box 628 -1152 15010 8321
use Universal_R_2R_Block2  x9
timestamp 1730992657
transform 0 1 15106 -1 0 29868
box 1610 -2760 7768 -198
use Universal_R_2R_Block2  x10
timestamp 1730992657
transform 0 1 12706 -1 0 29868
box 1610 -2760 7768 -198
use Universal_R_2R_Block2  x11
timestamp 1730992657
transform 0 1 7906 -1 0 29868
box 1610 -2760 7768 -198
use Universal_R_2R_Block2  x12
timestamp 1730992657
transform 0 1 22306 -1 0 29868
box 1610 -2760 7768 -198
use Universal_R_2R_Block2  x13
timestamp 1730992657
transform 0 1 27106 -1 0 29868
box 1610 -2760 7768 -198
<< labels >>
flabel metal1 2816 21760 3016 21960 0 FreeSans 256 0 0 0 VBIAS
port 17 nsew
flabel metal3 14660 -11380 14860 -11180 0 FreeSans 256 0 0 0 VOUT
port 8 nsew
flabel metal2 14894 21266 15094 21466 0 FreeSans 256 0 0 0 VO1
port 5 nsew
flabel metal3 2578 20814 2778 21014 0 FreeSans 256 0 0 0 AVSS
port 16 nsew
flabel metal3 726 21686 926 21886 0 FreeSans 256 0 0 0 AVDD
port 7 nsew
flabel metal2 24788 28058 24988 28258 0 FreeSans 256 270 0 0 V9
port 3 nsew
flabel metal2 22388 28058 22588 28258 0 FreeSans 256 270 0 0 V8
port 2 nsew
flabel metal2 19988 28058 20188 28258 0 FreeSans 256 270 0 0 V7
port 4 nsew
flabel metal2 17588 28058 17788 28258 0 FreeSans 256 270 0 0 V6
port 0 nsew
flabel metal2 15188 28058 15388 28258 0 FreeSans 256 270 0 0 V5
port 1 nsew
flabel metal2 12788 28058 12988 28258 0 FreeSans 256 270 0 0 V4
port 9 nsew
flabel metal2 10388 28058 10588 28258 0 FreeSans 256 270 0 0 V3
port 10 nsew
flabel metal2 7988 28058 8188 28258 0 FreeSans 256 270 0 0 V2
port 11 nsew
flabel metal2 5588 28058 5788 28258 0 FreeSans 256 270 0 0 V1
port 12 nsew
flabel metal2 3188 28058 3388 28258 0 FreeSans 256 270 0 0 V0
port 13 nsew
flabel metal1 26808 28030 27008 28230 0 FreeSans 256 0 0 0 DVSS
port 15 nsew
flabel metal1 26786 27546 26986 27746 0 FreeSans 256 0 0 0 DVDD
port 6 nsew
flabel metal3 26734 22090 26934 22290 0 FreeSans 256 0 0 0 VCM
port 14 nsew
<< end >>
