magic
tech sky130A
magscale 1 2
timestamp 1729620069
<< pwell >>
rect -235 -640582 235 640582
<< psubdiff >>
rect -199 640512 -103 640546
rect 103 640512 199 640546
rect -199 640450 -165 640512
rect 165 640450 199 640512
rect -199 -640512 -165 -640450
rect 165 -640512 199 -640450
rect -199 -640546 -103 -640512
rect 103 -640546 199 -640512
<< psubdiffcont >>
rect -103 640512 103 640546
rect -199 -640450 -165 640450
rect 165 -640450 199 640450
rect -103 -640546 103 -640512
<< xpolycontact >>
rect -69 639984 69 640416
rect -69 -640416 69 -639984
<< ppolyres >>
rect -69 -639984 69 639984
<< locali >>
rect -199 640512 -103 640546
rect 103 640512 199 640546
rect -199 640450 -165 640512
rect 165 640450 199 640512
rect -199 -640512 -165 -640450
rect 165 -640512 199 -640450
rect -199 -640546 -103 -640512
rect 103 -640546 199 -640512
<< viali >>
rect -53 640001 53 640398
rect -53 -640398 53 -640001
<< metal1 >>
rect -59 640398 59 640410
rect -59 640001 -53 640398
rect 53 640001 59 640398
rect -59 639989 59 640001
rect -59 -640001 59 -639989
rect -59 -640398 -53 -640001
rect 53 -640398 59 -640001
rect -59 -640410 59 -640398
<< properties >>
string FIXED_BBOX -182 -640529 182 640529
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 6400.0 m 1 nx 1 wmin 0.690 lmin 0.50 class resistor rho 319.8 val 2.966meg dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0 mult 1
<< end >>
