magic
tech sky130A
magscale 1 2
timestamp 1729620069
<< pwell >>
rect -3919 -758 3919 758
<< mvnmos >>
rect -3691 -500 -3491 500
rect -3313 -500 -3113 500
rect -2935 -500 -2735 500
rect -2557 -500 -2357 500
rect -2179 -500 -1979 500
rect -1801 -500 -1601 500
rect -1423 -500 -1223 500
rect -1045 -500 -845 500
rect -667 -500 -467 500
rect -289 -500 -89 500
rect 89 -500 289 500
rect 467 -500 667 500
rect 845 -500 1045 500
rect 1223 -500 1423 500
rect 1601 -500 1801 500
rect 1979 -500 2179 500
rect 2357 -500 2557 500
rect 2735 -500 2935 500
rect 3113 -500 3313 500
rect 3491 -500 3691 500
<< mvndiff >>
rect -3749 488 -3691 500
rect -3749 -488 -3737 488
rect -3703 -488 -3691 488
rect -3749 -500 -3691 -488
rect -3491 488 -3433 500
rect -3491 -488 -3479 488
rect -3445 -488 -3433 488
rect -3491 -500 -3433 -488
rect -3371 488 -3313 500
rect -3371 -488 -3359 488
rect -3325 -488 -3313 488
rect -3371 -500 -3313 -488
rect -3113 488 -3055 500
rect -3113 -488 -3101 488
rect -3067 -488 -3055 488
rect -3113 -500 -3055 -488
rect -2993 488 -2935 500
rect -2993 -488 -2981 488
rect -2947 -488 -2935 488
rect -2993 -500 -2935 -488
rect -2735 488 -2677 500
rect -2735 -488 -2723 488
rect -2689 -488 -2677 488
rect -2735 -500 -2677 -488
rect -2615 488 -2557 500
rect -2615 -488 -2603 488
rect -2569 -488 -2557 488
rect -2615 -500 -2557 -488
rect -2357 488 -2299 500
rect -2357 -488 -2345 488
rect -2311 -488 -2299 488
rect -2357 -500 -2299 -488
rect -2237 488 -2179 500
rect -2237 -488 -2225 488
rect -2191 -488 -2179 488
rect -2237 -500 -2179 -488
rect -1979 488 -1921 500
rect -1979 -488 -1967 488
rect -1933 -488 -1921 488
rect -1979 -500 -1921 -488
rect -1859 488 -1801 500
rect -1859 -488 -1847 488
rect -1813 -488 -1801 488
rect -1859 -500 -1801 -488
rect -1601 488 -1543 500
rect -1601 -488 -1589 488
rect -1555 -488 -1543 488
rect -1601 -500 -1543 -488
rect -1481 488 -1423 500
rect -1481 -488 -1469 488
rect -1435 -488 -1423 488
rect -1481 -500 -1423 -488
rect -1223 488 -1165 500
rect -1223 -488 -1211 488
rect -1177 -488 -1165 488
rect -1223 -500 -1165 -488
rect -1103 488 -1045 500
rect -1103 -488 -1091 488
rect -1057 -488 -1045 488
rect -1103 -500 -1045 -488
rect -845 488 -787 500
rect -845 -488 -833 488
rect -799 -488 -787 488
rect -845 -500 -787 -488
rect -725 488 -667 500
rect -725 -488 -713 488
rect -679 -488 -667 488
rect -725 -500 -667 -488
rect -467 488 -409 500
rect -467 -488 -455 488
rect -421 -488 -409 488
rect -467 -500 -409 -488
rect -347 488 -289 500
rect -347 -488 -335 488
rect -301 -488 -289 488
rect -347 -500 -289 -488
rect -89 488 -31 500
rect -89 -488 -77 488
rect -43 -488 -31 488
rect -89 -500 -31 -488
rect 31 488 89 500
rect 31 -488 43 488
rect 77 -488 89 488
rect 31 -500 89 -488
rect 289 488 347 500
rect 289 -488 301 488
rect 335 -488 347 488
rect 289 -500 347 -488
rect 409 488 467 500
rect 409 -488 421 488
rect 455 -488 467 488
rect 409 -500 467 -488
rect 667 488 725 500
rect 667 -488 679 488
rect 713 -488 725 488
rect 667 -500 725 -488
rect 787 488 845 500
rect 787 -488 799 488
rect 833 -488 845 488
rect 787 -500 845 -488
rect 1045 488 1103 500
rect 1045 -488 1057 488
rect 1091 -488 1103 488
rect 1045 -500 1103 -488
rect 1165 488 1223 500
rect 1165 -488 1177 488
rect 1211 -488 1223 488
rect 1165 -500 1223 -488
rect 1423 488 1481 500
rect 1423 -488 1435 488
rect 1469 -488 1481 488
rect 1423 -500 1481 -488
rect 1543 488 1601 500
rect 1543 -488 1555 488
rect 1589 -488 1601 488
rect 1543 -500 1601 -488
rect 1801 488 1859 500
rect 1801 -488 1813 488
rect 1847 -488 1859 488
rect 1801 -500 1859 -488
rect 1921 488 1979 500
rect 1921 -488 1933 488
rect 1967 -488 1979 488
rect 1921 -500 1979 -488
rect 2179 488 2237 500
rect 2179 -488 2191 488
rect 2225 -488 2237 488
rect 2179 -500 2237 -488
rect 2299 488 2357 500
rect 2299 -488 2311 488
rect 2345 -488 2357 488
rect 2299 -500 2357 -488
rect 2557 488 2615 500
rect 2557 -488 2569 488
rect 2603 -488 2615 488
rect 2557 -500 2615 -488
rect 2677 488 2735 500
rect 2677 -488 2689 488
rect 2723 -488 2735 488
rect 2677 -500 2735 -488
rect 2935 488 2993 500
rect 2935 -488 2947 488
rect 2981 -488 2993 488
rect 2935 -500 2993 -488
rect 3055 488 3113 500
rect 3055 -488 3067 488
rect 3101 -488 3113 488
rect 3055 -500 3113 -488
rect 3313 488 3371 500
rect 3313 -488 3325 488
rect 3359 -488 3371 488
rect 3313 -500 3371 -488
rect 3433 488 3491 500
rect 3433 -488 3445 488
rect 3479 -488 3491 488
rect 3433 -500 3491 -488
rect 3691 488 3749 500
rect 3691 -488 3703 488
rect 3737 -488 3749 488
rect 3691 -500 3749 -488
<< mvndiffc >>
rect -3737 -488 -3703 488
rect -3479 -488 -3445 488
rect -3359 -488 -3325 488
rect -3101 -488 -3067 488
rect -2981 -488 -2947 488
rect -2723 -488 -2689 488
rect -2603 -488 -2569 488
rect -2345 -488 -2311 488
rect -2225 -488 -2191 488
rect -1967 -488 -1933 488
rect -1847 -488 -1813 488
rect -1589 -488 -1555 488
rect -1469 -488 -1435 488
rect -1211 -488 -1177 488
rect -1091 -488 -1057 488
rect -833 -488 -799 488
rect -713 -488 -679 488
rect -455 -488 -421 488
rect -335 -488 -301 488
rect -77 -488 -43 488
rect 43 -488 77 488
rect 301 -488 335 488
rect 421 -488 455 488
rect 679 -488 713 488
rect 799 -488 833 488
rect 1057 -488 1091 488
rect 1177 -488 1211 488
rect 1435 -488 1469 488
rect 1555 -488 1589 488
rect 1813 -488 1847 488
rect 1933 -488 1967 488
rect 2191 -488 2225 488
rect 2311 -488 2345 488
rect 2569 -488 2603 488
rect 2689 -488 2723 488
rect 2947 -488 2981 488
rect 3067 -488 3101 488
rect 3325 -488 3359 488
rect 3445 -488 3479 488
rect 3703 -488 3737 488
<< mvpsubdiff >>
rect -3883 710 3883 722
rect -3883 676 -3775 710
rect 3775 676 3883 710
rect -3883 664 3883 676
rect -3883 614 -3825 664
rect -3883 -614 -3871 614
rect -3837 -614 -3825 614
rect 3825 614 3883 664
rect -3883 -664 -3825 -614
rect 3825 -614 3837 614
rect 3871 -614 3883 614
rect 3825 -664 3883 -614
rect -3883 -676 3883 -664
rect -3883 -710 -3775 -676
rect 3775 -710 3883 -676
rect -3883 -722 3883 -710
<< mvpsubdiffcont >>
rect -3775 676 3775 710
rect -3871 -614 -3837 614
rect 3837 -614 3871 614
rect -3775 -710 3775 -676
<< poly >>
rect -3691 572 -3491 588
rect -3691 538 -3675 572
rect -3507 538 -3491 572
rect -3691 500 -3491 538
rect -3313 572 -3113 588
rect -3313 538 -3297 572
rect -3129 538 -3113 572
rect -3313 500 -3113 538
rect -2935 572 -2735 588
rect -2935 538 -2919 572
rect -2751 538 -2735 572
rect -2935 500 -2735 538
rect -2557 572 -2357 588
rect -2557 538 -2541 572
rect -2373 538 -2357 572
rect -2557 500 -2357 538
rect -2179 572 -1979 588
rect -2179 538 -2163 572
rect -1995 538 -1979 572
rect -2179 500 -1979 538
rect -1801 572 -1601 588
rect -1801 538 -1785 572
rect -1617 538 -1601 572
rect -1801 500 -1601 538
rect -1423 572 -1223 588
rect -1423 538 -1407 572
rect -1239 538 -1223 572
rect -1423 500 -1223 538
rect -1045 572 -845 588
rect -1045 538 -1029 572
rect -861 538 -845 572
rect -1045 500 -845 538
rect -667 572 -467 588
rect -667 538 -651 572
rect -483 538 -467 572
rect -667 500 -467 538
rect -289 572 -89 588
rect -289 538 -273 572
rect -105 538 -89 572
rect -289 500 -89 538
rect 89 572 289 588
rect 89 538 105 572
rect 273 538 289 572
rect 89 500 289 538
rect 467 572 667 588
rect 467 538 483 572
rect 651 538 667 572
rect 467 500 667 538
rect 845 572 1045 588
rect 845 538 861 572
rect 1029 538 1045 572
rect 845 500 1045 538
rect 1223 572 1423 588
rect 1223 538 1239 572
rect 1407 538 1423 572
rect 1223 500 1423 538
rect 1601 572 1801 588
rect 1601 538 1617 572
rect 1785 538 1801 572
rect 1601 500 1801 538
rect 1979 572 2179 588
rect 1979 538 1995 572
rect 2163 538 2179 572
rect 1979 500 2179 538
rect 2357 572 2557 588
rect 2357 538 2373 572
rect 2541 538 2557 572
rect 2357 500 2557 538
rect 2735 572 2935 588
rect 2735 538 2751 572
rect 2919 538 2935 572
rect 2735 500 2935 538
rect 3113 572 3313 588
rect 3113 538 3129 572
rect 3297 538 3313 572
rect 3113 500 3313 538
rect 3491 572 3691 588
rect 3491 538 3507 572
rect 3675 538 3691 572
rect 3491 500 3691 538
rect -3691 -538 -3491 -500
rect -3691 -572 -3675 -538
rect -3507 -572 -3491 -538
rect -3691 -588 -3491 -572
rect -3313 -538 -3113 -500
rect -3313 -572 -3297 -538
rect -3129 -572 -3113 -538
rect -3313 -588 -3113 -572
rect -2935 -538 -2735 -500
rect -2935 -572 -2919 -538
rect -2751 -572 -2735 -538
rect -2935 -588 -2735 -572
rect -2557 -538 -2357 -500
rect -2557 -572 -2541 -538
rect -2373 -572 -2357 -538
rect -2557 -588 -2357 -572
rect -2179 -538 -1979 -500
rect -2179 -572 -2163 -538
rect -1995 -572 -1979 -538
rect -2179 -588 -1979 -572
rect -1801 -538 -1601 -500
rect -1801 -572 -1785 -538
rect -1617 -572 -1601 -538
rect -1801 -588 -1601 -572
rect -1423 -538 -1223 -500
rect -1423 -572 -1407 -538
rect -1239 -572 -1223 -538
rect -1423 -588 -1223 -572
rect -1045 -538 -845 -500
rect -1045 -572 -1029 -538
rect -861 -572 -845 -538
rect -1045 -588 -845 -572
rect -667 -538 -467 -500
rect -667 -572 -651 -538
rect -483 -572 -467 -538
rect -667 -588 -467 -572
rect -289 -538 -89 -500
rect -289 -572 -273 -538
rect -105 -572 -89 -538
rect -289 -588 -89 -572
rect 89 -538 289 -500
rect 89 -572 105 -538
rect 273 -572 289 -538
rect 89 -588 289 -572
rect 467 -538 667 -500
rect 467 -572 483 -538
rect 651 -572 667 -538
rect 467 -588 667 -572
rect 845 -538 1045 -500
rect 845 -572 861 -538
rect 1029 -572 1045 -538
rect 845 -588 1045 -572
rect 1223 -538 1423 -500
rect 1223 -572 1239 -538
rect 1407 -572 1423 -538
rect 1223 -588 1423 -572
rect 1601 -538 1801 -500
rect 1601 -572 1617 -538
rect 1785 -572 1801 -538
rect 1601 -588 1801 -572
rect 1979 -538 2179 -500
rect 1979 -572 1995 -538
rect 2163 -572 2179 -538
rect 1979 -588 2179 -572
rect 2357 -538 2557 -500
rect 2357 -572 2373 -538
rect 2541 -572 2557 -538
rect 2357 -588 2557 -572
rect 2735 -538 2935 -500
rect 2735 -572 2751 -538
rect 2919 -572 2935 -538
rect 2735 -588 2935 -572
rect 3113 -538 3313 -500
rect 3113 -572 3129 -538
rect 3297 -572 3313 -538
rect 3113 -588 3313 -572
rect 3491 -538 3691 -500
rect 3491 -572 3507 -538
rect 3675 -572 3691 -538
rect 3491 -588 3691 -572
<< polycont >>
rect -3675 538 -3507 572
rect -3297 538 -3129 572
rect -2919 538 -2751 572
rect -2541 538 -2373 572
rect -2163 538 -1995 572
rect -1785 538 -1617 572
rect -1407 538 -1239 572
rect -1029 538 -861 572
rect -651 538 -483 572
rect -273 538 -105 572
rect 105 538 273 572
rect 483 538 651 572
rect 861 538 1029 572
rect 1239 538 1407 572
rect 1617 538 1785 572
rect 1995 538 2163 572
rect 2373 538 2541 572
rect 2751 538 2919 572
rect 3129 538 3297 572
rect 3507 538 3675 572
rect -3675 -572 -3507 -538
rect -3297 -572 -3129 -538
rect -2919 -572 -2751 -538
rect -2541 -572 -2373 -538
rect -2163 -572 -1995 -538
rect -1785 -572 -1617 -538
rect -1407 -572 -1239 -538
rect -1029 -572 -861 -538
rect -651 -572 -483 -538
rect -273 -572 -105 -538
rect 105 -572 273 -538
rect 483 -572 651 -538
rect 861 -572 1029 -538
rect 1239 -572 1407 -538
rect 1617 -572 1785 -538
rect 1995 -572 2163 -538
rect 2373 -572 2541 -538
rect 2751 -572 2919 -538
rect 3129 -572 3297 -538
rect 3507 -572 3675 -538
<< locali >>
rect -3871 676 -3775 710
rect 3775 676 3871 710
rect -3871 614 -3837 676
rect 3837 614 3871 676
rect -3691 538 -3675 572
rect -3507 538 -3491 572
rect -3313 538 -3297 572
rect -3129 538 -3113 572
rect -2935 538 -2919 572
rect -2751 538 -2735 572
rect -2557 538 -2541 572
rect -2373 538 -2357 572
rect -2179 538 -2163 572
rect -1995 538 -1979 572
rect -1801 538 -1785 572
rect -1617 538 -1601 572
rect -1423 538 -1407 572
rect -1239 538 -1223 572
rect -1045 538 -1029 572
rect -861 538 -845 572
rect -667 538 -651 572
rect -483 538 -467 572
rect -289 538 -273 572
rect -105 538 -89 572
rect 89 538 105 572
rect 273 538 289 572
rect 467 538 483 572
rect 651 538 667 572
rect 845 538 861 572
rect 1029 538 1045 572
rect 1223 538 1239 572
rect 1407 538 1423 572
rect 1601 538 1617 572
rect 1785 538 1801 572
rect 1979 538 1995 572
rect 2163 538 2179 572
rect 2357 538 2373 572
rect 2541 538 2557 572
rect 2735 538 2751 572
rect 2919 538 2935 572
rect 3113 538 3129 572
rect 3297 538 3313 572
rect 3491 538 3507 572
rect 3675 538 3691 572
rect -3737 488 -3703 504
rect -3737 -504 -3703 -488
rect -3479 488 -3445 504
rect -3479 -504 -3445 -488
rect -3359 488 -3325 504
rect -3359 -504 -3325 -488
rect -3101 488 -3067 504
rect -3101 -504 -3067 -488
rect -2981 488 -2947 504
rect -2981 -504 -2947 -488
rect -2723 488 -2689 504
rect -2723 -504 -2689 -488
rect -2603 488 -2569 504
rect -2603 -504 -2569 -488
rect -2345 488 -2311 504
rect -2345 -504 -2311 -488
rect -2225 488 -2191 504
rect -2225 -504 -2191 -488
rect -1967 488 -1933 504
rect -1967 -504 -1933 -488
rect -1847 488 -1813 504
rect -1847 -504 -1813 -488
rect -1589 488 -1555 504
rect -1589 -504 -1555 -488
rect -1469 488 -1435 504
rect -1469 -504 -1435 -488
rect -1211 488 -1177 504
rect -1211 -504 -1177 -488
rect -1091 488 -1057 504
rect -1091 -504 -1057 -488
rect -833 488 -799 504
rect -833 -504 -799 -488
rect -713 488 -679 504
rect -713 -504 -679 -488
rect -455 488 -421 504
rect -455 -504 -421 -488
rect -335 488 -301 504
rect -335 -504 -301 -488
rect -77 488 -43 504
rect -77 -504 -43 -488
rect 43 488 77 504
rect 43 -504 77 -488
rect 301 488 335 504
rect 301 -504 335 -488
rect 421 488 455 504
rect 421 -504 455 -488
rect 679 488 713 504
rect 679 -504 713 -488
rect 799 488 833 504
rect 799 -504 833 -488
rect 1057 488 1091 504
rect 1057 -504 1091 -488
rect 1177 488 1211 504
rect 1177 -504 1211 -488
rect 1435 488 1469 504
rect 1435 -504 1469 -488
rect 1555 488 1589 504
rect 1555 -504 1589 -488
rect 1813 488 1847 504
rect 1813 -504 1847 -488
rect 1933 488 1967 504
rect 1933 -504 1967 -488
rect 2191 488 2225 504
rect 2191 -504 2225 -488
rect 2311 488 2345 504
rect 2311 -504 2345 -488
rect 2569 488 2603 504
rect 2569 -504 2603 -488
rect 2689 488 2723 504
rect 2689 -504 2723 -488
rect 2947 488 2981 504
rect 2947 -504 2981 -488
rect 3067 488 3101 504
rect 3067 -504 3101 -488
rect 3325 488 3359 504
rect 3325 -504 3359 -488
rect 3445 488 3479 504
rect 3445 -504 3479 -488
rect 3703 488 3737 504
rect 3703 -504 3737 -488
rect -3691 -572 -3675 -538
rect -3507 -572 -3491 -538
rect -3313 -572 -3297 -538
rect -3129 -572 -3113 -538
rect -2935 -572 -2919 -538
rect -2751 -572 -2735 -538
rect -2557 -572 -2541 -538
rect -2373 -572 -2357 -538
rect -2179 -572 -2163 -538
rect -1995 -572 -1979 -538
rect -1801 -572 -1785 -538
rect -1617 -572 -1601 -538
rect -1423 -572 -1407 -538
rect -1239 -572 -1223 -538
rect -1045 -572 -1029 -538
rect -861 -572 -845 -538
rect -667 -572 -651 -538
rect -483 -572 -467 -538
rect -289 -572 -273 -538
rect -105 -572 -89 -538
rect 89 -572 105 -538
rect 273 -572 289 -538
rect 467 -572 483 -538
rect 651 -572 667 -538
rect 845 -572 861 -538
rect 1029 -572 1045 -538
rect 1223 -572 1239 -538
rect 1407 -572 1423 -538
rect 1601 -572 1617 -538
rect 1785 -572 1801 -538
rect 1979 -572 1995 -538
rect 2163 -572 2179 -538
rect 2357 -572 2373 -538
rect 2541 -572 2557 -538
rect 2735 -572 2751 -538
rect 2919 -572 2935 -538
rect 3113 -572 3129 -538
rect 3297 -572 3313 -538
rect 3491 -572 3507 -538
rect 3675 -572 3691 -538
rect -3871 -676 -3837 -614
rect 3837 -676 3871 -614
rect -3871 -710 -3775 -676
rect 3775 -710 3871 -676
<< viali >>
rect -3675 538 -3507 572
rect -3297 538 -3129 572
rect -2919 538 -2751 572
rect -2541 538 -2373 572
rect -2163 538 -1995 572
rect -1785 538 -1617 572
rect -1407 538 -1239 572
rect -1029 538 -861 572
rect -651 538 -483 572
rect -273 538 -105 572
rect 105 538 273 572
rect 483 538 651 572
rect 861 538 1029 572
rect 1239 538 1407 572
rect 1617 538 1785 572
rect 1995 538 2163 572
rect 2373 538 2541 572
rect 2751 538 2919 572
rect 3129 538 3297 572
rect 3507 538 3675 572
rect -3737 -488 -3703 488
rect -3479 -488 -3445 488
rect -3359 -488 -3325 488
rect -3101 -488 -3067 488
rect -2981 -488 -2947 488
rect -2723 -488 -2689 488
rect -2603 -488 -2569 488
rect -2345 -488 -2311 488
rect -2225 -488 -2191 488
rect -1967 -488 -1933 488
rect -1847 -488 -1813 488
rect -1589 -488 -1555 488
rect -1469 -488 -1435 488
rect -1211 -488 -1177 488
rect -1091 -488 -1057 488
rect -833 -488 -799 488
rect -713 -488 -679 488
rect -455 -488 -421 488
rect -335 -488 -301 488
rect -77 -488 -43 488
rect 43 -488 77 488
rect 301 -488 335 488
rect 421 -488 455 488
rect 679 -488 713 488
rect 799 -488 833 488
rect 1057 -488 1091 488
rect 1177 -488 1211 488
rect 1435 -488 1469 488
rect 1555 -488 1589 488
rect 1813 -488 1847 488
rect 1933 -488 1967 488
rect 2191 -488 2225 488
rect 2311 -488 2345 488
rect 2569 -488 2603 488
rect 2689 -488 2723 488
rect 2947 -488 2981 488
rect 3067 -488 3101 488
rect 3325 -488 3359 488
rect 3445 -488 3479 488
rect 3703 -488 3737 488
rect -3675 -572 -3507 -538
rect -3297 -572 -3129 -538
rect -2919 -572 -2751 -538
rect -2541 -572 -2373 -538
rect -2163 -572 -1995 -538
rect -1785 -572 -1617 -538
rect -1407 -572 -1239 -538
rect -1029 -572 -861 -538
rect -651 -572 -483 -538
rect -273 -572 -105 -538
rect 105 -572 273 -538
rect 483 -572 651 -538
rect 861 -572 1029 -538
rect 1239 -572 1407 -538
rect 1617 -572 1785 -538
rect 1995 -572 2163 -538
rect 2373 -572 2541 -538
rect 2751 -572 2919 -538
rect 3129 -572 3297 -538
rect 3507 -572 3675 -538
<< metal1 >>
rect -3687 572 -3495 578
rect -3687 538 -3675 572
rect -3507 538 -3495 572
rect -3687 532 -3495 538
rect -3309 572 -3117 578
rect -3309 538 -3297 572
rect -3129 538 -3117 572
rect -3309 532 -3117 538
rect -2931 572 -2739 578
rect -2931 538 -2919 572
rect -2751 538 -2739 572
rect -2931 532 -2739 538
rect -2553 572 -2361 578
rect -2553 538 -2541 572
rect -2373 538 -2361 572
rect -2553 532 -2361 538
rect -2175 572 -1983 578
rect -2175 538 -2163 572
rect -1995 538 -1983 572
rect -2175 532 -1983 538
rect -1797 572 -1605 578
rect -1797 538 -1785 572
rect -1617 538 -1605 572
rect -1797 532 -1605 538
rect -1419 572 -1227 578
rect -1419 538 -1407 572
rect -1239 538 -1227 572
rect -1419 532 -1227 538
rect -1041 572 -849 578
rect -1041 538 -1029 572
rect -861 538 -849 572
rect -1041 532 -849 538
rect -663 572 -471 578
rect -663 538 -651 572
rect -483 538 -471 572
rect -663 532 -471 538
rect -285 572 -93 578
rect -285 538 -273 572
rect -105 538 -93 572
rect -285 532 -93 538
rect 93 572 285 578
rect 93 538 105 572
rect 273 538 285 572
rect 93 532 285 538
rect 471 572 663 578
rect 471 538 483 572
rect 651 538 663 572
rect 471 532 663 538
rect 849 572 1041 578
rect 849 538 861 572
rect 1029 538 1041 572
rect 849 532 1041 538
rect 1227 572 1419 578
rect 1227 538 1239 572
rect 1407 538 1419 572
rect 1227 532 1419 538
rect 1605 572 1797 578
rect 1605 538 1617 572
rect 1785 538 1797 572
rect 1605 532 1797 538
rect 1983 572 2175 578
rect 1983 538 1995 572
rect 2163 538 2175 572
rect 1983 532 2175 538
rect 2361 572 2553 578
rect 2361 538 2373 572
rect 2541 538 2553 572
rect 2361 532 2553 538
rect 2739 572 2931 578
rect 2739 538 2751 572
rect 2919 538 2931 572
rect 2739 532 2931 538
rect 3117 572 3309 578
rect 3117 538 3129 572
rect 3297 538 3309 572
rect 3117 532 3309 538
rect 3495 572 3687 578
rect 3495 538 3507 572
rect 3675 538 3687 572
rect 3495 532 3687 538
rect -3743 488 -3697 500
rect -3743 -488 -3737 488
rect -3703 -488 -3697 488
rect -3743 -500 -3697 -488
rect -3485 488 -3439 500
rect -3485 -488 -3479 488
rect -3445 -488 -3439 488
rect -3485 -500 -3439 -488
rect -3365 488 -3319 500
rect -3365 -488 -3359 488
rect -3325 -488 -3319 488
rect -3365 -500 -3319 -488
rect -3107 488 -3061 500
rect -3107 -488 -3101 488
rect -3067 -488 -3061 488
rect -3107 -500 -3061 -488
rect -2987 488 -2941 500
rect -2987 -488 -2981 488
rect -2947 -488 -2941 488
rect -2987 -500 -2941 -488
rect -2729 488 -2683 500
rect -2729 -488 -2723 488
rect -2689 -488 -2683 488
rect -2729 -500 -2683 -488
rect -2609 488 -2563 500
rect -2609 -488 -2603 488
rect -2569 -488 -2563 488
rect -2609 -500 -2563 -488
rect -2351 488 -2305 500
rect -2351 -488 -2345 488
rect -2311 -488 -2305 488
rect -2351 -500 -2305 -488
rect -2231 488 -2185 500
rect -2231 -488 -2225 488
rect -2191 -488 -2185 488
rect -2231 -500 -2185 -488
rect -1973 488 -1927 500
rect -1973 -488 -1967 488
rect -1933 -488 -1927 488
rect -1973 -500 -1927 -488
rect -1853 488 -1807 500
rect -1853 -488 -1847 488
rect -1813 -488 -1807 488
rect -1853 -500 -1807 -488
rect -1595 488 -1549 500
rect -1595 -488 -1589 488
rect -1555 -488 -1549 488
rect -1595 -500 -1549 -488
rect -1475 488 -1429 500
rect -1475 -488 -1469 488
rect -1435 -488 -1429 488
rect -1475 -500 -1429 -488
rect -1217 488 -1171 500
rect -1217 -488 -1211 488
rect -1177 -488 -1171 488
rect -1217 -500 -1171 -488
rect -1097 488 -1051 500
rect -1097 -488 -1091 488
rect -1057 -488 -1051 488
rect -1097 -500 -1051 -488
rect -839 488 -793 500
rect -839 -488 -833 488
rect -799 -488 -793 488
rect -839 -500 -793 -488
rect -719 488 -673 500
rect -719 -488 -713 488
rect -679 -488 -673 488
rect -719 -500 -673 -488
rect -461 488 -415 500
rect -461 -488 -455 488
rect -421 -488 -415 488
rect -461 -500 -415 -488
rect -341 488 -295 500
rect -341 -488 -335 488
rect -301 -488 -295 488
rect -341 -500 -295 -488
rect -83 488 -37 500
rect -83 -488 -77 488
rect -43 -488 -37 488
rect -83 -500 -37 -488
rect 37 488 83 500
rect 37 -488 43 488
rect 77 -488 83 488
rect 37 -500 83 -488
rect 295 488 341 500
rect 295 -488 301 488
rect 335 -488 341 488
rect 295 -500 341 -488
rect 415 488 461 500
rect 415 -488 421 488
rect 455 -488 461 488
rect 415 -500 461 -488
rect 673 488 719 500
rect 673 -488 679 488
rect 713 -488 719 488
rect 673 -500 719 -488
rect 793 488 839 500
rect 793 -488 799 488
rect 833 -488 839 488
rect 793 -500 839 -488
rect 1051 488 1097 500
rect 1051 -488 1057 488
rect 1091 -488 1097 488
rect 1051 -500 1097 -488
rect 1171 488 1217 500
rect 1171 -488 1177 488
rect 1211 -488 1217 488
rect 1171 -500 1217 -488
rect 1429 488 1475 500
rect 1429 -488 1435 488
rect 1469 -488 1475 488
rect 1429 -500 1475 -488
rect 1549 488 1595 500
rect 1549 -488 1555 488
rect 1589 -488 1595 488
rect 1549 -500 1595 -488
rect 1807 488 1853 500
rect 1807 -488 1813 488
rect 1847 -488 1853 488
rect 1807 -500 1853 -488
rect 1927 488 1973 500
rect 1927 -488 1933 488
rect 1967 -488 1973 488
rect 1927 -500 1973 -488
rect 2185 488 2231 500
rect 2185 -488 2191 488
rect 2225 -488 2231 488
rect 2185 -500 2231 -488
rect 2305 488 2351 500
rect 2305 -488 2311 488
rect 2345 -488 2351 488
rect 2305 -500 2351 -488
rect 2563 488 2609 500
rect 2563 -488 2569 488
rect 2603 -488 2609 488
rect 2563 -500 2609 -488
rect 2683 488 2729 500
rect 2683 -488 2689 488
rect 2723 -488 2729 488
rect 2683 -500 2729 -488
rect 2941 488 2987 500
rect 2941 -488 2947 488
rect 2981 -488 2987 488
rect 2941 -500 2987 -488
rect 3061 488 3107 500
rect 3061 -488 3067 488
rect 3101 -488 3107 488
rect 3061 -500 3107 -488
rect 3319 488 3365 500
rect 3319 -488 3325 488
rect 3359 -488 3365 488
rect 3319 -500 3365 -488
rect 3439 488 3485 500
rect 3439 -488 3445 488
rect 3479 -488 3485 488
rect 3439 -500 3485 -488
rect 3697 488 3743 500
rect 3697 -488 3703 488
rect 3737 -488 3743 488
rect 3697 -500 3743 -488
rect -3687 -538 -3495 -532
rect -3687 -572 -3675 -538
rect -3507 -572 -3495 -538
rect -3687 -578 -3495 -572
rect -3309 -538 -3117 -532
rect -3309 -572 -3297 -538
rect -3129 -572 -3117 -538
rect -3309 -578 -3117 -572
rect -2931 -538 -2739 -532
rect -2931 -572 -2919 -538
rect -2751 -572 -2739 -538
rect -2931 -578 -2739 -572
rect -2553 -538 -2361 -532
rect -2553 -572 -2541 -538
rect -2373 -572 -2361 -538
rect -2553 -578 -2361 -572
rect -2175 -538 -1983 -532
rect -2175 -572 -2163 -538
rect -1995 -572 -1983 -538
rect -2175 -578 -1983 -572
rect -1797 -538 -1605 -532
rect -1797 -572 -1785 -538
rect -1617 -572 -1605 -538
rect -1797 -578 -1605 -572
rect -1419 -538 -1227 -532
rect -1419 -572 -1407 -538
rect -1239 -572 -1227 -538
rect -1419 -578 -1227 -572
rect -1041 -538 -849 -532
rect -1041 -572 -1029 -538
rect -861 -572 -849 -538
rect -1041 -578 -849 -572
rect -663 -538 -471 -532
rect -663 -572 -651 -538
rect -483 -572 -471 -538
rect -663 -578 -471 -572
rect -285 -538 -93 -532
rect -285 -572 -273 -538
rect -105 -572 -93 -538
rect -285 -578 -93 -572
rect 93 -538 285 -532
rect 93 -572 105 -538
rect 273 -572 285 -538
rect 93 -578 285 -572
rect 471 -538 663 -532
rect 471 -572 483 -538
rect 651 -572 663 -538
rect 471 -578 663 -572
rect 849 -538 1041 -532
rect 849 -572 861 -538
rect 1029 -572 1041 -538
rect 849 -578 1041 -572
rect 1227 -538 1419 -532
rect 1227 -572 1239 -538
rect 1407 -572 1419 -538
rect 1227 -578 1419 -572
rect 1605 -538 1797 -532
rect 1605 -572 1617 -538
rect 1785 -572 1797 -538
rect 1605 -578 1797 -572
rect 1983 -538 2175 -532
rect 1983 -572 1995 -538
rect 2163 -572 2175 -538
rect 1983 -578 2175 -572
rect 2361 -538 2553 -532
rect 2361 -572 2373 -538
rect 2541 -572 2553 -538
rect 2361 -578 2553 -572
rect 2739 -538 2931 -532
rect 2739 -572 2751 -538
rect 2919 -572 2931 -538
rect 2739 -578 2931 -572
rect 3117 -538 3309 -532
rect 3117 -572 3129 -538
rect 3297 -572 3309 -538
rect 3117 -578 3309 -572
rect 3495 -538 3687 -532
rect 3495 -572 3507 -538
rect 3675 -572 3687 -538
rect 3495 -578 3687 -572
<< properties >>
string FIXED_BBOX -3854 -693 3854 693
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 1.0 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
