magic
tech sky130A
magscale 1 2
timestamp 1730992408
<< locali >>
rect 896 -500 992 -300
rect 884 -1802 986 -1602
<< metal1 >>
rect 704 -260 904 -134
rect 562 -938 646 -550
rect 718 -816 766 -260
rect 562 -1138 658 -938
rect 820 -952 904 -550
rect 562 -1556 646 -1138
rect 794 -1152 904 -952
rect 706 -1830 754 -1286
rect 820 -1556 904 -1152
rect 704 -1926 904 -1830
use sky130_fd_pr__nfet_g5v0d10v5_92HZNS  XM1 paramcells
timestamp 1730992408
transform 1 0 740 0 1 -646
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_TUFYNQ  XM2 paramcells
timestamp 1730992408
transform 1 0 730 0 1 -1459
box -308 -397 308 397
<< labels >>
flabel metal1 704 -260 904 -134 0 FreeSans 256 0 0 0 NGATE
port 2 nsew
flabel metal1 704 -1926 904 -1830 0 FreeSans 256 0 0 0 PGATE
port 1 nsew
flabel metal1 796 -1152 904 -952 0 FreeSans 256 0 0 0 LOWER
port 3 nsew
flabel metal1 562 -1138 656 -938 0 FreeSans 256 0 0 0 UPPER
port 0 nsew
flabel locali 884 -1802 986 -1602 0 FreeSans 256 0 0 0 AVDD
port 5 nsew
flabel locali 896 -500 992 -300 0 FreeSans 256 0 0 0 AVSS
port 4 nsew
<< end >>
