magic
tech sky130A
magscale 1 2
timestamp 1729620069
<< pwell >>
rect -4864 -2585 4864 2585
<< mvnmos >>
rect -4636 1327 -4436 2327
rect -4258 1327 -4058 2327
rect -3880 1327 -3680 2327
rect -3502 1327 -3302 2327
rect -3124 1327 -2924 2327
rect -2746 1327 -2546 2327
rect -2368 1327 -2168 2327
rect -1990 1327 -1790 2327
rect -1612 1327 -1412 2327
rect -1234 1327 -1034 2327
rect -856 1327 -656 2327
rect -478 1327 -278 2327
rect -100 1327 100 2327
rect 278 1327 478 2327
rect 656 1327 856 2327
rect 1034 1327 1234 2327
rect 1412 1327 1612 2327
rect 1790 1327 1990 2327
rect 2168 1327 2368 2327
rect 2546 1327 2746 2327
rect 2924 1327 3124 2327
rect 3302 1327 3502 2327
rect 3680 1327 3880 2327
rect 4058 1327 4258 2327
rect 4436 1327 4636 2327
rect -4636 109 -4436 1109
rect -4258 109 -4058 1109
rect -3880 109 -3680 1109
rect -3502 109 -3302 1109
rect -3124 109 -2924 1109
rect -2746 109 -2546 1109
rect -2368 109 -2168 1109
rect -1990 109 -1790 1109
rect -1612 109 -1412 1109
rect -1234 109 -1034 1109
rect -856 109 -656 1109
rect -478 109 -278 1109
rect -100 109 100 1109
rect 278 109 478 1109
rect 656 109 856 1109
rect 1034 109 1234 1109
rect 1412 109 1612 1109
rect 1790 109 1990 1109
rect 2168 109 2368 1109
rect 2546 109 2746 1109
rect 2924 109 3124 1109
rect 3302 109 3502 1109
rect 3680 109 3880 1109
rect 4058 109 4258 1109
rect 4436 109 4636 1109
rect -4636 -1109 -4436 -109
rect -4258 -1109 -4058 -109
rect -3880 -1109 -3680 -109
rect -3502 -1109 -3302 -109
rect -3124 -1109 -2924 -109
rect -2746 -1109 -2546 -109
rect -2368 -1109 -2168 -109
rect -1990 -1109 -1790 -109
rect -1612 -1109 -1412 -109
rect -1234 -1109 -1034 -109
rect -856 -1109 -656 -109
rect -478 -1109 -278 -109
rect -100 -1109 100 -109
rect 278 -1109 478 -109
rect 656 -1109 856 -109
rect 1034 -1109 1234 -109
rect 1412 -1109 1612 -109
rect 1790 -1109 1990 -109
rect 2168 -1109 2368 -109
rect 2546 -1109 2746 -109
rect 2924 -1109 3124 -109
rect 3302 -1109 3502 -109
rect 3680 -1109 3880 -109
rect 4058 -1109 4258 -109
rect 4436 -1109 4636 -109
rect -4636 -2327 -4436 -1327
rect -4258 -2327 -4058 -1327
rect -3880 -2327 -3680 -1327
rect -3502 -2327 -3302 -1327
rect -3124 -2327 -2924 -1327
rect -2746 -2327 -2546 -1327
rect -2368 -2327 -2168 -1327
rect -1990 -2327 -1790 -1327
rect -1612 -2327 -1412 -1327
rect -1234 -2327 -1034 -1327
rect -856 -2327 -656 -1327
rect -478 -2327 -278 -1327
rect -100 -2327 100 -1327
rect 278 -2327 478 -1327
rect 656 -2327 856 -1327
rect 1034 -2327 1234 -1327
rect 1412 -2327 1612 -1327
rect 1790 -2327 1990 -1327
rect 2168 -2327 2368 -1327
rect 2546 -2327 2746 -1327
rect 2924 -2327 3124 -1327
rect 3302 -2327 3502 -1327
rect 3680 -2327 3880 -1327
rect 4058 -2327 4258 -1327
rect 4436 -2327 4636 -1327
<< mvndiff >>
rect -4694 2315 -4636 2327
rect -4694 1339 -4682 2315
rect -4648 1339 -4636 2315
rect -4694 1327 -4636 1339
rect -4436 2315 -4378 2327
rect -4436 1339 -4424 2315
rect -4390 1339 -4378 2315
rect -4436 1327 -4378 1339
rect -4316 2315 -4258 2327
rect -4316 1339 -4304 2315
rect -4270 1339 -4258 2315
rect -4316 1327 -4258 1339
rect -4058 2315 -4000 2327
rect -4058 1339 -4046 2315
rect -4012 1339 -4000 2315
rect -4058 1327 -4000 1339
rect -3938 2315 -3880 2327
rect -3938 1339 -3926 2315
rect -3892 1339 -3880 2315
rect -3938 1327 -3880 1339
rect -3680 2315 -3622 2327
rect -3680 1339 -3668 2315
rect -3634 1339 -3622 2315
rect -3680 1327 -3622 1339
rect -3560 2315 -3502 2327
rect -3560 1339 -3548 2315
rect -3514 1339 -3502 2315
rect -3560 1327 -3502 1339
rect -3302 2315 -3244 2327
rect -3302 1339 -3290 2315
rect -3256 1339 -3244 2315
rect -3302 1327 -3244 1339
rect -3182 2315 -3124 2327
rect -3182 1339 -3170 2315
rect -3136 1339 -3124 2315
rect -3182 1327 -3124 1339
rect -2924 2315 -2866 2327
rect -2924 1339 -2912 2315
rect -2878 1339 -2866 2315
rect -2924 1327 -2866 1339
rect -2804 2315 -2746 2327
rect -2804 1339 -2792 2315
rect -2758 1339 -2746 2315
rect -2804 1327 -2746 1339
rect -2546 2315 -2488 2327
rect -2546 1339 -2534 2315
rect -2500 1339 -2488 2315
rect -2546 1327 -2488 1339
rect -2426 2315 -2368 2327
rect -2426 1339 -2414 2315
rect -2380 1339 -2368 2315
rect -2426 1327 -2368 1339
rect -2168 2315 -2110 2327
rect -2168 1339 -2156 2315
rect -2122 1339 -2110 2315
rect -2168 1327 -2110 1339
rect -2048 2315 -1990 2327
rect -2048 1339 -2036 2315
rect -2002 1339 -1990 2315
rect -2048 1327 -1990 1339
rect -1790 2315 -1732 2327
rect -1790 1339 -1778 2315
rect -1744 1339 -1732 2315
rect -1790 1327 -1732 1339
rect -1670 2315 -1612 2327
rect -1670 1339 -1658 2315
rect -1624 1339 -1612 2315
rect -1670 1327 -1612 1339
rect -1412 2315 -1354 2327
rect -1412 1339 -1400 2315
rect -1366 1339 -1354 2315
rect -1412 1327 -1354 1339
rect -1292 2315 -1234 2327
rect -1292 1339 -1280 2315
rect -1246 1339 -1234 2315
rect -1292 1327 -1234 1339
rect -1034 2315 -976 2327
rect -1034 1339 -1022 2315
rect -988 1339 -976 2315
rect -1034 1327 -976 1339
rect -914 2315 -856 2327
rect -914 1339 -902 2315
rect -868 1339 -856 2315
rect -914 1327 -856 1339
rect -656 2315 -598 2327
rect -656 1339 -644 2315
rect -610 1339 -598 2315
rect -656 1327 -598 1339
rect -536 2315 -478 2327
rect -536 1339 -524 2315
rect -490 1339 -478 2315
rect -536 1327 -478 1339
rect -278 2315 -220 2327
rect -278 1339 -266 2315
rect -232 1339 -220 2315
rect -278 1327 -220 1339
rect -158 2315 -100 2327
rect -158 1339 -146 2315
rect -112 1339 -100 2315
rect -158 1327 -100 1339
rect 100 2315 158 2327
rect 100 1339 112 2315
rect 146 1339 158 2315
rect 100 1327 158 1339
rect 220 2315 278 2327
rect 220 1339 232 2315
rect 266 1339 278 2315
rect 220 1327 278 1339
rect 478 2315 536 2327
rect 478 1339 490 2315
rect 524 1339 536 2315
rect 478 1327 536 1339
rect 598 2315 656 2327
rect 598 1339 610 2315
rect 644 1339 656 2315
rect 598 1327 656 1339
rect 856 2315 914 2327
rect 856 1339 868 2315
rect 902 1339 914 2315
rect 856 1327 914 1339
rect 976 2315 1034 2327
rect 976 1339 988 2315
rect 1022 1339 1034 2315
rect 976 1327 1034 1339
rect 1234 2315 1292 2327
rect 1234 1339 1246 2315
rect 1280 1339 1292 2315
rect 1234 1327 1292 1339
rect 1354 2315 1412 2327
rect 1354 1339 1366 2315
rect 1400 1339 1412 2315
rect 1354 1327 1412 1339
rect 1612 2315 1670 2327
rect 1612 1339 1624 2315
rect 1658 1339 1670 2315
rect 1612 1327 1670 1339
rect 1732 2315 1790 2327
rect 1732 1339 1744 2315
rect 1778 1339 1790 2315
rect 1732 1327 1790 1339
rect 1990 2315 2048 2327
rect 1990 1339 2002 2315
rect 2036 1339 2048 2315
rect 1990 1327 2048 1339
rect 2110 2315 2168 2327
rect 2110 1339 2122 2315
rect 2156 1339 2168 2315
rect 2110 1327 2168 1339
rect 2368 2315 2426 2327
rect 2368 1339 2380 2315
rect 2414 1339 2426 2315
rect 2368 1327 2426 1339
rect 2488 2315 2546 2327
rect 2488 1339 2500 2315
rect 2534 1339 2546 2315
rect 2488 1327 2546 1339
rect 2746 2315 2804 2327
rect 2746 1339 2758 2315
rect 2792 1339 2804 2315
rect 2746 1327 2804 1339
rect 2866 2315 2924 2327
rect 2866 1339 2878 2315
rect 2912 1339 2924 2315
rect 2866 1327 2924 1339
rect 3124 2315 3182 2327
rect 3124 1339 3136 2315
rect 3170 1339 3182 2315
rect 3124 1327 3182 1339
rect 3244 2315 3302 2327
rect 3244 1339 3256 2315
rect 3290 1339 3302 2315
rect 3244 1327 3302 1339
rect 3502 2315 3560 2327
rect 3502 1339 3514 2315
rect 3548 1339 3560 2315
rect 3502 1327 3560 1339
rect 3622 2315 3680 2327
rect 3622 1339 3634 2315
rect 3668 1339 3680 2315
rect 3622 1327 3680 1339
rect 3880 2315 3938 2327
rect 3880 1339 3892 2315
rect 3926 1339 3938 2315
rect 3880 1327 3938 1339
rect 4000 2315 4058 2327
rect 4000 1339 4012 2315
rect 4046 1339 4058 2315
rect 4000 1327 4058 1339
rect 4258 2315 4316 2327
rect 4258 1339 4270 2315
rect 4304 1339 4316 2315
rect 4258 1327 4316 1339
rect 4378 2315 4436 2327
rect 4378 1339 4390 2315
rect 4424 1339 4436 2315
rect 4378 1327 4436 1339
rect 4636 2315 4694 2327
rect 4636 1339 4648 2315
rect 4682 1339 4694 2315
rect 4636 1327 4694 1339
rect -4694 1097 -4636 1109
rect -4694 121 -4682 1097
rect -4648 121 -4636 1097
rect -4694 109 -4636 121
rect -4436 1097 -4378 1109
rect -4436 121 -4424 1097
rect -4390 121 -4378 1097
rect -4436 109 -4378 121
rect -4316 1097 -4258 1109
rect -4316 121 -4304 1097
rect -4270 121 -4258 1097
rect -4316 109 -4258 121
rect -4058 1097 -4000 1109
rect -4058 121 -4046 1097
rect -4012 121 -4000 1097
rect -4058 109 -4000 121
rect -3938 1097 -3880 1109
rect -3938 121 -3926 1097
rect -3892 121 -3880 1097
rect -3938 109 -3880 121
rect -3680 1097 -3622 1109
rect -3680 121 -3668 1097
rect -3634 121 -3622 1097
rect -3680 109 -3622 121
rect -3560 1097 -3502 1109
rect -3560 121 -3548 1097
rect -3514 121 -3502 1097
rect -3560 109 -3502 121
rect -3302 1097 -3244 1109
rect -3302 121 -3290 1097
rect -3256 121 -3244 1097
rect -3302 109 -3244 121
rect -3182 1097 -3124 1109
rect -3182 121 -3170 1097
rect -3136 121 -3124 1097
rect -3182 109 -3124 121
rect -2924 1097 -2866 1109
rect -2924 121 -2912 1097
rect -2878 121 -2866 1097
rect -2924 109 -2866 121
rect -2804 1097 -2746 1109
rect -2804 121 -2792 1097
rect -2758 121 -2746 1097
rect -2804 109 -2746 121
rect -2546 1097 -2488 1109
rect -2546 121 -2534 1097
rect -2500 121 -2488 1097
rect -2546 109 -2488 121
rect -2426 1097 -2368 1109
rect -2426 121 -2414 1097
rect -2380 121 -2368 1097
rect -2426 109 -2368 121
rect -2168 1097 -2110 1109
rect -2168 121 -2156 1097
rect -2122 121 -2110 1097
rect -2168 109 -2110 121
rect -2048 1097 -1990 1109
rect -2048 121 -2036 1097
rect -2002 121 -1990 1097
rect -2048 109 -1990 121
rect -1790 1097 -1732 1109
rect -1790 121 -1778 1097
rect -1744 121 -1732 1097
rect -1790 109 -1732 121
rect -1670 1097 -1612 1109
rect -1670 121 -1658 1097
rect -1624 121 -1612 1097
rect -1670 109 -1612 121
rect -1412 1097 -1354 1109
rect -1412 121 -1400 1097
rect -1366 121 -1354 1097
rect -1412 109 -1354 121
rect -1292 1097 -1234 1109
rect -1292 121 -1280 1097
rect -1246 121 -1234 1097
rect -1292 109 -1234 121
rect -1034 1097 -976 1109
rect -1034 121 -1022 1097
rect -988 121 -976 1097
rect -1034 109 -976 121
rect -914 1097 -856 1109
rect -914 121 -902 1097
rect -868 121 -856 1097
rect -914 109 -856 121
rect -656 1097 -598 1109
rect -656 121 -644 1097
rect -610 121 -598 1097
rect -656 109 -598 121
rect -536 1097 -478 1109
rect -536 121 -524 1097
rect -490 121 -478 1097
rect -536 109 -478 121
rect -278 1097 -220 1109
rect -278 121 -266 1097
rect -232 121 -220 1097
rect -278 109 -220 121
rect -158 1097 -100 1109
rect -158 121 -146 1097
rect -112 121 -100 1097
rect -158 109 -100 121
rect 100 1097 158 1109
rect 100 121 112 1097
rect 146 121 158 1097
rect 100 109 158 121
rect 220 1097 278 1109
rect 220 121 232 1097
rect 266 121 278 1097
rect 220 109 278 121
rect 478 1097 536 1109
rect 478 121 490 1097
rect 524 121 536 1097
rect 478 109 536 121
rect 598 1097 656 1109
rect 598 121 610 1097
rect 644 121 656 1097
rect 598 109 656 121
rect 856 1097 914 1109
rect 856 121 868 1097
rect 902 121 914 1097
rect 856 109 914 121
rect 976 1097 1034 1109
rect 976 121 988 1097
rect 1022 121 1034 1097
rect 976 109 1034 121
rect 1234 1097 1292 1109
rect 1234 121 1246 1097
rect 1280 121 1292 1097
rect 1234 109 1292 121
rect 1354 1097 1412 1109
rect 1354 121 1366 1097
rect 1400 121 1412 1097
rect 1354 109 1412 121
rect 1612 1097 1670 1109
rect 1612 121 1624 1097
rect 1658 121 1670 1097
rect 1612 109 1670 121
rect 1732 1097 1790 1109
rect 1732 121 1744 1097
rect 1778 121 1790 1097
rect 1732 109 1790 121
rect 1990 1097 2048 1109
rect 1990 121 2002 1097
rect 2036 121 2048 1097
rect 1990 109 2048 121
rect 2110 1097 2168 1109
rect 2110 121 2122 1097
rect 2156 121 2168 1097
rect 2110 109 2168 121
rect 2368 1097 2426 1109
rect 2368 121 2380 1097
rect 2414 121 2426 1097
rect 2368 109 2426 121
rect 2488 1097 2546 1109
rect 2488 121 2500 1097
rect 2534 121 2546 1097
rect 2488 109 2546 121
rect 2746 1097 2804 1109
rect 2746 121 2758 1097
rect 2792 121 2804 1097
rect 2746 109 2804 121
rect 2866 1097 2924 1109
rect 2866 121 2878 1097
rect 2912 121 2924 1097
rect 2866 109 2924 121
rect 3124 1097 3182 1109
rect 3124 121 3136 1097
rect 3170 121 3182 1097
rect 3124 109 3182 121
rect 3244 1097 3302 1109
rect 3244 121 3256 1097
rect 3290 121 3302 1097
rect 3244 109 3302 121
rect 3502 1097 3560 1109
rect 3502 121 3514 1097
rect 3548 121 3560 1097
rect 3502 109 3560 121
rect 3622 1097 3680 1109
rect 3622 121 3634 1097
rect 3668 121 3680 1097
rect 3622 109 3680 121
rect 3880 1097 3938 1109
rect 3880 121 3892 1097
rect 3926 121 3938 1097
rect 3880 109 3938 121
rect 4000 1097 4058 1109
rect 4000 121 4012 1097
rect 4046 121 4058 1097
rect 4000 109 4058 121
rect 4258 1097 4316 1109
rect 4258 121 4270 1097
rect 4304 121 4316 1097
rect 4258 109 4316 121
rect 4378 1097 4436 1109
rect 4378 121 4390 1097
rect 4424 121 4436 1097
rect 4378 109 4436 121
rect 4636 1097 4694 1109
rect 4636 121 4648 1097
rect 4682 121 4694 1097
rect 4636 109 4694 121
rect -4694 -121 -4636 -109
rect -4694 -1097 -4682 -121
rect -4648 -1097 -4636 -121
rect -4694 -1109 -4636 -1097
rect -4436 -121 -4378 -109
rect -4436 -1097 -4424 -121
rect -4390 -1097 -4378 -121
rect -4436 -1109 -4378 -1097
rect -4316 -121 -4258 -109
rect -4316 -1097 -4304 -121
rect -4270 -1097 -4258 -121
rect -4316 -1109 -4258 -1097
rect -4058 -121 -4000 -109
rect -4058 -1097 -4046 -121
rect -4012 -1097 -4000 -121
rect -4058 -1109 -4000 -1097
rect -3938 -121 -3880 -109
rect -3938 -1097 -3926 -121
rect -3892 -1097 -3880 -121
rect -3938 -1109 -3880 -1097
rect -3680 -121 -3622 -109
rect -3680 -1097 -3668 -121
rect -3634 -1097 -3622 -121
rect -3680 -1109 -3622 -1097
rect -3560 -121 -3502 -109
rect -3560 -1097 -3548 -121
rect -3514 -1097 -3502 -121
rect -3560 -1109 -3502 -1097
rect -3302 -121 -3244 -109
rect -3302 -1097 -3290 -121
rect -3256 -1097 -3244 -121
rect -3302 -1109 -3244 -1097
rect -3182 -121 -3124 -109
rect -3182 -1097 -3170 -121
rect -3136 -1097 -3124 -121
rect -3182 -1109 -3124 -1097
rect -2924 -121 -2866 -109
rect -2924 -1097 -2912 -121
rect -2878 -1097 -2866 -121
rect -2924 -1109 -2866 -1097
rect -2804 -121 -2746 -109
rect -2804 -1097 -2792 -121
rect -2758 -1097 -2746 -121
rect -2804 -1109 -2746 -1097
rect -2546 -121 -2488 -109
rect -2546 -1097 -2534 -121
rect -2500 -1097 -2488 -121
rect -2546 -1109 -2488 -1097
rect -2426 -121 -2368 -109
rect -2426 -1097 -2414 -121
rect -2380 -1097 -2368 -121
rect -2426 -1109 -2368 -1097
rect -2168 -121 -2110 -109
rect -2168 -1097 -2156 -121
rect -2122 -1097 -2110 -121
rect -2168 -1109 -2110 -1097
rect -2048 -121 -1990 -109
rect -2048 -1097 -2036 -121
rect -2002 -1097 -1990 -121
rect -2048 -1109 -1990 -1097
rect -1790 -121 -1732 -109
rect -1790 -1097 -1778 -121
rect -1744 -1097 -1732 -121
rect -1790 -1109 -1732 -1097
rect -1670 -121 -1612 -109
rect -1670 -1097 -1658 -121
rect -1624 -1097 -1612 -121
rect -1670 -1109 -1612 -1097
rect -1412 -121 -1354 -109
rect -1412 -1097 -1400 -121
rect -1366 -1097 -1354 -121
rect -1412 -1109 -1354 -1097
rect -1292 -121 -1234 -109
rect -1292 -1097 -1280 -121
rect -1246 -1097 -1234 -121
rect -1292 -1109 -1234 -1097
rect -1034 -121 -976 -109
rect -1034 -1097 -1022 -121
rect -988 -1097 -976 -121
rect -1034 -1109 -976 -1097
rect -914 -121 -856 -109
rect -914 -1097 -902 -121
rect -868 -1097 -856 -121
rect -914 -1109 -856 -1097
rect -656 -121 -598 -109
rect -656 -1097 -644 -121
rect -610 -1097 -598 -121
rect -656 -1109 -598 -1097
rect -536 -121 -478 -109
rect -536 -1097 -524 -121
rect -490 -1097 -478 -121
rect -536 -1109 -478 -1097
rect -278 -121 -220 -109
rect -278 -1097 -266 -121
rect -232 -1097 -220 -121
rect -278 -1109 -220 -1097
rect -158 -121 -100 -109
rect -158 -1097 -146 -121
rect -112 -1097 -100 -121
rect -158 -1109 -100 -1097
rect 100 -121 158 -109
rect 100 -1097 112 -121
rect 146 -1097 158 -121
rect 100 -1109 158 -1097
rect 220 -121 278 -109
rect 220 -1097 232 -121
rect 266 -1097 278 -121
rect 220 -1109 278 -1097
rect 478 -121 536 -109
rect 478 -1097 490 -121
rect 524 -1097 536 -121
rect 478 -1109 536 -1097
rect 598 -121 656 -109
rect 598 -1097 610 -121
rect 644 -1097 656 -121
rect 598 -1109 656 -1097
rect 856 -121 914 -109
rect 856 -1097 868 -121
rect 902 -1097 914 -121
rect 856 -1109 914 -1097
rect 976 -121 1034 -109
rect 976 -1097 988 -121
rect 1022 -1097 1034 -121
rect 976 -1109 1034 -1097
rect 1234 -121 1292 -109
rect 1234 -1097 1246 -121
rect 1280 -1097 1292 -121
rect 1234 -1109 1292 -1097
rect 1354 -121 1412 -109
rect 1354 -1097 1366 -121
rect 1400 -1097 1412 -121
rect 1354 -1109 1412 -1097
rect 1612 -121 1670 -109
rect 1612 -1097 1624 -121
rect 1658 -1097 1670 -121
rect 1612 -1109 1670 -1097
rect 1732 -121 1790 -109
rect 1732 -1097 1744 -121
rect 1778 -1097 1790 -121
rect 1732 -1109 1790 -1097
rect 1990 -121 2048 -109
rect 1990 -1097 2002 -121
rect 2036 -1097 2048 -121
rect 1990 -1109 2048 -1097
rect 2110 -121 2168 -109
rect 2110 -1097 2122 -121
rect 2156 -1097 2168 -121
rect 2110 -1109 2168 -1097
rect 2368 -121 2426 -109
rect 2368 -1097 2380 -121
rect 2414 -1097 2426 -121
rect 2368 -1109 2426 -1097
rect 2488 -121 2546 -109
rect 2488 -1097 2500 -121
rect 2534 -1097 2546 -121
rect 2488 -1109 2546 -1097
rect 2746 -121 2804 -109
rect 2746 -1097 2758 -121
rect 2792 -1097 2804 -121
rect 2746 -1109 2804 -1097
rect 2866 -121 2924 -109
rect 2866 -1097 2878 -121
rect 2912 -1097 2924 -121
rect 2866 -1109 2924 -1097
rect 3124 -121 3182 -109
rect 3124 -1097 3136 -121
rect 3170 -1097 3182 -121
rect 3124 -1109 3182 -1097
rect 3244 -121 3302 -109
rect 3244 -1097 3256 -121
rect 3290 -1097 3302 -121
rect 3244 -1109 3302 -1097
rect 3502 -121 3560 -109
rect 3502 -1097 3514 -121
rect 3548 -1097 3560 -121
rect 3502 -1109 3560 -1097
rect 3622 -121 3680 -109
rect 3622 -1097 3634 -121
rect 3668 -1097 3680 -121
rect 3622 -1109 3680 -1097
rect 3880 -121 3938 -109
rect 3880 -1097 3892 -121
rect 3926 -1097 3938 -121
rect 3880 -1109 3938 -1097
rect 4000 -121 4058 -109
rect 4000 -1097 4012 -121
rect 4046 -1097 4058 -121
rect 4000 -1109 4058 -1097
rect 4258 -121 4316 -109
rect 4258 -1097 4270 -121
rect 4304 -1097 4316 -121
rect 4258 -1109 4316 -1097
rect 4378 -121 4436 -109
rect 4378 -1097 4390 -121
rect 4424 -1097 4436 -121
rect 4378 -1109 4436 -1097
rect 4636 -121 4694 -109
rect 4636 -1097 4648 -121
rect 4682 -1097 4694 -121
rect 4636 -1109 4694 -1097
rect -4694 -1339 -4636 -1327
rect -4694 -2315 -4682 -1339
rect -4648 -2315 -4636 -1339
rect -4694 -2327 -4636 -2315
rect -4436 -1339 -4378 -1327
rect -4436 -2315 -4424 -1339
rect -4390 -2315 -4378 -1339
rect -4436 -2327 -4378 -2315
rect -4316 -1339 -4258 -1327
rect -4316 -2315 -4304 -1339
rect -4270 -2315 -4258 -1339
rect -4316 -2327 -4258 -2315
rect -4058 -1339 -4000 -1327
rect -4058 -2315 -4046 -1339
rect -4012 -2315 -4000 -1339
rect -4058 -2327 -4000 -2315
rect -3938 -1339 -3880 -1327
rect -3938 -2315 -3926 -1339
rect -3892 -2315 -3880 -1339
rect -3938 -2327 -3880 -2315
rect -3680 -1339 -3622 -1327
rect -3680 -2315 -3668 -1339
rect -3634 -2315 -3622 -1339
rect -3680 -2327 -3622 -2315
rect -3560 -1339 -3502 -1327
rect -3560 -2315 -3548 -1339
rect -3514 -2315 -3502 -1339
rect -3560 -2327 -3502 -2315
rect -3302 -1339 -3244 -1327
rect -3302 -2315 -3290 -1339
rect -3256 -2315 -3244 -1339
rect -3302 -2327 -3244 -2315
rect -3182 -1339 -3124 -1327
rect -3182 -2315 -3170 -1339
rect -3136 -2315 -3124 -1339
rect -3182 -2327 -3124 -2315
rect -2924 -1339 -2866 -1327
rect -2924 -2315 -2912 -1339
rect -2878 -2315 -2866 -1339
rect -2924 -2327 -2866 -2315
rect -2804 -1339 -2746 -1327
rect -2804 -2315 -2792 -1339
rect -2758 -2315 -2746 -1339
rect -2804 -2327 -2746 -2315
rect -2546 -1339 -2488 -1327
rect -2546 -2315 -2534 -1339
rect -2500 -2315 -2488 -1339
rect -2546 -2327 -2488 -2315
rect -2426 -1339 -2368 -1327
rect -2426 -2315 -2414 -1339
rect -2380 -2315 -2368 -1339
rect -2426 -2327 -2368 -2315
rect -2168 -1339 -2110 -1327
rect -2168 -2315 -2156 -1339
rect -2122 -2315 -2110 -1339
rect -2168 -2327 -2110 -2315
rect -2048 -1339 -1990 -1327
rect -2048 -2315 -2036 -1339
rect -2002 -2315 -1990 -1339
rect -2048 -2327 -1990 -2315
rect -1790 -1339 -1732 -1327
rect -1790 -2315 -1778 -1339
rect -1744 -2315 -1732 -1339
rect -1790 -2327 -1732 -2315
rect -1670 -1339 -1612 -1327
rect -1670 -2315 -1658 -1339
rect -1624 -2315 -1612 -1339
rect -1670 -2327 -1612 -2315
rect -1412 -1339 -1354 -1327
rect -1412 -2315 -1400 -1339
rect -1366 -2315 -1354 -1339
rect -1412 -2327 -1354 -2315
rect -1292 -1339 -1234 -1327
rect -1292 -2315 -1280 -1339
rect -1246 -2315 -1234 -1339
rect -1292 -2327 -1234 -2315
rect -1034 -1339 -976 -1327
rect -1034 -2315 -1022 -1339
rect -988 -2315 -976 -1339
rect -1034 -2327 -976 -2315
rect -914 -1339 -856 -1327
rect -914 -2315 -902 -1339
rect -868 -2315 -856 -1339
rect -914 -2327 -856 -2315
rect -656 -1339 -598 -1327
rect -656 -2315 -644 -1339
rect -610 -2315 -598 -1339
rect -656 -2327 -598 -2315
rect -536 -1339 -478 -1327
rect -536 -2315 -524 -1339
rect -490 -2315 -478 -1339
rect -536 -2327 -478 -2315
rect -278 -1339 -220 -1327
rect -278 -2315 -266 -1339
rect -232 -2315 -220 -1339
rect -278 -2327 -220 -2315
rect -158 -1339 -100 -1327
rect -158 -2315 -146 -1339
rect -112 -2315 -100 -1339
rect -158 -2327 -100 -2315
rect 100 -1339 158 -1327
rect 100 -2315 112 -1339
rect 146 -2315 158 -1339
rect 100 -2327 158 -2315
rect 220 -1339 278 -1327
rect 220 -2315 232 -1339
rect 266 -2315 278 -1339
rect 220 -2327 278 -2315
rect 478 -1339 536 -1327
rect 478 -2315 490 -1339
rect 524 -2315 536 -1339
rect 478 -2327 536 -2315
rect 598 -1339 656 -1327
rect 598 -2315 610 -1339
rect 644 -2315 656 -1339
rect 598 -2327 656 -2315
rect 856 -1339 914 -1327
rect 856 -2315 868 -1339
rect 902 -2315 914 -1339
rect 856 -2327 914 -2315
rect 976 -1339 1034 -1327
rect 976 -2315 988 -1339
rect 1022 -2315 1034 -1339
rect 976 -2327 1034 -2315
rect 1234 -1339 1292 -1327
rect 1234 -2315 1246 -1339
rect 1280 -2315 1292 -1339
rect 1234 -2327 1292 -2315
rect 1354 -1339 1412 -1327
rect 1354 -2315 1366 -1339
rect 1400 -2315 1412 -1339
rect 1354 -2327 1412 -2315
rect 1612 -1339 1670 -1327
rect 1612 -2315 1624 -1339
rect 1658 -2315 1670 -1339
rect 1612 -2327 1670 -2315
rect 1732 -1339 1790 -1327
rect 1732 -2315 1744 -1339
rect 1778 -2315 1790 -1339
rect 1732 -2327 1790 -2315
rect 1990 -1339 2048 -1327
rect 1990 -2315 2002 -1339
rect 2036 -2315 2048 -1339
rect 1990 -2327 2048 -2315
rect 2110 -1339 2168 -1327
rect 2110 -2315 2122 -1339
rect 2156 -2315 2168 -1339
rect 2110 -2327 2168 -2315
rect 2368 -1339 2426 -1327
rect 2368 -2315 2380 -1339
rect 2414 -2315 2426 -1339
rect 2368 -2327 2426 -2315
rect 2488 -1339 2546 -1327
rect 2488 -2315 2500 -1339
rect 2534 -2315 2546 -1339
rect 2488 -2327 2546 -2315
rect 2746 -1339 2804 -1327
rect 2746 -2315 2758 -1339
rect 2792 -2315 2804 -1339
rect 2746 -2327 2804 -2315
rect 2866 -1339 2924 -1327
rect 2866 -2315 2878 -1339
rect 2912 -2315 2924 -1339
rect 2866 -2327 2924 -2315
rect 3124 -1339 3182 -1327
rect 3124 -2315 3136 -1339
rect 3170 -2315 3182 -1339
rect 3124 -2327 3182 -2315
rect 3244 -1339 3302 -1327
rect 3244 -2315 3256 -1339
rect 3290 -2315 3302 -1339
rect 3244 -2327 3302 -2315
rect 3502 -1339 3560 -1327
rect 3502 -2315 3514 -1339
rect 3548 -2315 3560 -1339
rect 3502 -2327 3560 -2315
rect 3622 -1339 3680 -1327
rect 3622 -2315 3634 -1339
rect 3668 -2315 3680 -1339
rect 3622 -2327 3680 -2315
rect 3880 -1339 3938 -1327
rect 3880 -2315 3892 -1339
rect 3926 -2315 3938 -1339
rect 3880 -2327 3938 -2315
rect 4000 -1339 4058 -1327
rect 4000 -2315 4012 -1339
rect 4046 -2315 4058 -1339
rect 4000 -2327 4058 -2315
rect 4258 -1339 4316 -1327
rect 4258 -2315 4270 -1339
rect 4304 -2315 4316 -1339
rect 4258 -2327 4316 -2315
rect 4378 -1339 4436 -1327
rect 4378 -2315 4390 -1339
rect 4424 -2315 4436 -1339
rect 4378 -2327 4436 -2315
rect 4636 -1339 4694 -1327
rect 4636 -2315 4648 -1339
rect 4682 -2315 4694 -1339
rect 4636 -2327 4694 -2315
<< mvndiffc >>
rect -4682 1339 -4648 2315
rect -4424 1339 -4390 2315
rect -4304 1339 -4270 2315
rect -4046 1339 -4012 2315
rect -3926 1339 -3892 2315
rect -3668 1339 -3634 2315
rect -3548 1339 -3514 2315
rect -3290 1339 -3256 2315
rect -3170 1339 -3136 2315
rect -2912 1339 -2878 2315
rect -2792 1339 -2758 2315
rect -2534 1339 -2500 2315
rect -2414 1339 -2380 2315
rect -2156 1339 -2122 2315
rect -2036 1339 -2002 2315
rect -1778 1339 -1744 2315
rect -1658 1339 -1624 2315
rect -1400 1339 -1366 2315
rect -1280 1339 -1246 2315
rect -1022 1339 -988 2315
rect -902 1339 -868 2315
rect -644 1339 -610 2315
rect -524 1339 -490 2315
rect -266 1339 -232 2315
rect -146 1339 -112 2315
rect 112 1339 146 2315
rect 232 1339 266 2315
rect 490 1339 524 2315
rect 610 1339 644 2315
rect 868 1339 902 2315
rect 988 1339 1022 2315
rect 1246 1339 1280 2315
rect 1366 1339 1400 2315
rect 1624 1339 1658 2315
rect 1744 1339 1778 2315
rect 2002 1339 2036 2315
rect 2122 1339 2156 2315
rect 2380 1339 2414 2315
rect 2500 1339 2534 2315
rect 2758 1339 2792 2315
rect 2878 1339 2912 2315
rect 3136 1339 3170 2315
rect 3256 1339 3290 2315
rect 3514 1339 3548 2315
rect 3634 1339 3668 2315
rect 3892 1339 3926 2315
rect 4012 1339 4046 2315
rect 4270 1339 4304 2315
rect 4390 1339 4424 2315
rect 4648 1339 4682 2315
rect -4682 121 -4648 1097
rect -4424 121 -4390 1097
rect -4304 121 -4270 1097
rect -4046 121 -4012 1097
rect -3926 121 -3892 1097
rect -3668 121 -3634 1097
rect -3548 121 -3514 1097
rect -3290 121 -3256 1097
rect -3170 121 -3136 1097
rect -2912 121 -2878 1097
rect -2792 121 -2758 1097
rect -2534 121 -2500 1097
rect -2414 121 -2380 1097
rect -2156 121 -2122 1097
rect -2036 121 -2002 1097
rect -1778 121 -1744 1097
rect -1658 121 -1624 1097
rect -1400 121 -1366 1097
rect -1280 121 -1246 1097
rect -1022 121 -988 1097
rect -902 121 -868 1097
rect -644 121 -610 1097
rect -524 121 -490 1097
rect -266 121 -232 1097
rect -146 121 -112 1097
rect 112 121 146 1097
rect 232 121 266 1097
rect 490 121 524 1097
rect 610 121 644 1097
rect 868 121 902 1097
rect 988 121 1022 1097
rect 1246 121 1280 1097
rect 1366 121 1400 1097
rect 1624 121 1658 1097
rect 1744 121 1778 1097
rect 2002 121 2036 1097
rect 2122 121 2156 1097
rect 2380 121 2414 1097
rect 2500 121 2534 1097
rect 2758 121 2792 1097
rect 2878 121 2912 1097
rect 3136 121 3170 1097
rect 3256 121 3290 1097
rect 3514 121 3548 1097
rect 3634 121 3668 1097
rect 3892 121 3926 1097
rect 4012 121 4046 1097
rect 4270 121 4304 1097
rect 4390 121 4424 1097
rect 4648 121 4682 1097
rect -4682 -1097 -4648 -121
rect -4424 -1097 -4390 -121
rect -4304 -1097 -4270 -121
rect -4046 -1097 -4012 -121
rect -3926 -1097 -3892 -121
rect -3668 -1097 -3634 -121
rect -3548 -1097 -3514 -121
rect -3290 -1097 -3256 -121
rect -3170 -1097 -3136 -121
rect -2912 -1097 -2878 -121
rect -2792 -1097 -2758 -121
rect -2534 -1097 -2500 -121
rect -2414 -1097 -2380 -121
rect -2156 -1097 -2122 -121
rect -2036 -1097 -2002 -121
rect -1778 -1097 -1744 -121
rect -1658 -1097 -1624 -121
rect -1400 -1097 -1366 -121
rect -1280 -1097 -1246 -121
rect -1022 -1097 -988 -121
rect -902 -1097 -868 -121
rect -644 -1097 -610 -121
rect -524 -1097 -490 -121
rect -266 -1097 -232 -121
rect -146 -1097 -112 -121
rect 112 -1097 146 -121
rect 232 -1097 266 -121
rect 490 -1097 524 -121
rect 610 -1097 644 -121
rect 868 -1097 902 -121
rect 988 -1097 1022 -121
rect 1246 -1097 1280 -121
rect 1366 -1097 1400 -121
rect 1624 -1097 1658 -121
rect 1744 -1097 1778 -121
rect 2002 -1097 2036 -121
rect 2122 -1097 2156 -121
rect 2380 -1097 2414 -121
rect 2500 -1097 2534 -121
rect 2758 -1097 2792 -121
rect 2878 -1097 2912 -121
rect 3136 -1097 3170 -121
rect 3256 -1097 3290 -121
rect 3514 -1097 3548 -121
rect 3634 -1097 3668 -121
rect 3892 -1097 3926 -121
rect 4012 -1097 4046 -121
rect 4270 -1097 4304 -121
rect 4390 -1097 4424 -121
rect 4648 -1097 4682 -121
rect -4682 -2315 -4648 -1339
rect -4424 -2315 -4390 -1339
rect -4304 -2315 -4270 -1339
rect -4046 -2315 -4012 -1339
rect -3926 -2315 -3892 -1339
rect -3668 -2315 -3634 -1339
rect -3548 -2315 -3514 -1339
rect -3290 -2315 -3256 -1339
rect -3170 -2315 -3136 -1339
rect -2912 -2315 -2878 -1339
rect -2792 -2315 -2758 -1339
rect -2534 -2315 -2500 -1339
rect -2414 -2315 -2380 -1339
rect -2156 -2315 -2122 -1339
rect -2036 -2315 -2002 -1339
rect -1778 -2315 -1744 -1339
rect -1658 -2315 -1624 -1339
rect -1400 -2315 -1366 -1339
rect -1280 -2315 -1246 -1339
rect -1022 -2315 -988 -1339
rect -902 -2315 -868 -1339
rect -644 -2315 -610 -1339
rect -524 -2315 -490 -1339
rect -266 -2315 -232 -1339
rect -146 -2315 -112 -1339
rect 112 -2315 146 -1339
rect 232 -2315 266 -1339
rect 490 -2315 524 -1339
rect 610 -2315 644 -1339
rect 868 -2315 902 -1339
rect 988 -2315 1022 -1339
rect 1246 -2315 1280 -1339
rect 1366 -2315 1400 -1339
rect 1624 -2315 1658 -1339
rect 1744 -2315 1778 -1339
rect 2002 -2315 2036 -1339
rect 2122 -2315 2156 -1339
rect 2380 -2315 2414 -1339
rect 2500 -2315 2534 -1339
rect 2758 -2315 2792 -1339
rect 2878 -2315 2912 -1339
rect 3136 -2315 3170 -1339
rect 3256 -2315 3290 -1339
rect 3514 -2315 3548 -1339
rect 3634 -2315 3668 -1339
rect 3892 -2315 3926 -1339
rect 4012 -2315 4046 -1339
rect 4270 -2315 4304 -1339
rect 4390 -2315 4424 -1339
rect 4648 -2315 4682 -1339
<< mvpsubdiff >>
rect -4828 2537 4828 2549
rect -4828 2503 -4720 2537
rect 4720 2503 4828 2537
rect -4828 2491 4828 2503
rect -4828 2441 -4770 2491
rect -4828 -2441 -4816 2441
rect -4782 -2441 -4770 2441
rect 4770 2441 4828 2491
rect -4828 -2491 -4770 -2441
rect 4770 -2441 4782 2441
rect 4816 -2441 4828 2441
rect 4770 -2491 4828 -2441
rect -4828 -2503 4828 -2491
rect -4828 -2537 -4720 -2503
rect 4720 -2537 4828 -2503
rect -4828 -2549 4828 -2537
<< mvpsubdiffcont >>
rect -4720 2503 4720 2537
rect -4816 -2441 -4782 2441
rect 4782 -2441 4816 2441
rect -4720 -2537 4720 -2503
<< poly >>
rect -4636 2399 -4436 2415
rect -4636 2365 -4620 2399
rect -4452 2365 -4436 2399
rect -4636 2327 -4436 2365
rect -4258 2399 -4058 2415
rect -4258 2365 -4242 2399
rect -4074 2365 -4058 2399
rect -4258 2327 -4058 2365
rect -3880 2399 -3680 2415
rect -3880 2365 -3864 2399
rect -3696 2365 -3680 2399
rect -3880 2327 -3680 2365
rect -3502 2399 -3302 2415
rect -3502 2365 -3486 2399
rect -3318 2365 -3302 2399
rect -3502 2327 -3302 2365
rect -3124 2399 -2924 2415
rect -3124 2365 -3108 2399
rect -2940 2365 -2924 2399
rect -3124 2327 -2924 2365
rect -2746 2399 -2546 2415
rect -2746 2365 -2730 2399
rect -2562 2365 -2546 2399
rect -2746 2327 -2546 2365
rect -2368 2399 -2168 2415
rect -2368 2365 -2352 2399
rect -2184 2365 -2168 2399
rect -2368 2327 -2168 2365
rect -1990 2399 -1790 2415
rect -1990 2365 -1974 2399
rect -1806 2365 -1790 2399
rect -1990 2327 -1790 2365
rect -1612 2399 -1412 2415
rect -1612 2365 -1596 2399
rect -1428 2365 -1412 2399
rect -1612 2327 -1412 2365
rect -1234 2399 -1034 2415
rect -1234 2365 -1218 2399
rect -1050 2365 -1034 2399
rect -1234 2327 -1034 2365
rect -856 2399 -656 2415
rect -856 2365 -840 2399
rect -672 2365 -656 2399
rect -856 2327 -656 2365
rect -478 2399 -278 2415
rect -478 2365 -462 2399
rect -294 2365 -278 2399
rect -478 2327 -278 2365
rect -100 2399 100 2415
rect -100 2365 -84 2399
rect 84 2365 100 2399
rect -100 2327 100 2365
rect 278 2399 478 2415
rect 278 2365 294 2399
rect 462 2365 478 2399
rect 278 2327 478 2365
rect 656 2399 856 2415
rect 656 2365 672 2399
rect 840 2365 856 2399
rect 656 2327 856 2365
rect 1034 2399 1234 2415
rect 1034 2365 1050 2399
rect 1218 2365 1234 2399
rect 1034 2327 1234 2365
rect 1412 2399 1612 2415
rect 1412 2365 1428 2399
rect 1596 2365 1612 2399
rect 1412 2327 1612 2365
rect 1790 2399 1990 2415
rect 1790 2365 1806 2399
rect 1974 2365 1990 2399
rect 1790 2327 1990 2365
rect 2168 2399 2368 2415
rect 2168 2365 2184 2399
rect 2352 2365 2368 2399
rect 2168 2327 2368 2365
rect 2546 2399 2746 2415
rect 2546 2365 2562 2399
rect 2730 2365 2746 2399
rect 2546 2327 2746 2365
rect 2924 2399 3124 2415
rect 2924 2365 2940 2399
rect 3108 2365 3124 2399
rect 2924 2327 3124 2365
rect 3302 2399 3502 2415
rect 3302 2365 3318 2399
rect 3486 2365 3502 2399
rect 3302 2327 3502 2365
rect 3680 2399 3880 2415
rect 3680 2365 3696 2399
rect 3864 2365 3880 2399
rect 3680 2327 3880 2365
rect 4058 2399 4258 2415
rect 4058 2365 4074 2399
rect 4242 2365 4258 2399
rect 4058 2327 4258 2365
rect 4436 2399 4636 2415
rect 4436 2365 4452 2399
rect 4620 2365 4636 2399
rect 4436 2327 4636 2365
rect -4636 1289 -4436 1327
rect -4636 1255 -4620 1289
rect -4452 1255 -4436 1289
rect -4636 1239 -4436 1255
rect -4258 1289 -4058 1327
rect -4258 1255 -4242 1289
rect -4074 1255 -4058 1289
rect -4258 1239 -4058 1255
rect -3880 1289 -3680 1327
rect -3880 1255 -3864 1289
rect -3696 1255 -3680 1289
rect -3880 1239 -3680 1255
rect -3502 1289 -3302 1327
rect -3502 1255 -3486 1289
rect -3318 1255 -3302 1289
rect -3502 1239 -3302 1255
rect -3124 1289 -2924 1327
rect -3124 1255 -3108 1289
rect -2940 1255 -2924 1289
rect -3124 1239 -2924 1255
rect -2746 1289 -2546 1327
rect -2746 1255 -2730 1289
rect -2562 1255 -2546 1289
rect -2746 1239 -2546 1255
rect -2368 1289 -2168 1327
rect -2368 1255 -2352 1289
rect -2184 1255 -2168 1289
rect -2368 1239 -2168 1255
rect -1990 1289 -1790 1327
rect -1990 1255 -1974 1289
rect -1806 1255 -1790 1289
rect -1990 1239 -1790 1255
rect -1612 1289 -1412 1327
rect -1612 1255 -1596 1289
rect -1428 1255 -1412 1289
rect -1612 1239 -1412 1255
rect -1234 1289 -1034 1327
rect -1234 1255 -1218 1289
rect -1050 1255 -1034 1289
rect -1234 1239 -1034 1255
rect -856 1289 -656 1327
rect -856 1255 -840 1289
rect -672 1255 -656 1289
rect -856 1239 -656 1255
rect -478 1289 -278 1327
rect -478 1255 -462 1289
rect -294 1255 -278 1289
rect -478 1239 -278 1255
rect -100 1289 100 1327
rect -100 1255 -84 1289
rect 84 1255 100 1289
rect -100 1239 100 1255
rect 278 1289 478 1327
rect 278 1255 294 1289
rect 462 1255 478 1289
rect 278 1239 478 1255
rect 656 1289 856 1327
rect 656 1255 672 1289
rect 840 1255 856 1289
rect 656 1239 856 1255
rect 1034 1289 1234 1327
rect 1034 1255 1050 1289
rect 1218 1255 1234 1289
rect 1034 1239 1234 1255
rect 1412 1289 1612 1327
rect 1412 1255 1428 1289
rect 1596 1255 1612 1289
rect 1412 1239 1612 1255
rect 1790 1289 1990 1327
rect 1790 1255 1806 1289
rect 1974 1255 1990 1289
rect 1790 1239 1990 1255
rect 2168 1289 2368 1327
rect 2168 1255 2184 1289
rect 2352 1255 2368 1289
rect 2168 1239 2368 1255
rect 2546 1289 2746 1327
rect 2546 1255 2562 1289
rect 2730 1255 2746 1289
rect 2546 1239 2746 1255
rect 2924 1289 3124 1327
rect 2924 1255 2940 1289
rect 3108 1255 3124 1289
rect 2924 1239 3124 1255
rect 3302 1289 3502 1327
rect 3302 1255 3318 1289
rect 3486 1255 3502 1289
rect 3302 1239 3502 1255
rect 3680 1289 3880 1327
rect 3680 1255 3696 1289
rect 3864 1255 3880 1289
rect 3680 1239 3880 1255
rect 4058 1289 4258 1327
rect 4058 1255 4074 1289
rect 4242 1255 4258 1289
rect 4058 1239 4258 1255
rect 4436 1289 4636 1327
rect 4436 1255 4452 1289
rect 4620 1255 4636 1289
rect 4436 1239 4636 1255
rect -4636 1181 -4436 1197
rect -4636 1147 -4620 1181
rect -4452 1147 -4436 1181
rect -4636 1109 -4436 1147
rect -4258 1181 -4058 1197
rect -4258 1147 -4242 1181
rect -4074 1147 -4058 1181
rect -4258 1109 -4058 1147
rect -3880 1181 -3680 1197
rect -3880 1147 -3864 1181
rect -3696 1147 -3680 1181
rect -3880 1109 -3680 1147
rect -3502 1181 -3302 1197
rect -3502 1147 -3486 1181
rect -3318 1147 -3302 1181
rect -3502 1109 -3302 1147
rect -3124 1181 -2924 1197
rect -3124 1147 -3108 1181
rect -2940 1147 -2924 1181
rect -3124 1109 -2924 1147
rect -2746 1181 -2546 1197
rect -2746 1147 -2730 1181
rect -2562 1147 -2546 1181
rect -2746 1109 -2546 1147
rect -2368 1181 -2168 1197
rect -2368 1147 -2352 1181
rect -2184 1147 -2168 1181
rect -2368 1109 -2168 1147
rect -1990 1181 -1790 1197
rect -1990 1147 -1974 1181
rect -1806 1147 -1790 1181
rect -1990 1109 -1790 1147
rect -1612 1181 -1412 1197
rect -1612 1147 -1596 1181
rect -1428 1147 -1412 1181
rect -1612 1109 -1412 1147
rect -1234 1181 -1034 1197
rect -1234 1147 -1218 1181
rect -1050 1147 -1034 1181
rect -1234 1109 -1034 1147
rect -856 1181 -656 1197
rect -856 1147 -840 1181
rect -672 1147 -656 1181
rect -856 1109 -656 1147
rect -478 1181 -278 1197
rect -478 1147 -462 1181
rect -294 1147 -278 1181
rect -478 1109 -278 1147
rect -100 1181 100 1197
rect -100 1147 -84 1181
rect 84 1147 100 1181
rect -100 1109 100 1147
rect 278 1181 478 1197
rect 278 1147 294 1181
rect 462 1147 478 1181
rect 278 1109 478 1147
rect 656 1181 856 1197
rect 656 1147 672 1181
rect 840 1147 856 1181
rect 656 1109 856 1147
rect 1034 1181 1234 1197
rect 1034 1147 1050 1181
rect 1218 1147 1234 1181
rect 1034 1109 1234 1147
rect 1412 1181 1612 1197
rect 1412 1147 1428 1181
rect 1596 1147 1612 1181
rect 1412 1109 1612 1147
rect 1790 1181 1990 1197
rect 1790 1147 1806 1181
rect 1974 1147 1990 1181
rect 1790 1109 1990 1147
rect 2168 1181 2368 1197
rect 2168 1147 2184 1181
rect 2352 1147 2368 1181
rect 2168 1109 2368 1147
rect 2546 1181 2746 1197
rect 2546 1147 2562 1181
rect 2730 1147 2746 1181
rect 2546 1109 2746 1147
rect 2924 1181 3124 1197
rect 2924 1147 2940 1181
rect 3108 1147 3124 1181
rect 2924 1109 3124 1147
rect 3302 1181 3502 1197
rect 3302 1147 3318 1181
rect 3486 1147 3502 1181
rect 3302 1109 3502 1147
rect 3680 1181 3880 1197
rect 3680 1147 3696 1181
rect 3864 1147 3880 1181
rect 3680 1109 3880 1147
rect 4058 1181 4258 1197
rect 4058 1147 4074 1181
rect 4242 1147 4258 1181
rect 4058 1109 4258 1147
rect 4436 1181 4636 1197
rect 4436 1147 4452 1181
rect 4620 1147 4636 1181
rect 4436 1109 4636 1147
rect -4636 71 -4436 109
rect -4636 37 -4620 71
rect -4452 37 -4436 71
rect -4636 21 -4436 37
rect -4258 71 -4058 109
rect -4258 37 -4242 71
rect -4074 37 -4058 71
rect -4258 21 -4058 37
rect -3880 71 -3680 109
rect -3880 37 -3864 71
rect -3696 37 -3680 71
rect -3880 21 -3680 37
rect -3502 71 -3302 109
rect -3502 37 -3486 71
rect -3318 37 -3302 71
rect -3502 21 -3302 37
rect -3124 71 -2924 109
rect -3124 37 -3108 71
rect -2940 37 -2924 71
rect -3124 21 -2924 37
rect -2746 71 -2546 109
rect -2746 37 -2730 71
rect -2562 37 -2546 71
rect -2746 21 -2546 37
rect -2368 71 -2168 109
rect -2368 37 -2352 71
rect -2184 37 -2168 71
rect -2368 21 -2168 37
rect -1990 71 -1790 109
rect -1990 37 -1974 71
rect -1806 37 -1790 71
rect -1990 21 -1790 37
rect -1612 71 -1412 109
rect -1612 37 -1596 71
rect -1428 37 -1412 71
rect -1612 21 -1412 37
rect -1234 71 -1034 109
rect -1234 37 -1218 71
rect -1050 37 -1034 71
rect -1234 21 -1034 37
rect -856 71 -656 109
rect -856 37 -840 71
rect -672 37 -656 71
rect -856 21 -656 37
rect -478 71 -278 109
rect -478 37 -462 71
rect -294 37 -278 71
rect -478 21 -278 37
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect 278 71 478 109
rect 278 37 294 71
rect 462 37 478 71
rect 278 21 478 37
rect 656 71 856 109
rect 656 37 672 71
rect 840 37 856 71
rect 656 21 856 37
rect 1034 71 1234 109
rect 1034 37 1050 71
rect 1218 37 1234 71
rect 1034 21 1234 37
rect 1412 71 1612 109
rect 1412 37 1428 71
rect 1596 37 1612 71
rect 1412 21 1612 37
rect 1790 71 1990 109
rect 1790 37 1806 71
rect 1974 37 1990 71
rect 1790 21 1990 37
rect 2168 71 2368 109
rect 2168 37 2184 71
rect 2352 37 2368 71
rect 2168 21 2368 37
rect 2546 71 2746 109
rect 2546 37 2562 71
rect 2730 37 2746 71
rect 2546 21 2746 37
rect 2924 71 3124 109
rect 2924 37 2940 71
rect 3108 37 3124 71
rect 2924 21 3124 37
rect 3302 71 3502 109
rect 3302 37 3318 71
rect 3486 37 3502 71
rect 3302 21 3502 37
rect 3680 71 3880 109
rect 3680 37 3696 71
rect 3864 37 3880 71
rect 3680 21 3880 37
rect 4058 71 4258 109
rect 4058 37 4074 71
rect 4242 37 4258 71
rect 4058 21 4258 37
rect 4436 71 4636 109
rect 4436 37 4452 71
rect 4620 37 4636 71
rect 4436 21 4636 37
rect -4636 -37 -4436 -21
rect -4636 -71 -4620 -37
rect -4452 -71 -4436 -37
rect -4636 -109 -4436 -71
rect -4258 -37 -4058 -21
rect -4258 -71 -4242 -37
rect -4074 -71 -4058 -37
rect -4258 -109 -4058 -71
rect -3880 -37 -3680 -21
rect -3880 -71 -3864 -37
rect -3696 -71 -3680 -37
rect -3880 -109 -3680 -71
rect -3502 -37 -3302 -21
rect -3502 -71 -3486 -37
rect -3318 -71 -3302 -37
rect -3502 -109 -3302 -71
rect -3124 -37 -2924 -21
rect -3124 -71 -3108 -37
rect -2940 -71 -2924 -37
rect -3124 -109 -2924 -71
rect -2746 -37 -2546 -21
rect -2746 -71 -2730 -37
rect -2562 -71 -2546 -37
rect -2746 -109 -2546 -71
rect -2368 -37 -2168 -21
rect -2368 -71 -2352 -37
rect -2184 -71 -2168 -37
rect -2368 -109 -2168 -71
rect -1990 -37 -1790 -21
rect -1990 -71 -1974 -37
rect -1806 -71 -1790 -37
rect -1990 -109 -1790 -71
rect -1612 -37 -1412 -21
rect -1612 -71 -1596 -37
rect -1428 -71 -1412 -37
rect -1612 -109 -1412 -71
rect -1234 -37 -1034 -21
rect -1234 -71 -1218 -37
rect -1050 -71 -1034 -37
rect -1234 -109 -1034 -71
rect -856 -37 -656 -21
rect -856 -71 -840 -37
rect -672 -71 -656 -37
rect -856 -109 -656 -71
rect -478 -37 -278 -21
rect -478 -71 -462 -37
rect -294 -71 -278 -37
rect -478 -109 -278 -71
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect 278 -37 478 -21
rect 278 -71 294 -37
rect 462 -71 478 -37
rect 278 -109 478 -71
rect 656 -37 856 -21
rect 656 -71 672 -37
rect 840 -71 856 -37
rect 656 -109 856 -71
rect 1034 -37 1234 -21
rect 1034 -71 1050 -37
rect 1218 -71 1234 -37
rect 1034 -109 1234 -71
rect 1412 -37 1612 -21
rect 1412 -71 1428 -37
rect 1596 -71 1612 -37
rect 1412 -109 1612 -71
rect 1790 -37 1990 -21
rect 1790 -71 1806 -37
rect 1974 -71 1990 -37
rect 1790 -109 1990 -71
rect 2168 -37 2368 -21
rect 2168 -71 2184 -37
rect 2352 -71 2368 -37
rect 2168 -109 2368 -71
rect 2546 -37 2746 -21
rect 2546 -71 2562 -37
rect 2730 -71 2746 -37
rect 2546 -109 2746 -71
rect 2924 -37 3124 -21
rect 2924 -71 2940 -37
rect 3108 -71 3124 -37
rect 2924 -109 3124 -71
rect 3302 -37 3502 -21
rect 3302 -71 3318 -37
rect 3486 -71 3502 -37
rect 3302 -109 3502 -71
rect 3680 -37 3880 -21
rect 3680 -71 3696 -37
rect 3864 -71 3880 -37
rect 3680 -109 3880 -71
rect 4058 -37 4258 -21
rect 4058 -71 4074 -37
rect 4242 -71 4258 -37
rect 4058 -109 4258 -71
rect 4436 -37 4636 -21
rect 4436 -71 4452 -37
rect 4620 -71 4636 -37
rect 4436 -109 4636 -71
rect -4636 -1147 -4436 -1109
rect -4636 -1181 -4620 -1147
rect -4452 -1181 -4436 -1147
rect -4636 -1197 -4436 -1181
rect -4258 -1147 -4058 -1109
rect -4258 -1181 -4242 -1147
rect -4074 -1181 -4058 -1147
rect -4258 -1197 -4058 -1181
rect -3880 -1147 -3680 -1109
rect -3880 -1181 -3864 -1147
rect -3696 -1181 -3680 -1147
rect -3880 -1197 -3680 -1181
rect -3502 -1147 -3302 -1109
rect -3502 -1181 -3486 -1147
rect -3318 -1181 -3302 -1147
rect -3502 -1197 -3302 -1181
rect -3124 -1147 -2924 -1109
rect -3124 -1181 -3108 -1147
rect -2940 -1181 -2924 -1147
rect -3124 -1197 -2924 -1181
rect -2746 -1147 -2546 -1109
rect -2746 -1181 -2730 -1147
rect -2562 -1181 -2546 -1147
rect -2746 -1197 -2546 -1181
rect -2368 -1147 -2168 -1109
rect -2368 -1181 -2352 -1147
rect -2184 -1181 -2168 -1147
rect -2368 -1197 -2168 -1181
rect -1990 -1147 -1790 -1109
rect -1990 -1181 -1974 -1147
rect -1806 -1181 -1790 -1147
rect -1990 -1197 -1790 -1181
rect -1612 -1147 -1412 -1109
rect -1612 -1181 -1596 -1147
rect -1428 -1181 -1412 -1147
rect -1612 -1197 -1412 -1181
rect -1234 -1147 -1034 -1109
rect -1234 -1181 -1218 -1147
rect -1050 -1181 -1034 -1147
rect -1234 -1197 -1034 -1181
rect -856 -1147 -656 -1109
rect -856 -1181 -840 -1147
rect -672 -1181 -656 -1147
rect -856 -1197 -656 -1181
rect -478 -1147 -278 -1109
rect -478 -1181 -462 -1147
rect -294 -1181 -278 -1147
rect -478 -1197 -278 -1181
rect -100 -1147 100 -1109
rect -100 -1181 -84 -1147
rect 84 -1181 100 -1147
rect -100 -1197 100 -1181
rect 278 -1147 478 -1109
rect 278 -1181 294 -1147
rect 462 -1181 478 -1147
rect 278 -1197 478 -1181
rect 656 -1147 856 -1109
rect 656 -1181 672 -1147
rect 840 -1181 856 -1147
rect 656 -1197 856 -1181
rect 1034 -1147 1234 -1109
rect 1034 -1181 1050 -1147
rect 1218 -1181 1234 -1147
rect 1034 -1197 1234 -1181
rect 1412 -1147 1612 -1109
rect 1412 -1181 1428 -1147
rect 1596 -1181 1612 -1147
rect 1412 -1197 1612 -1181
rect 1790 -1147 1990 -1109
rect 1790 -1181 1806 -1147
rect 1974 -1181 1990 -1147
rect 1790 -1197 1990 -1181
rect 2168 -1147 2368 -1109
rect 2168 -1181 2184 -1147
rect 2352 -1181 2368 -1147
rect 2168 -1197 2368 -1181
rect 2546 -1147 2746 -1109
rect 2546 -1181 2562 -1147
rect 2730 -1181 2746 -1147
rect 2546 -1197 2746 -1181
rect 2924 -1147 3124 -1109
rect 2924 -1181 2940 -1147
rect 3108 -1181 3124 -1147
rect 2924 -1197 3124 -1181
rect 3302 -1147 3502 -1109
rect 3302 -1181 3318 -1147
rect 3486 -1181 3502 -1147
rect 3302 -1197 3502 -1181
rect 3680 -1147 3880 -1109
rect 3680 -1181 3696 -1147
rect 3864 -1181 3880 -1147
rect 3680 -1197 3880 -1181
rect 4058 -1147 4258 -1109
rect 4058 -1181 4074 -1147
rect 4242 -1181 4258 -1147
rect 4058 -1197 4258 -1181
rect 4436 -1147 4636 -1109
rect 4436 -1181 4452 -1147
rect 4620 -1181 4636 -1147
rect 4436 -1197 4636 -1181
rect -4636 -1255 -4436 -1239
rect -4636 -1289 -4620 -1255
rect -4452 -1289 -4436 -1255
rect -4636 -1327 -4436 -1289
rect -4258 -1255 -4058 -1239
rect -4258 -1289 -4242 -1255
rect -4074 -1289 -4058 -1255
rect -4258 -1327 -4058 -1289
rect -3880 -1255 -3680 -1239
rect -3880 -1289 -3864 -1255
rect -3696 -1289 -3680 -1255
rect -3880 -1327 -3680 -1289
rect -3502 -1255 -3302 -1239
rect -3502 -1289 -3486 -1255
rect -3318 -1289 -3302 -1255
rect -3502 -1327 -3302 -1289
rect -3124 -1255 -2924 -1239
rect -3124 -1289 -3108 -1255
rect -2940 -1289 -2924 -1255
rect -3124 -1327 -2924 -1289
rect -2746 -1255 -2546 -1239
rect -2746 -1289 -2730 -1255
rect -2562 -1289 -2546 -1255
rect -2746 -1327 -2546 -1289
rect -2368 -1255 -2168 -1239
rect -2368 -1289 -2352 -1255
rect -2184 -1289 -2168 -1255
rect -2368 -1327 -2168 -1289
rect -1990 -1255 -1790 -1239
rect -1990 -1289 -1974 -1255
rect -1806 -1289 -1790 -1255
rect -1990 -1327 -1790 -1289
rect -1612 -1255 -1412 -1239
rect -1612 -1289 -1596 -1255
rect -1428 -1289 -1412 -1255
rect -1612 -1327 -1412 -1289
rect -1234 -1255 -1034 -1239
rect -1234 -1289 -1218 -1255
rect -1050 -1289 -1034 -1255
rect -1234 -1327 -1034 -1289
rect -856 -1255 -656 -1239
rect -856 -1289 -840 -1255
rect -672 -1289 -656 -1255
rect -856 -1327 -656 -1289
rect -478 -1255 -278 -1239
rect -478 -1289 -462 -1255
rect -294 -1289 -278 -1255
rect -478 -1327 -278 -1289
rect -100 -1255 100 -1239
rect -100 -1289 -84 -1255
rect 84 -1289 100 -1255
rect -100 -1327 100 -1289
rect 278 -1255 478 -1239
rect 278 -1289 294 -1255
rect 462 -1289 478 -1255
rect 278 -1327 478 -1289
rect 656 -1255 856 -1239
rect 656 -1289 672 -1255
rect 840 -1289 856 -1255
rect 656 -1327 856 -1289
rect 1034 -1255 1234 -1239
rect 1034 -1289 1050 -1255
rect 1218 -1289 1234 -1255
rect 1034 -1327 1234 -1289
rect 1412 -1255 1612 -1239
rect 1412 -1289 1428 -1255
rect 1596 -1289 1612 -1255
rect 1412 -1327 1612 -1289
rect 1790 -1255 1990 -1239
rect 1790 -1289 1806 -1255
rect 1974 -1289 1990 -1255
rect 1790 -1327 1990 -1289
rect 2168 -1255 2368 -1239
rect 2168 -1289 2184 -1255
rect 2352 -1289 2368 -1255
rect 2168 -1327 2368 -1289
rect 2546 -1255 2746 -1239
rect 2546 -1289 2562 -1255
rect 2730 -1289 2746 -1255
rect 2546 -1327 2746 -1289
rect 2924 -1255 3124 -1239
rect 2924 -1289 2940 -1255
rect 3108 -1289 3124 -1255
rect 2924 -1327 3124 -1289
rect 3302 -1255 3502 -1239
rect 3302 -1289 3318 -1255
rect 3486 -1289 3502 -1255
rect 3302 -1327 3502 -1289
rect 3680 -1255 3880 -1239
rect 3680 -1289 3696 -1255
rect 3864 -1289 3880 -1255
rect 3680 -1327 3880 -1289
rect 4058 -1255 4258 -1239
rect 4058 -1289 4074 -1255
rect 4242 -1289 4258 -1255
rect 4058 -1327 4258 -1289
rect 4436 -1255 4636 -1239
rect 4436 -1289 4452 -1255
rect 4620 -1289 4636 -1255
rect 4436 -1327 4636 -1289
rect -4636 -2365 -4436 -2327
rect -4636 -2399 -4620 -2365
rect -4452 -2399 -4436 -2365
rect -4636 -2415 -4436 -2399
rect -4258 -2365 -4058 -2327
rect -4258 -2399 -4242 -2365
rect -4074 -2399 -4058 -2365
rect -4258 -2415 -4058 -2399
rect -3880 -2365 -3680 -2327
rect -3880 -2399 -3864 -2365
rect -3696 -2399 -3680 -2365
rect -3880 -2415 -3680 -2399
rect -3502 -2365 -3302 -2327
rect -3502 -2399 -3486 -2365
rect -3318 -2399 -3302 -2365
rect -3502 -2415 -3302 -2399
rect -3124 -2365 -2924 -2327
rect -3124 -2399 -3108 -2365
rect -2940 -2399 -2924 -2365
rect -3124 -2415 -2924 -2399
rect -2746 -2365 -2546 -2327
rect -2746 -2399 -2730 -2365
rect -2562 -2399 -2546 -2365
rect -2746 -2415 -2546 -2399
rect -2368 -2365 -2168 -2327
rect -2368 -2399 -2352 -2365
rect -2184 -2399 -2168 -2365
rect -2368 -2415 -2168 -2399
rect -1990 -2365 -1790 -2327
rect -1990 -2399 -1974 -2365
rect -1806 -2399 -1790 -2365
rect -1990 -2415 -1790 -2399
rect -1612 -2365 -1412 -2327
rect -1612 -2399 -1596 -2365
rect -1428 -2399 -1412 -2365
rect -1612 -2415 -1412 -2399
rect -1234 -2365 -1034 -2327
rect -1234 -2399 -1218 -2365
rect -1050 -2399 -1034 -2365
rect -1234 -2415 -1034 -2399
rect -856 -2365 -656 -2327
rect -856 -2399 -840 -2365
rect -672 -2399 -656 -2365
rect -856 -2415 -656 -2399
rect -478 -2365 -278 -2327
rect -478 -2399 -462 -2365
rect -294 -2399 -278 -2365
rect -478 -2415 -278 -2399
rect -100 -2365 100 -2327
rect -100 -2399 -84 -2365
rect 84 -2399 100 -2365
rect -100 -2415 100 -2399
rect 278 -2365 478 -2327
rect 278 -2399 294 -2365
rect 462 -2399 478 -2365
rect 278 -2415 478 -2399
rect 656 -2365 856 -2327
rect 656 -2399 672 -2365
rect 840 -2399 856 -2365
rect 656 -2415 856 -2399
rect 1034 -2365 1234 -2327
rect 1034 -2399 1050 -2365
rect 1218 -2399 1234 -2365
rect 1034 -2415 1234 -2399
rect 1412 -2365 1612 -2327
rect 1412 -2399 1428 -2365
rect 1596 -2399 1612 -2365
rect 1412 -2415 1612 -2399
rect 1790 -2365 1990 -2327
rect 1790 -2399 1806 -2365
rect 1974 -2399 1990 -2365
rect 1790 -2415 1990 -2399
rect 2168 -2365 2368 -2327
rect 2168 -2399 2184 -2365
rect 2352 -2399 2368 -2365
rect 2168 -2415 2368 -2399
rect 2546 -2365 2746 -2327
rect 2546 -2399 2562 -2365
rect 2730 -2399 2746 -2365
rect 2546 -2415 2746 -2399
rect 2924 -2365 3124 -2327
rect 2924 -2399 2940 -2365
rect 3108 -2399 3124 -2365
rect 2924 -2415 3124 -2399
rect 3302 -2365 3502 -2327
rect 3302 -2399 3318 -2365
rect 3486 -2399 3502 -2365
rect 3302 -2415 3502 -2399
rect 3680 -2365 3880 -2327
rect 3680 -2399 3696 -2365
rect 3864 -2399 3880 -2365
rect 3680 -2415 3880 -2399
rect 4058 -2365 4258 -2327
rect 4058 -2399 4074 -2365
rect 4242 -2399 4258 -2365
rect 4058 -2415 4258 -2399
rect 4436 -2365 4636 -2327
rect 4436 -2399 4452 -2365
rect 4620 -2399 4636 -2365
rect 4436 -2415 4636 -2399
<< polycont >>
rect -4620 2365 -4452 2399
rect -4242 2365 -4074 2399
rect -3864 2365 -3696 2399
rect -3486 2365 -3318 2399
rect -3108 2365 -2940 2399
rect -2730 2365 -2562 2399
rect -2352 2365 -2184 2399
rect -1974 2365 -1806 2399
rect -1596 2365 -1428 2399
rect -1218 2365 -1050 2399
rect -840 2365 -672 2399
rect -462 2365 -294 2399
rect -84 2365 84 2399
rect 294 2365 462 2399
rect 672 2365 840 2399
rect 1050 2365 1218 2399
rect 1428 2365 1596 2399
rect 1806 2365 1974 2399
rect 2184 2365 2352 2399
rect 2562 2365 2730 2399
rect 2940 2365 3108 2399
rect 3318 2365 3486 2399
rect 3696 2365 3864 2399
rect 4074 2365 4242 2399
rect 4452 2365 4620 2399
rect -4620 1255 -4452 1289
rect -4242 1255 -4074 1289
rect -3864 1255 -3696 1289
rect -3486 1255 -3318 1289
rect -3108 1255 -2940 1289
rect -2730 1255 -2562 1289
rect -2352 1255 -2184 1289
rect -1974 1255 -1806 1289
rect -1596 1255 -1428 1289
rect -1218 1255 -1050 1289
rect -840 1255 -672 1289
rect -462 1255 -294 1289
rect -84 1255 84 1289
rect 294 1255 462 1289
rect 672 1255 840 1289
rect 1050 1255 1218 1289
rect 1428 1255 1596 1289
rect 1806 1255 1974 1289
rect 2184 1255 2352 1289
rect 2562 1255 2730 1289
rect 2940 1255 3108 1289
rect 3318 1255 3486 1289
rect 3696 1255 3864 1289
rect 4074 1255 4242 1289
rect 4452 1255 4620 1289
rect -4620 1147 -4452 1181
rect -4242 1147 -4074 1181
rect -3864 1147 -3696 1181
rect -3486 1147 -3318 1181
rect -3108 1147 -2940 1181
rect -2730 1147 -2562 1181
rect -2352 1147 -2184 1181
rect -1974 1147 -1806 1181
rect -1596 1147 -1428 1181
rect -1218 1147 -1050 1181
rect -840 1147 -672 1181
rect -462 1147 -294 1181
rect -84 1147 84 1181
rect 294 1147 462 1181
rect 672 1147 840 1181
rect 1050 1147 1218 1181
rect 1428 1147 1596 1181
rect 1806 1147 1974 1181
rect 2184 1147 2352 1181
rect 2562 1147 2730 1181
rect 2940 1147 3108 1181
rect 3318 1147 3486 1181
rect 3696 1147 3864 1181
rect 4074 1147 4242 1181
rect 4452 1147 4620 1181
rect -4620 37 -4452 71
rect -4242 37 -4074 71
rect -3864 37 -3696 71
rect -3486 37 -3318 71
rect -3108 37 -2940 71
rect -2730 37 -2562 71
rect -2352 37 -2184 71
rect -1974 37 -1806 71
rect -1596 37 -1428 71
rect -1218 37 -1050 71
rect -840 37 -672 71
rect -462 37 -294 71
rect -84 37 84 71
rect 294 37 462 71
rect 672 37 840 71
rect 1050 37 1218 71
rect 1428 37 1596 71
rect 1806 37 1974 71
rect 2184 37 2352 71
rect 2562 37 2730 71
rect 2940 37 3108 71
rect 3318 37 3486 71
rect 3696 37 3864 71
rect 4074 37 4242 71
rect 4452 37 4620 71
rect -4620 -71 -4452 -37
rect -4242 -71 -4074 -37
rect -3864 -71 -3696 -37
rect -3486 -71 -3318 -37
rect -3108 -71 -2940 -37
rect -2730 -71 -2562 -37
rect -2352 -71 -2184 -37
rect -1974 -71 -1806 -37
rect -1596 -71 -1428 -37
rect -1218 -71 -1050 -37
rect -840 -71 -672 -37
rect -462 -71 -294 -37
rect -84 -71 84 -37
rect 294 -71 462 -37
rect 672 -71 840 -37
rect 1050 -71 1218 -37
rect 1428 -71 1596 -37
rect 1806 -71 1974 -37
rect 2184 -71 2352 -37
rect 2562 -71 2730 -37
rect 2940 -71 3108 -37
rect 3318 -71 3486 -37
rect 3696 -71 3864 -37
rect 4074 -71 4242 -37
rect 4452 -71 4620 -37
rect -4620 -1181 -4452 -1147
rect -4242 -1181 -4074 -1147
rect -3864 -1181 -3696 -1147
rect -3486 -1181 -3318 -1147
rect -3108 -1181 -2940 -1147
rect -2730 -1181 -2562 -1147
rect -2352 -1181 -2184 -1147
rect -1974 -1181 -1806 -1147
rect -1596 -1181 -1428 -1147
rect -1218 -1181 -1050 -1147
rect -840 -1181 -672 -1147
rect -462 -1181 -294 -1147
rect -84 -1181 84 -1147
rect 294 -1181 462 -1147
rect 672 -1181 840 -1147
rect 1050 -1181 1218 -1147
rect 1428 -1181 1596 -1147
rect 1806 -1181 1974 -1147
rect 2184 -1181 2352 -1147
rect 2562 -1181 2730 -1147
rect 2940 -1181 3108 -1147
rect 3318 -1181 3486 -1147
rect 3696 -1181 3864 -1147
rect 4074 -1181 4242 -1147
rect 4452 -1181 4620 -1147
rect -4620 -1289 -4452 -1255
rect -4242 -1289 -4074 -1255
rect -3864 -1289 -3696 -1255
rect -3486 -1289 -3318 -1255
rect -3108 -1289 -2940 -1255
rect -2730 -1289 -2562 -1255
rect -2352 -1289 -2184 -1255
rect -1974 -1289 -1806 -1255
rect -1596 -1289 -1428 -1255
rect -1218 -1289 -1050 -1255
rect -840 -1289 -672 -1255
rect -462 -1289 -294 -1255
rect -84 -1289 84 -1255
rect 294 -1289 462 -1255
rect 672 -1289 840 -1255
rect 1050 -1289 1218 -1255
rect 1428 -1289 1596 -1255
rect 1806 -1289 1974 -1255
rect 2184 -1289 2352 -1255
rect 2562 -1289 2730 -1255
rect 2940 -1289 3108 -1255
rect 3318 -1289 3486 -1255
rect 3696 -1289 3864 -1255
rect 4074 -1289 4242 -1255
rect 4452 -1289 4620 -1255
rect -4620 -2399 -4452 -2365
rect -4242 -2399 -4074 -2365
rect -3864 -2399 -3696 -2365
rect -3486 -2399 -3318 -2365
rect -3108 -2399 -2940 -2365
rect -2730 -2399 -2562 -2365
rect -2352 -2399 -2184 -2365
rect -1974 -2399 -1806 -2365
rect -1596 -2399 -1428 -2365
rect -1218 -2399 -1050 -2365
rect -840 -2399 -672 -2365
rect -462 -2399 -294 -2365
rect -84 -2399 84 -2365
rect 294 -2399 462 -2365
rect 672 -2399 840 -2365
rect 1050 -2399 1218 -2365
rect 1428 -2399 1596 -2365
rect 1806 -2399 1974 -2365
rect 2184 -2399 2352 -2365
rect 2562 -2399 2730 -2365
rect 2940 -2399 3108 -2365
rect 3318 -2399 3486 -2365
rect 3696 -2399 3864 -2365
rect 4074 -2399 4242 -2365
rect 4452 -2399 4620 -2365
<< locali >>
rect -4816 2503 -4720 2537
rect 4720 2503 4816 2537
rect -4816 2441 -4782 2503
rect 4782 2441 4816 2503
rect -4636 2365 -4620 2399
rect -4452 2365 -4436 2399
rect -4258 2365 -4242 2399
rect -4074 2365 -4058 2399
rect -3880 2365 -3864 2399
rect -3696 2365 -3680 2399
rect -3502 2365 -3486 2399
rect -3318 2365 -3302 2399
rect -3124 2365 -3108 2399
rect -2940 2365 -2924 2399
rect -2746 2365 -2730 2399
rect -2562 2365 -2546 2399
rect -2368 2365 -2352 2399
rect -2184 2365 -2168 2399
rect -1990 2365 -1974 2399
rect -1806 2365 -1790 2399
rect -1612 2365 -1596 2399
rect -1428 2365 -1412 2399
rect -1234 2365 -1218 2399
rect -1050 2365 -1034 2399
rect -856 2365 -840 2399
rect -672 2365 -656 2399
rect -478 2365 -462 2399
rect -294 2365 -278 2399
rect -100 2365 -84 2399
rect 84 2365 100 2399
rect 278 2365 294 2399
rect 462 2365 478 2399
rect 656 2365 672 2399
rect 840 2365 856 2399
rect 1034 2365 1050 2399
rect 1218 2365 1234 2399
rect 1412 2365 1428 2399
rect 1596 2365 1612 2399
rect 1790 2365 1806 2399
rect 1974 2365 1990 2399
rect 2168 2365 2184 2399
rect 2352 2365 2368 2399
rect 2546 2365 2562 2399
rect 2730 2365 2746 2399
rect 2924 2365 2940 2399
rect 3108 2365 3124 2399
rect 3302 2365 3318 2399
rect 3486 2365 3502 2399
rect 3680 2365 3696 2399
rect 3864 2365 3880 2399
rect 4058 2365 4074 2399
rect 4242 2365 4258 2399
rect 4436 2365 4452 2399
rect 4620 2365 4636 2399
rect -4682 2315 -4648 2331
rect -4682 1323 -4648 1339
rect -4424 2315 -4390 2331
rect -4424 1323 -4390 1339
rect -4304 2315 -4270 2331
rect -4304 1323 -4270 1339
rect -4046 2315 -4012 2331
rect -4046 1323 -4012 1339
rect -3926 2315 -3892 2331
rect -3926 1323 -3892 1339
rect -3668 2315 -3634 2331
rect -3668 1323 -3634 1339
rect -3548 2315 -3514 2331
rect -3548 1323 -3514 1339
rect -3290 2315 -3256 2331
rect -3290 1323 -3256 1339
rect -3170 2315 -3136 2331
rect -3170 1323 -3136 1339
rect -2912 2315 -2878 2331
rect -2912 1323 -2878 1339
rect -2792 2315 -2758 2331
rect -2792 1323 -2758 1339
rect -2534 2315 -2500 2331
rect -2534 1323 -2500 1339
rect -2414 2315 -2380 2331
rect -2414 1323 -2380 1339
rect -2156 2315 -2122 2331
rect -2156 1323 -2122 1339
rect -2036 2315 -2002 2331
rect -2036 1323 -2002 1339
rect -1778 2315 -1744 2331
rect -1778 1323 -1744 1339
rect -1658 2315 -1624 2331
rect -1658 1323 -1624 1339
rect -1400 2315 -1366 2331
rect -1400 1323 -1366 1339
rect -1280 2315 -1246 2331
rect -1280 1323 -1246 1339
rect -1022 2315 -988 2331
rect -1022 1323 -988 1339
rect -902 2315 -868 2331
rect -902 1323 -868 1339
rect -644 2315 -610 2331
rect -644 1323 -610 1339
rect -524 2315 -490 2331
rect -524 1323 -490 1339
rect -266 2315 -232 2331
rect -266 1323 -232 1339
rect -146 2315 -112 2331
rect -146 1323 -112 1339
rect 112 2315 146 2331
rect 112 1323 146 1339
rect 232 2315 266 2331
rect 232 1323 266 1339
rect 490 2315 524 2331
rect 490 1323 524 1339
rect 610 2315 644 2331
rect 610 1323 644 1339
rect 868 2315 902 2331
rect 868 1323 902 1339
rect 988 2315 1022 2331
rect 988 1323 1022 1339
rect 1246 2315 1280 2331
rect 1246 1323 1280 1339
rect 1366 2315 1400 2331
rect 1366 1323 1400 1339
rect 1624 2315 1658 2331
rect 1624 1323 1658 1339
rect 1744 2315 1778 2331
rect 1744 1323 1778 1339
rect 2002 2315 2036 2331
rect 2002 1323 2036 1339
rect 2122 2315 2156 2331
rect 2122 1323 2156 1339
rect 2380 2315 2414 2331
rect 2380 1323 2414 1339
rect 2500 2315 2534 2331
rect 2500 1323 2534 1339
rect 2758 2315 2792 2331
rect 2758 1323 2792 1339
rect 2878 2315 2912 2331
rect 2878 1323 2912 1339
rect 3136 2315 3170 2331
rect 3136 1323 3170 1339
rect 3256 2315 3290 2331
rect 3256 1323 3290 1339
rect 3514 2315 3548 2331
rect 3514 1323 3548 1339
rect 3634 2315 3668 2331
rect 3634 1323 3668 1339
rect 3892 2315 3926 2331
rect 3892 1323 3926 1339
rect 4012 2315 4046 2331
rect 4012 1323 4046 1339
rect 4270 2315 4304 2331
rect 4270 1323 4304 1339
rect 4390 2315 4424 2331
rect 4390 1323 4424 1339
rect 4648 2315 4682 2331
rect 4648 1323 4682 1339
rect -4636 1255 -4620 1289
rect -4452 1255 -4436 1289
rect -4258 1255 -4242 1289
rect -4074 1255 -4058 1289
rect -3880 1255 -3864 1289
rect -3696 1255 -3680 1289
rect -3502 1255 -3486 1289
rect -3318 1255 -3302 1289
rect -3124 1255 -3108 1289
rect -2940 1255 -2924 1289
rect -2746 1255 -2730 1289
rect -2562 1255 -2546 1289
rect -2368 1255 -2352 1289
rect -2184 1255 -2168 1289
rect -1990 1255 -1974 1289
rect -1806 1255 -1790 1289
rect -1612 1255 -1596 1289
rect -1428 1255 -1412 1289
rect -1234 1255 -1218 1289
rect -1050 1255 -1034 1289
rect -856 1255 -840 1289
rect -672 1255 -656 1289
rect -478 1255 -462 1289
rect -294 1255 -278 1289
rect -100 1255 -84 1289
rect 84 1255 100 1289
rect 278 1255 294 1289
rect 462 1255 478 1289
rect 656 1255 672 1289
rect 840 1255 856 1289
rect 1034 1255 1050 1289
rect 1218 1255 1234 1289
rect 1412 1255 1428 1289
rect 1596 1255 1612 1289
rect 1790 1255 1806 1289
rect 1974 1255 1990 1289
rect 2168 1255 2184 1289
rect 2352 1255 2368 1289
rect 2546 1255 2562 1289
rect 2730 1255 2746 1289
rect 2924 1255 2940 1289
rect 3108 1255 3124 1289
rect 3302 1255 3318 1289
rect 3486 1255 3502 1289
rect 3680 1255 3696 1289
rect 3864 1255 3880 1289
rect 4058 1255 4074 1289
rect 4242 1255 4258 1289
rect 4436 1255 4452 1289
rect 4620 1255 4636 1289
rect -4636 1147 -4620 1181
rect -4452 1147 -4436 1181
rect -4258 1147 -4242 1181
rect -4074 1147 -4058 1181
rect -3880 1147 -3864 1181
rect -3696 1147 -3680 1181
rect -3502 1147 -3486 1181
rect -3318 1147 -3302 1181
rect -3124 1147 -3108 1181
rect -2940 1147 -2924 1181
rect -2746 1147 -2730 1181
rect -2562 1147 -2546 1181
rect -2368 1147 -2352 1181
rect -2184 1147 -2168 1181
rect -1990 1147 -1974 1181
rect -1806 1147 -1790 1181
rect -1612 1147 -1596 1181
rect -1428 1147 -1412 1181
rect -1234 1147 -1218 1181
rect -1050 1147 -1034 1181
rect -856 1147 -840 1181
rect -672 1147 -656 1181
rect -478 1147 -462 1181
rect -294 1147 -278 1181
rect -100 1147 -84 1181
rect 84 1147 100 1181
rect 278 1147 294 1181
rect 462 1147 478 1181
rect 656 1147 672 1181
rect 840 1147 856 1181
rect 1034 1147 1050 1181
rect 1218 1147 1234 1181
rect 1412 1147 1428 1181
rect 1596 1147 1612 1181
rect 1790 1147 1806 1181
rect 1974 1147 1990 1181
rect 2168 1147 2184 1181
rect 2352 1147 2368 1181
rect 2546 1147 2562 1181
rect 2730 1147 2746 1181
rect 2924 1147 2940 1181
rect 3108 1147 3124 1181
rect 3302 1147 3318 1181
rect 3486 1147 3502 1181
rect 3680 1147 3696 1181
rect 3864 1147 3880 1181
rect 4058 1147 4074 1181
rect 4242 1147 4258 1181
rect 4436 1147 4452 1181
rect 4620 1147 4636 1181
rect -4682 1097 -4648 1113
rect -4682 105 -4648 121
rect -4424 1097 -4390 1113
rect -4424 105 -4390 121
rect -4304 1097 -4270 1113
rect -4304 105 -4270 121
rect -4046 1097 -4012 1113
rect -4046 105 -4012 121
rect -3926 1097 -3892 1113
rect -3926 105 -3892 121
rect -3668 1097 -3634 1113
rect -3668 105 -3634 121
rect -3548 1097 -3514 1113
rect -3548 105 -3514 121
rect -3290 1097 -3256 1113
rect -3290 105 -3256 121
rect -3170 1097 -3136 1113
rect -3170 105 -3136 121
rect -2912 1097 -2878 1113
rect -2912 105 -2878 121
rect -2792 1097 -2758 1113
rect -2792 105 -2758 121
rect -2534 1097 -2500 1113
rect -2534 105 -2500 121
rect -2414 1097 -2380 1113
rect -2414 105 -2380 121
rect -2156 1097 -2122 1113
rect -2156 105 -2122 121
rect -2036 1097 -2002 1113
rect -2036 105 -2002 121
rect -1778 1097 -1744 1113
rect -1778 105 -1744 121
rect -1658 1097 -1624 1113
rect -1658 105 -1624 121
rect -1400 1097 -1366 1113
rect -1400 105 -1366 121
rect -1280 1097 -1246 1113
rect -1280 105 -1246 121
rect -1022 1097 -988 1113
rect -1022 105 -988 121
rect -902 1097 -868 1113
rect -902 105 -868 121
rect -644 1097 -610 1113
rect -644 105 -610 121
rect -524 1097 -490 1113
rect -524 105 -490 121
rect -266 1097 -232 1113
rect -266 105 -232 121
rect -146 1097 -112 1113
rect -146 105 -112 121
rect 112 1097 146 1113
rect 112 105 146 121
rect 232 1097 266 1113
rect 232 105 266 121
rect 490 1097 524 1113
rect 490 105 524 121
rect 610 1097 644 1113
rect 610 105 644 121
rect 868 1097 902 1113
rect 868 105 902 121
rect 988 1097 1022 1113
rect 988 105 1022 121
rect 1246 1097 1280 1113
rect 1246 105 1280 121
rect 1366 1097 1400 1113
rect 1366 105 1400 121
rect 1624 1097 1658 1113
rect 1624 105 1658 121
rect 1744 1097 1778 1113
rect 1744 105 1778 121
rect 2002 1097 2036 1113
rect 2002 105 2036 121
rect 2122 1097 2156 1113
rect 2122 105 2156 121
rect 2380 1097 2414 1113
rect 2380 105 2414 121
rect 2500 1097 2534 1113
rect 2500 105 2534 121
rect 2758 1097 2792 1113
rect 2758 105 2792 121
rect 2878 1097 2912 1113
rect 2878 105 2912 121
rect 3136 1097 3170 1113
rect 3136 105 3170 121
rect 3256 1097 3290 1113
rect 3256 105 3290 121
rect 3514 1097 3548 1113
rect 3514 105 3548 121
rect 3634 1097 3668 1113
rect 3634 105 3668 121
rect 3892 1097 3926 1113
rect 3892 105 3926 121
rect 4012 1097 4046 1113
rect 4012 105 4046 121
rect 4270 1097 4304 1113
rect 4270 105 4304 121
rect 4390 1097 4424 1113
rect 4390 105 4424 121
rect 4648 1097 4682 1113
rect 4648 105 4682 121
rect -4636 37 -4620 71
rect -4452 37 -4436 71
rect -4258 37 -4242 71
rect -4074 37 -4058 71
rect -3880 37 -3864 71
rect -3696 37 -3680 71
rect -3502 37 -3486 71
rect -3318 37 -3302 71
rect -3124 37 -3108 71
rect -2940 37 -2924 71
rect -2746 37 -2730 71
rect -2562 37 -2546 71
rect -2368 37 -2352 71
rect -2184 37 -2168 71
rect -1990 37 -1974 71
rect -1806 37 -1790 71
rect -1612 37 -1596 71
rect -1428 37 -1412 71
rect -1234 37 -1218 71
rect -1050 37 -1034 71
rect -856 37 -840 71
rect -672 37 -656 71
rect -478 37 -462 71
rect -294 37 -278 71
rect -100 37 -84 71
rect 84 37 100 71
rect 278 37 294 71
rect 462 37 478 71
rect 656 37 672 71
rect 840 37 856 71
rect 1034 37 1050 71
rect 1218 37 1234 71
rect 1412 37 1428 71
rect 1596 37 1612 71
rect 1790 37 1806 71
rect 1974 37 1990 71
rect 2168 37 2184 71
rect 2352 37 2368 71
rect 2546 37 2562 71
rect 2730 37 2746 71
rect 2924 37 2940 71
rect 3108 37 3124 71
rect 3302 37 3318 71
rect 3486 37 3502 71
rect 3680 37 3696 71
rect 3864 37 3880 71
rect 4058 37 4074 71
rect 4242 37 4258 71
rect 4436 37 4452 71
rect 4620 37 4636 71
rect -4636 -71 -4620 -37
rect -4452 -71 -4436 -37
rect -4258 -71 -4242 -37
rect -4074 -71 -4058 -37
rect -3880 -71 -3864 -37
rect -3696 -71 -3680 -37
rect -3502 -71 -3486 -37
rect -3318 -71 -3302 -37
rect -3124 -71 -3108 -37
rect -2940 -71 -2924 -37
rect -2746 -71 -2730 -37
rect -2562 -71 -2546 -37
rect -2368 -71 -2352 -37
rect -2184 -71 -2168 -37
rect -1990 -71 -1974 -37
rect -1806 -71 -1790 -37
rect -1612 -71 -1596 -37
rect -1428 -71 -1412 -37
rect -1234 -71 -1218 -37
rect -1050 -71 -1034 -37
rect -856 -71 -840 -37
rect -672 -71 -656 -37
rect -478 -71 -462 -37
rect -294 -71 -278 -37
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect 278 -71 294 -37
rect 462 -71 478 -37
rect 656 -71 672 -37
rect 840 -71 856 -37
rect 1034 -71 1050 -37
rect 1218 -71 1234 -37
rect 1412 -71 1428 -37
rect 1596 -71 1612 -37
rect 1790 -71 1806 -37
rect 1974 -71 1990 -37
rect 2168 -71 2184 -37
rect 2352 -71 2368 -37
rect 2546 -71 2562 -37
rect 2730 -71 2746 -37
rect 2924 -71 2940 -37
rect 3108 -71 3124 -37
rect 3302 -71 3318 -37
rect 3486 -71 3502 -37
rect 3680 -71 3696 -37
rect 3864 -71 3880 -37
rect 4058 -71 4074 -37
rect 4242 -71 4258 -37
rect 4436 -71 4452 -37
rect 4620 -71 4636 -37
rect -4682 -121 -4648 -105
rect -4682 -1113 -4648 -1097
rect -4424 -121 -4390 -105
rect -4424 -1113 -4390 -1097
rect -4304 -121 -4270 -105
rect -4304 -1113 -4270 -1097
rect -4046 -121 -4012 -105
rect -4046 -1113 -4012 -1097
rect -3926 -121 -3892 -105
rect -3926 -1113 -3892 -1097
rect -3668 -121 -3634 -105
rect -3668 -1113 -3634 -1097
rect -3548 -121 -3514 -105
rect -3548 -1113 -3514 -1097
rect -3290 -121 -3256 -105
rect -3290 -1113 -3256 -1097
rect -3170 -121 -3136 -105
rect -3170 -1113 -3136 -1097
rect -2912 -121 -2878 -105
rect -2912 -1113 -2878 -1097
rect -2792 -121 -2758 -105
rect -2792 -1113 -2758 -1097
rect -2534 -121 -2500 -105
rect -2534 -1113 -2500 -1097
rect -2414 -121 -2380 -105
rect -2414 -1113 -2380 -1097
rect -2156 -121 -2122 -105
rect -2156 -1113 -2122 -1097
rect -2036 -121 -2002 -105
rect -2036 -1113 -2002 -1097
rect -1778 -121 -1744 -105
rect -1778 -1113 -1744 -1097
rect -1658 -121 -1624 -105
rect -1658 -1113 -1624 -1097
rect -1400 -121 -1366 -105
rect -1400 -1113 -1366 -1097
rect -1280 -121 -1246 -105
rect -1280 -1113 -1246 -1097
rect -1022 -121 -988 -105
rect -1022 -1113 -988 -1097
rect -902 -121 -868 -105
rect -902 -1113 -868 -1097
rect -644 -121 -610 -105
rect -644 -1113 -610 -1097
rect -524 -121 -490 -105
rect -524 -1113 -490 -1097
rect -266 -121 -232 -105
rect -266 -1113 -232 -1097
rect -146 -121 -112 -105
rect -146 -1113 -112 -1097
rect 112 -121 146 -105
rect 112 -1113 146 -1097
rect 232 -121 266 -105
rect 232 -1113 266 -1097
rect 490 -121 524 -105
rect 490 -1113 524 -1097
rect 610 -121 644 -105
rect 610 -1113 644 -1097
rect 868 -121 902 -105
rect 868 -1113 902 -1097
rect 988 -121 1022 -105
rect 988 -1113 1022 -1097
rect 1246 -121 1280 -105
rect 1246 -1113 1280 -1097
rect 1366 -121 1400 -105
rect 1366 -1113 1400 -1097
rect 1624 -121 1658 -105
rect 1624 -1113 1658 -1097
rect 1744 -121 1778 -105
rect 1744 -1113 1778 -1097
rect 2002 -121 2036 -105
rect 2002 -1113 2036 -1097
rect 2122 -121 2156 -105
rect 2122 -1113 2156 -1097
rect 2380 -121 2414 -105
rect 2380 -1113 2414 -1097
rect 2500 -121 2534 -105
rect 2500 -1113 2534 -1097
rect 2758 -121 2792 -105
rect 2758 -1113 2792 -1097
rect 2878 -121 2912 -105
rect 2878 -1113 2912 -1097
rect 3136 -121 3170 -105
rect 3136 -1113 3170 -1097
rect 3256 -121 3290 -105
rect 3256 -1113 3290 -1097
rect 3514 -121 3548 -105
rect 3514 -1113 3548 -1097
rect 3634 -121 3668 -105
rect 3634 -1113 3668 -1097
rect 3892 -121 3926 -105
rect 3892 -1113 3926 -1097
rect 4012 -121 4046 -105
rect 4012 -1113 4046 -1097
rect 4270 -121 4304 -105
rect 4270 -1113 4304 -1097
rect 4390 -121 4424 -105
rect 4390 -1113 4424 -1097
rect 4648 -121 4682 -105
rect 4648 -1113 4682 -1097
rect -4636 -1181 -4620 -1147
rect -4452 -1181 -4436 -1147
rect -4258 -1181 -4242 -1147
rect -4074 -1181 -4058 -1147
rect -3880 -1181 -3864 -1147
rect -3696 -1181 -3680 -1147
rect -3502 -1181 -3486 -1147
rect -3318 -1181 -3302 -1147
rect -3124 -1181 -3108 -1147
rect -2940 -1181 -2924 -1147
rect -2746 -1181 -2730 -1147
rect -2562 -1181 -2546 -1147
rect -2368 -1181 -2352 -1147
rect -2184 -1181 -2168 -1147
rect -1990 -1181 -1974 -1147
rect -1806 -1181 -1790 -1147
rect -1612 -1181 -1596 -1147
rect -1428 -1181 -1412 -1147
rect -1234 -1181 -1218 -1147
rect -1050 -1181 -1034 -1147
rect -856 -1181 -840 -1147
rect -672 -1181 -656 -1147
rect -478 -1181 -462 -1147
rect -294 -1181 -278 -1147
rect -100 -1181 -84 -1147
rect 84 -1181 100 -1147
rect 278 -1181 294 -1147
rect 462 -1181 478 -1147
rect 656 -1181 672 -1147
rect 840 -1181 856 -1147
rect 1034 -1181 1050 -1147
rect 1218 -1181 1234 -1147
rect 1412 -1181 1428 -1147
rect 1596 -1181 1612 -1147
rect 1790 -1181 1806 -1147
rect 1974 -1181 1990 -1147
rect 2168 -1181 2184 -1147
rect 2352 -1181 2368 -1147
rect 2546 -1181 2562 -1147
rect 2730 -1181 2746 -1147
rect 2924 -1181 2940 -1147
rect 3108 -1181 3124 -1147
rect 3302 -1181 3318 -1147
rect 3486 -1181 3502 -1147
rect 3680 -1181 3696 -1147
rect 3864 -1181 3880 -1147
rect 4058 -1181 4074 -1147
rect 4242 -1181 4258 -1147
rect 4436 -1181 4452 -1147
rect 4620 -1181 4636 -1147
rect -4636 -1289 -4620 -1255
rect -4452 -1289 -4436 -1255
rect -4258 -1289 -4242 -1255
rect -4074 -1289 -4058 -1255
rect -3880 -1289 -3864 -1255
rect -3696 -1289 -3680 -1255
rect -3502 -1289 -3486 -1255
rect -3318 -1289 -3302 -1255
rect -3124 -1289 -3108 -1255
rect -2940 -1289 -2924 -1255
rect -2746 -1289 -2730 -1255
rect -2562 -1289 -2546 -1255
rect -2368 -1289 -2352 -1255
rect -2184 -1289 -2168 -1255
rect -1990 -1289 -1974 -1255
rect -1806 -1289 -1790 -1255
rect -1612 -1289 -1596 -1255
rect -1428 -1289 -1412 -1255
rect -1234 -1289 -1218 -1255
rect -1050 -1289 -1034 -1255
rect -856 -1289 -840 -1255
rect -672 -1289 -656 -1255
rect -478 -1289 -462 -1255
rect -294 -1289 -278 -1255
rect -100 -1289 -84 -1255
rect 84 -1289 100 -1255
rect 278 -1289 294 -1255
rect 462 -1289 478 -1255
rect 656 -1289 672 -1255
rect 840 -1289 856 -1255
rect 1034 -1289 1050 -1255
rect 1218 -1289 1234 -1255
rect 1412 -1289 1428 -1255
rect 1596 -1289 1612 -1255
rect 1790 -1289 1806 -1255
rect 1974 -1289 1990 -1255
rect 2168 -1289 2184 -1255
rect 2352 -1289 2368 -1255
rect 2546 -1289 2562 -1255
rect 2730 -1289 2746 -1255
rect 2924 -1289 2940 -1255
rect 3108 -1289 3124 -1255
rect 3302 -1289 3318 -1255
rect 3486 -1289 3502 -1255
rect 3680 -1289 3696 -1255
rect 3864 -1289 3880 -1255
rect 4058 -1289 4074 -1255
rect 4242 -1289 4258 -1255
rect 4436 -1289 4452 -1255
rect 4620 -1289 4636 -1255
rect -4682 -1339 -4648 -1323
rect -4682 -2331 -4648 -2315
rect -4424 -1339 -4390 -1323
rect -4424 -2331 -4390 -2315
rect -4304 -1339 -4270 -1323
rect -4304 -2331 -4270 -2315
rect -4046 -1339 -4012 -1323
rect -4046 -2331 -4012 -2315
rect -3926 -1339 -3892 -1323
rect -3926 -2331 -3892 -2315
rect -3668 -1339 -3634 -1323
rect -3668 -2331 -3634 -2315
rect -3548 -1339 -3514 -1323
rect -3548 -2331 -3514 -2315
rect -3290 -1339 -3256 -1323
rect -3290 -2331 -3256 -2315
rect -3170 -1339 -3136 -1323
rect -3170 -2331 -3136 -2315
rect -2912 -1339 -2878 -1323
rect -2912 -2331 -2878 -2315
rect -2792 -1339 -2758 -1323
rect -2792 -2331 -2758 -2315
rect -2534 -1339 -2500 -1323
rect -2534 -2331 -2500 -2315
rect -2414 -1339 -2380 -1323
rect -2414 -2331 -2380 -2315
rect -2156 -1339 -2122 -1323
rect -2156 -2331 -2122 -2315
rect -2036 -1339 -2002 -1323
rect -2036 -2331 -2002 -2315
rect -1778 -1339 -1744 -1323
rect -1778 -2331 -1744 -2315
rect -1658 -1339 -1624 -1323
rect -1658 -2331 -1624 -2315
rect -1400 -1339 -1366 -1323
rect -1400 -2331 -1366 -2315
rect -1280 -1339 -1246 -1323
rect -1280 -2331 -1246 -2315
rect -1022 -1339 -988 -1323
rect -1022 -2331 -988 -2315
rect -902 -1339 -868 -1323
rect -902 -2331 -868 -2315
rect -644 -1339 -610 -1323
rect -644 -2331 -610 -2315
rect -524 -1339 -490 -1323
rect -524 -2331 -490 -2315
rect -266 -1339 -232 -1323
rect -266 -2331 -232 -2315
rect -146 -1339 -112 -1323
rect -146 -2331 -112 -2315
rect 112 -1339 146 -1323
rect 112 -2331 146 -2315
rect 232 -1339 266 -1323
rect 232 -2331 266 -2315
rect 490 -1339 524 -1323
rect 490 -2331 524 -2315
rect 610 -1339 644 -1323
rect 610 -2331 644 -2315
rect 868 -1339 902 -1323
rect 868 -2331 902 -2315
rect 988 -1339 1022 -1323
rect 988 -2331 1022 -2315
rect 1246 -1339 1280 -1323
rect 1246 -2331 1280 -2315
rect 1366 -1339 1400 -1323
rect 1366 -2331 1400 -2315
rect 1624 -1339 1658 -1323
rect 1624 -2331 1658 -2315
rect 1744 -1339 1778 -1323
rect 1744 -2331 1778 -2315
rect 2002 -1339 2036 -1323
rect 2002 -2331 2036 -2315
rect 2122 -1339 2156 -1323
rect 2122 -2331 2156 -2315
rect 2380 -1339 2414 -1323
rect 2380 -2331 2414 -2315
rect 2500 -1339 2534 -1323
rect 2500 -2331 2534 -2315
rect 2758 -1339 2792 -1323
rect 2758 -2331 2792 -2315
rect 2878 -1339 2912 -1323
rect 2878 -2331 2912 -2315
rect 3136 -1339 3170 -1323
rect 3136 -2331 3170 -2315
rect 3256 -1339 3290 -1323
rect 3256 -2331 3290 -2315
rect 3514 -1339 3548 -1323
rect 3514 -2331 3548 -2315
rect 3634 -1339 3668 -1323
rect 3634 -2331 3668 -2315
rect 3892 -1339 3926 -1323
rect 3892 -2331 3926 -2315
rect 4012 -1339 4046 -1323
rect 4012 -2331 4046 -2315
rect 4270 -1339 4304 -1323
rect 4270 -2331 4304 -2315
rect 4390 -1339 4424 -1323
rect 4390 -2331 4424 -2315
rect 4648 -1339 4682 -1323
rect 4648 -2331 4682 -2315
rect -4636 -2399 -4620 -2365
rect -4452 -2399 -4436 -2365
rect -4258 -2399 -4242 -2365
rect -4074 -2399 -4058 -2365
rect -3880 -2399 -3864 -2365
rect -3696 -2399 -3680 -2365
rect -3502 -2399 -3486 -2365
rect -3318 -2399 -3302 -2365
rect -3124 -2399 -3108 -2365
rect -2940 -2399 -2924 -2365
rect -2746 -2399 -2730 -2365
rect -2562 -2399 -2546 -2365
rect -2368 -2399 -2352 -2365
rect -2184 -2399 -2168 -2365
rect -1990 -2399 -1974 -2365
rect -1806 -2399 -1790 -2365
rect -1612 -2399 -1596 -2365
rect -1428 -2399 -1412 -2365
rect -1234 -2399 -1218 -2365
rect -1050 -2399 -1034 -2365
rect -856 -2399 -840 -2365
rect -672 -2399 -656 -2365
rect -478 -2399 -462 -2365
rect -294 -2399 -278 -2365
rect -100 -2399 -84 -2365
rect 84 -2399 100 -2365
rect 278 -2399 294 -2365
rect 462 -2399 478 -2365
rect 656 -2399 672 -2365
rect 840 -2399 856 -2365
rect 1034 -2399 1050 -2365
rect 1218 -2399 1234 -2365
rect 1412 -2399 1428 -2365
rect 1596 -2399 1612 -2365
rect 1790 -2399 1806 -2365
rect 1974 -2399 1990 -2365
rect 2168 -2399 2184 -2365
rect 2352 -2399 2368 -2365
rect 2546 -2399 2562 -2365
rect 2730 -2399 2746 -2365
rect 2924 -2399 2940 -2365
rect 3108 -2399 3124 -2365
rect 3302 -2399 3318 -2365
rect 3486 -2399 3502 -2365
rect 3680 -2399 3696 -2365
rect 3864 -2399 3880 -2365
rect 4058 -2399 4074 -2365
rect 4242 -2399 4258 -2365
rect 4436 -2399 4452 -2365
rect 4620 -2399 4636 -2365
rect -4816 -2503 -4782 -2441
rect 4782 -2503 4816 -2441
rect -4816 -2537 -4720 -2503
rect 4720 -2537 4816 -2503
<< viali >>
rect -4620 2365 -4452 2399
rect -4242 2365 -4074 2399
rect -3864 2365 -3696 2399
rect -3486 2365 -3318 2399
rect -3108 2365 -2940 2399
rect -2730 2365 -2562 2399
rect -2352 2365 -2184 2399
rect -1974 2365 -1806 2399
rect -1596 2365 -1428 2399
rect -1218 2365 -1050 2399
rect -840 2365 -672 2399
rect -462 2365 -294 2399
rect -84 2365 84 2399
rect 294 2365 462 2399
rect 672 2365 840 2399
rect 1050 2365 1218 2399
rect 1428 2365 1596 2399
rect 1806 2365 1974 2399
rect 2184 2365 2352 2399
rect 2562 2365 2730 2399
rect 2940 2365 3108 2399
rect 3318 2365 3486 2399
rect 3696 2365 3864 2399
rect 4074 2365 4242 2399
rect 4452 2365 4620 2399
rect -4682 1339 -4648 2315
rect -4424 1339 -4390 2315
rect -4304 1339 -4270 2315
rect -4046 1339 -4012 2315
rect -3926 1339 -3892 2315
rect -3668 1339 -3634 2315
rect -3548 1339 -3514 2315
rect -3290 1339 -3256 2315
rect -3170 1339 -3136 2315
rect -2912 1339 -2878 2315
rect -2792 1339 -2758 2315
rect -2534 1339 -2500 2315
rect -2414 1339 -2380 2315
rect -2156 1339 -2122 2315
rect -2036 1339 -2002 2315
rect -1778 1339 -1744 2315
rect -1658 1339 -1624 2315
rect -1400 1339 -1366 2315
rect -1280 1339 -1246 2315
rect -1022 1339 -988 2315
rect -902 1339 -868 2315
rect -644 1339 -610 2315
rect -524 1339 -490 2315
rect -266 1339 -232 2315
rect -146 1339 -112 2315
rect 112 1339 146 2315
rect 232 1339 266 2315
rect 490 1339 524 2315
rect 610 1339 644 2315
rect 868 1339 902 2315
rect 988 1339 1022 2315
rect 1246 1339 1280 2315
rect 1366 1339 1400 2315
rect 1624 1339 1658 2315
rect 1744 1339 1778 2315
rect 2002 1339 2036 2315
rect 2122 1339 2156 2315
rect 2380 1339 2414 2315
rect 2500 1339 2534 2315
rect 2758 1339 2792 2315
rect 2878 1339 2912 2315
rect 3136 1339 3170 2315
rect 3256 1339 3290 2315
rect 3514 1339 3548 2315
rect 3634 1339 3668 2315
rect 3892 1339 3926 2315
rect 4012 1339 4046 2315
rect 4270 1339 4304 2315
rect 4390 1339 4424 2315
rect 4648 1339 4682 2315
rect -4620 1255 -4452 1289
rect -4242 1255 -4074 1289
rect -3864 1255 -3696 1289
rect -3486 1255 -3318 1289
rect -3108 1255 -2940 1289
rect -2730 1255 -2562 1289
rect -2352 1255 -2184 1289
rect -1974 1255 -1806 1289
rect -1596 1255 -1428 1289
rect -1218 1255 -1050 1289
rect -840 1255 -672 1289
rect -462 1255 -294 1289
rect -84 1255 84 1289
rect 294 1255 462 1289
rect 672 1255 840 1289
rect 1050 1255 1218 1289
rect 1428 1255 1596 1289
rect 1806 1255 1974 1289
rect 2184 1255 2352 1289
rect 2562 1255 2730 1289
rect 2940 1255 3108 1289
rect 3318 1255 3486 1289
rect 3696 1255 3864 1289
rect 4074 1255 4242 1289
rect 4452 1255 4620 1289
rect -4620 1147 -4452 1181
rect -4242 1147 -4074 1181
rect -3864 1147 -3696 1181
rect -3486 1147 -3318 1181
rect -3108 1147 -2940 1181
rect -2730 1147 -2562 1181
rect -2352 1147 -2184 1181
rect -1974 1147 -1806 1181
rect -1596 1147 -1428 1181
rect -1218 1147 -1050 1181
rect -840 1147 -672 1181
rect -462 1147 -294 1181
rect -84 1147 84 1181
rect 294 1147 462 1181
rect 672 1147 840 1181
rect 1050 1147 1218 1181
rect 1428 1147 1596 1181
rect 1806 1147 1974 1181
rect 2184 1147 2352 1181
rect 2562 1147 2730 1181
rect 2940 1147 3108 1181
rect 3318 1147 3486 1181
rect 3696 1147 3864 1181
rect 4074 1147 4242 1181
rect 4452 1147 4620 1181
rect -4682 121 -4648 1097
rect -4424 121 -4390 1097
rect -4304 121 -4270 1097
rect -4046 121 -4012 1097
rect -3926 121 -3892 1097
rect -3668 121 -3634 1097
rect -3548 121 -3514 1097
rect -3290 121 -3256 1097
rect -3170 121 -3136 1097
rect -2912 121 -2878 1097
rect -2792 121 -2758 1097
rect -2534 121 -2500 1097
rect -2414 121 -2380 1097
rect -2156 121 -2122 1097
rect -2036 121 -2002 1097
rect -1778 121 -1744 1097
rect -1658 121 -1624 1097
rect -1400 121 -1366 1097
rect -1280 121 -1246 1097
rect -1022 121 -988 1097
rect -902 121 -868 1097
rect -644 121 -610 1097
rect -524 121 -490 1097
rect -266 121 -232 1097
rect -146 121 -112 1097
rect 112 121 146 1097
rect 232 121 266 1097
rect 490 121 524 1097
rect 610 121 644 1097
rect 868 121 902 1097
rect 988 121 1022 1097
rect 1246 121 1280 1097
rect 1366 121 1400 1097
rect 1624 121 1658 1097
rect 1744 121 1778 1097
rect 2002 121 2036 1097
rect 2122 121 2156 1097
rect 2380 121 2414 1097
rect 2500 121 2534 1097
rect 2758 121 2792 1097
rect 2878 121 2912 1097
rect 3136 121 3170 1097
rect 3256 121 3290 1097
rect 3514 121 3548 1097
rect 3634 121 3668 1097
rect 3892 121 3926 1097
rect 4012 121 4046 1097
rect 4270 121 4304 1097
rect 4390 121 4424 1097
rect 4648 121 4682 1097
rect -4620 37 -4452 71
rect -4242 37 -4074 71
rect -3864 37 -3696 71
rect -3486 37 -3318 71
rect -3108 37 -2940 71
rect -2730 37 -2562 71
rect -2352 37 -2184 71
rect -1974 37 -1806 71
rect -1596 37 -1428 71
rect -1218 37 -1050 71
rect -840 37 -672 71
rect -462 37 -294 71
rect -84 37 84 71
rect 294 37 462 71
rect 672 37 840 71
rect 1050 37 1218 71
rect 1428 37 1596 71
rect 1806 37 1974 71
rect 2184 37 2352 71
rect 2562 37 2730 71
rect 2940 37 3108 71
rect 3318 37 3486 71
rect 3696 37 3864 71
rect 4074 37 4242 71
rect 4452 37 4620 71
rect -4620 -71 -4452 -37
rect -4242 -71 -4074 -37
rect -3864 -71 -3696 -37
rect -3486 -71 -3318 -37
rect -3108 -71 -2940 -37
rect -2730 -71 -2562 -37
rect -2352 -71 -2184 -37
rect -1974 -71 -1806 -37
rect -1596 -71 -1428 -37
rect -1218 -71 -1050 -37
rect -840 -71 -672 -37
rect -462 -71 -294 -37
rect -84 -71 84 -37
rect 294 -71 462 -37
rect 672 -71 840 -37
rect 1050 -71 1218 -37
rect 1428 -71 1596 -37
rect 1806 -71 1974 -37
rect 2184 -71 2352 -37
rect 2562 -71 2730 -37
rect 2940 -71 3108 -37
rect 3318 -71 3486 -37
rect 3696 -71 3864 -37
rect 4074 -71 4242 -37
rect 4452 -71 4620 -37
rect -4682 -1097 -4648 -121
rect -4424 -1097 -4390 -121
rect -4304 -1097 -4270 -121
rect -4046 -1097 -4012 -121
rect -3926 -1097 -3892 -121
rect -3668 -1097 -3634 -121
rect -3548 -1097 -3514 -121
rect -3290 -1097 -3256 -121
rect -3170 -1097 -3136 -121
rect -2912 -1097 -2878 -121
rect -2792 -1097 -2758 -121
rect -2534 -1097 -2500 -121
rect -2414 -1097 -2380 -121
rect -2156 -1097 -2122 -121
rect -2036 -1097 -2002 -121
rect -1778 -1097 -1744 -121
rect -1658 -1097 -1624 -121
rect -1400 -1097 -1366 -121
rect -1280 -1097 -1246 -121
rect -1022 -1097 -988 -121
rect -902 -1097 -868 -121
rect -644 -1097 -610 -121
rect -524 -1097 -490 -121
rect -266 -1097 -232 -121
rect -146 -1097 -112 -121
rect 112 -1097 146 -121
rect 232 -1097 266 -121
rect 490 -1097 524 -121
rect 610 -1097 644 -121
rect 868 -1097 902 -121
rect 988 -1097 1022 -121
rect 1246 -1097 1280 -121
rect 1366 -1097 1400 -121
rect 1624 -1097 1658 -121
rect 1744 -1097 1778 -121
rect 2002 -1097 2036 -121
rect 2122 -1097 2156 -121
rect 2380 -1097 2414 -121
rect 2500 -1097 2534 -121
rect 2758 -1097 2792 -121
rect 2878 -1097 2912 -121
rect 3136 -1097 3170 -121
rect 3256 -1097 3290 -121
rect 3514 -1097 3548 -121
rect 3634 -1097 3668 -121
rect 3892 -1097 3926 -121
rect 4012 -1097 4046 -121
rect 4270 -1097 4304 -121
rect 4390 -1097 4424 -121
rect 4648 -1097 4682 -121
rect -4620 -1181 -4452 -1147
rect -4242 -1181 -4074 -1147
rect -3864 -1181 -3696 -1147
rect -3486 -1181 -3318 -1147
rect -3108 -1181 -2940 -1147
rect -2730 -1181 -2562 -1147
rect -2352 -1181 -2184 -1147
rect -1974 -1181 -1806 -1147
rect -1596 -1181 -1428 -1147
rect -1218 -1181 -1050 -1147
rect -840 -1181 -672 -1147
rect -462 -1181 -294 -1147
rect -84 -1181 84 -1147
rect 294 -1181 462 -1147
rect 672 -1181 840 -1147
rect 1050 -1181 1218 -1147
rect 1428 -1181 1596 -1147
rect 1806 -1181 1974 -1147
rect 2184 -1181 2352 -1147
rect 2562 -1181 2730 -1147
rect 2940 -1181 3108 -1147
rect 3318 -1181 3486 -1147
rect 3696 -1181 3864 -1147
rect 4074 -1181 4242 -1147
rect 4452 -1181 4620 -1147
rect -4620 -1289 -4452 -1255
rect -4242 -1289 -4074 -1255
rect -3864 -1289 -3696 -1255
rect -3486 -1289 -3318 -1255
rect -3108 -1289 -2940 -1255
rect -2730 -1289 -2562 -1255
rect -2352 -1289 -2184 -1255
rect -1974 -1289 -1806 -1255
rect -1596 -1289 -1428 -1255
rect -1218 -1289 -1050 -1255
rect -840 -1289 -672 -1255
rect -462 -1289 -294 -1255
rect -84 -1289 84 -1255
rect 294 -1289 462 -1255
rect 672 -1289 840 -1255
rect 1050 -1289 1218 -1255
rect 1428 -1289 1596 -1255
rect 1806 -1289 1974 -1255
rect 2184 -1289 2352 -1255
rect 2562 -1289 2730 -1255
rect 2940 -1289 3108 -1255
rect 3318 -1289 3486 -1255
rect 3696 -1289 3864 -1255
rect 4074 -1289 4242 -1255
rect 4452 -1289 4620 -1255
rect -4682 -2315 -4648 -1339
rect -4424 -2315 -4390 -1339
rect -4304 -2315 -4270 -1339
rect -4046 -2315 -4012 -1339
rect -3926 -2315 -3892 -1339
rect -3668 -2315 -3634 -1339
rect -3548 -2315 -3514 -1339
rect -3290 -2315 -3256 -1339
rect -3170 -2315 -3136 -1339
rect -2912 -2315 -2878 -1339
rect -2792 -2315 -2758 -1339
rect -2534 -2315 -2500 -1339
rect -2414 -2315 -2380 -1339
rect -2156 -2315 -2122 -1339
rect -2036 -2315 -2002 -1339
rect -1778 -2315 -1744 -1339
rect -1658 -2315 -1624 -1339
rect -1400 -2315 -1366 -1339
rect -1280 -2315 -1246 -1339
rect -1022 -2315 -988 -1339
rect -902 -2315 -868 -1339
rect -644 -2315 -610 -1339
rect -524 -2315 -490 -1339
rect -266 -2315 -232 -1339
rect -146 -2315 -112 -1339
rect 112 -2315 146 -1339
rect 232 -2315 266 -1339
rect 490 -2315 524 -1339
rect 610 -2315 644 -1339
rect 868 -2315 902 -1339
rect 988 -2315 1022 -1339
rect 1246 -2315 1280 -1339
rect 1366 -2315 1400 -1339
rect 1624 -2315 1658 -1339
rect 1744 -2315 1778 -1339
rect 2002 -2315 2036 -1339
rect 2122 -2315 2156 -1339
rect 2380 -2315 2414 -1339
rect 2500 -2315 2534 -1339
rect 2758 -2315 2792 -1339
rect 2878 -2315 2912 -1339
rect 3136 -2315 3170 -1339
rect 3256 -2315 3290 -1339
rect 3514 -2315 3548 -1339
rect 3634 -2315 3668 -1339
rect 3892 -2315 3926 -1339
rect 4012 -2315 4046 -1339
rect 4270 -2315 4304 -1339
rect 4390 -2315 4424 -1339
rect 4648 -2315 4682 -1339
rect -4620 -2399 -4452 -2365
rect -4242 -2399 -4074 -2365
rect -3864 -2399 -3696 -2365
rect -3486 -2399 -3318 -2365
rect -3108 -2399 -2940 -2365
rect -2730 -2399 -2562 -2365
rect -2352 -2399 -2184 -2365
rect -1974 -2399 -1806 -2365
rect -1596 -2399 -1428 -2365
rect -1218 -2399 -1050 -2365
rect -840 -2399 -672 -2365
rect -462 -2399 -294 -2365
rect -84 -2399 84 -2365
rect 294 -2399 462 -2365
rect 672 -2399 840 -2365
rect 1050 -2399 1218 -2365
rect 1428 -2399 1596 -2365
rect 1806 -2399 1974 -2365
rect 2184 -2399 2352 -2365
rect 2562 -2399 2730 -2365
rect 2940 -2399 3108 -2365
rect 3318 -2399 3486 -2365
rect 3696 -2399 3864 -2365
rect 4074 -2399 4242 -2365
rect 4452 -2399 4620 -2365
<< metal1 >>
rect -4632 2399 -4440 2405
rect -4632 2365 -4620 2399
rect -4452 2365 -4440 2399
rect -4632 2359 -4440 2365
rect -4254 2399 -4062 2405
rect -4254 2365 -4242 2399
rect -4074 2365 -4062 2399
rect -4254 2359 -4062 2365
rect -3876 2399 -3684 2405
rect -3876 2365 -3864 2399
rect -3696 2365 -3684 2399
rect -3876 2359 -3684 2365
rect -3498 2399 -3306 2405
rect -3498 2365 -3486 2399
rect -3318 2365 -3306 2399
rect -3498 2359 -3306 2365
rect -3120 2399 -2928 2405
rect -3120 2365 -3108 2399
rect -2940 2365 -2928 2399
rect -3120 2359 -2928 2365
rect -2742 2399 -2550 2405
rect -2742 2365 -2730 2399
rect -2562 2365 -2550 2399
rect -2742 2359 -2550 2365
rect -2364 2399 -2172 2405
rect -2364 2365 -2352 2399
rect -2184 2365 -2172 2399
rect -2364 2359 -2172 2365
rect -1986 2399 -1794 2405
rect -1986 2365 -1974 2399
rect -1806 2365 -1794 2399
rect -1986 2359 -1794 2365
rect -1608 2399 -1416 2405
rect -1608 2365 -1596 2399
rect -1428 2365 -1416 2399
rect -1608 2359 -1416 2365
rect -1230 2399 -1038 2405
rect -1230 2365 -1218 2399
rect -1050 2365 -1038 2399
rect -1230 2359 -1038 2365
rect -852 2399 -660 2405
rect -852 2365 -840 2399
rect -672 2365 -660 2399
rect -852 2359 -660 2365
rect -474 2399 -282 2405
rect -474 2365 -462 2399
rect -294 2365 -282 2399
rect -474 2359 -282 2365
rect -96 2399 96 2405
rect -96 2365 -84 2399
rect 84 2365 96 2399
rect -96 2359 96 2365
rect 282 2399 474 2405
rect 282 2365 294 2399
rect 462 2365 474 2399
rect 282 2359 474 2365
rect 660 2399 852 2405
rect 660 2365 672 2399
rect 840 2365 852 2399
rect 660 2359 852 2365
rect 1038 2399 1230 2405
rect 1038 2365 1050 2399
rect 1218 2365 1230 2399
rect 1038 2359 1230 2365
rect 1416 2399 1608 2405
rect 1416 2365 1428 2399
rect 1596 2365 1608 2399
rect 1416 2359 1608 2365
rect 1794 2399 1986 2405
rect 1794 2365 1806 2399
rect 1974 2365 1986 2399
rect 1794 2359 1986 2365
rect 2172 2399 2364 2405
rect 2172 2365 2184 2399
rect 2352 2365 2364 2399
rect 2172 2359 2364 2365
rect 2550 2399 2742 2405
rect 2550 2365 2562 2399
rect 2730 2365 2742 2399
rect 2550 2359 2742 2365
rect 2928 2399 3120 2405
rect 2928 2365 2940 2399
rect 3108 2365 3120 2399
rect 2928 2359 3120 2365
rect 3306 2399 3498 2405
rect 3306 2365 3318 2399
rect 3486 2365 3498 2399
rect 3306 2359 3498 2365
rect 3684 2399 3876 2405
rect 3684 2365 3696 2399
rect 3864 2365 3876 2399
rect 3684 2359 3876 2365
rect 4062 2399 4254 2405
rect 4062 2365 4074 2399
rect 4242 2365 4254 2399
rect 4062 2359 4254 2365
rect 4440 2399 4632 2405
rect 4440 2365 4452 2399
rect 4620 2365 4632 2399
rect 4440 2359 4632 2365
rect -4688 2315 -4642 2327
rect -4688 1339 -4682 2315
rect -4648 1339 -4642 2315
rect -4688 1327 -4642 1339
rect -4430 2315 -4384 2327
rect -4430 1339 -4424 2315
rect -4390 1339 -4384 2315
rect -4430 1327 -4384 1339
rect -4310 2315 -4264 2327
rect -4310 1339 -4304 2315
rect -4270 1339 -4264 2315
rect -4310 1327 -4264 1339
rect -4052 2315 -4006 2327
rect -4052 1339 -4046 2315
rect -4012 1339 -4006 2315
rect -4052 1327 -4006 1339
rect -3932 2315 -3886 2327
rect -3932 1339 -3926 2315
rect -3892 1339 -3886 2315
rect -3932 1327 -3886 1339
rect -3674 2315 -3628 2327
rect -3674 1339 -3668 2315
rect -3634 1339 -3628 2315
rect -3674 1327 -3628 1339
rect -3554 2315 -3508 2327
rect -3554 1339 -3548 2315
rect -3514 1339 -3508 2315
rect -3554 1327 -3508 1339
rect -3296 2315 -3250 2327
rect -3296 1339 -3290 2315
rect -3256 1339 -3250 2315
rect -3296 1327 -3250 1339
rect -3176 2315 -3130 2327
rect -3176 1339 -3170 2315
rect -3136 1339 -3130 2315
rect -3176 1327 -3130 1339
rect -2918 2315 -2872 2327
rect -2918 1339 -2912 2315
rect -2878 1339 -2872 2315
rect -2918 1327 -2872 1339
rect -2798 2315 -2752 2327
rect -2798 1339 -2792 2315
rect -2758 1339 -2752 2315
rect -2798 1327 -2752 1339
rect -2540 2315 -2494 2327
rect -2540 1339 -2534 2315
rect -2500 1339 -2494 2315
rect -2540 1327 -2494 1339
rect -2420 2315 -2374 2327
rect -2420 1339 -2414 2315
rect -2380 1339 -2374 2315
rect -2420 1327 -2374 1339
rect -2162 2315 -2116 2327
rect -2162 1339 -2156 2315
rect -2122 1339 -2116 2315
rect -2162 1327 -2116 1339
rect -2042 2315 -1996 2327
rect -2042 1339 -2036 2315
rect -2002 1339 -1996 2315
rect -2042 1327 -1996 1339
rect -1784 2315 -1738 2327
rect -1784 1339 -1778 2315
rect -1744 1339 -1738 2315
rect -1784 1327 -1738 1339
rect -1664 2315 -1618 2327
rect -1664 1339 -1658 2315
rect -1624 1339 -1618 2315
rect -1664 1327 -1618 1339
rect -1406 2315 -1360 2327
rect -1406 1339 -1400 2315
rect -1366 1339 -1360 2315
rect -1406 1327 -1360 1339
rect -1286 2315 -1240 2327
rect -1286 1339 -1280 2315
rect -1246 1339 -1240 2315
rect -1286 1327 -1240 1339
rect -1028 2315 -982 2327
rect -1028 1339 -1022 2315
rect -988 1339 -982 2315
rect -1028 1327 -982 1339
rect -908 2315 -862 2327
rect -908 1339 -902 2315
rect -868 1339 -862 2315
rect -908 1327 -862 1339
rect -650 2315 -604 2327
rect -650 1339 -644 2315
rect -610 1339 -604 2315
rect -650 1327 -604 1339
rect -530 2315 -484 2327
rect -530 1339 -524 2315
rect -490 1339 -484 2315
rect -530 1327 -484 1339
rect -272 2315 -226 2327
rect -272 1339 -266 2315
rect -232 1339 -226 2315
rect -272 1327 -226 1339
rect -152 2315 -106 2327
rect -152 1339 -146 2315
rect -112 1339 -106 2315
rect -152 1327 -106 1339
rect 106 2315 152 2327
rect 106 1339 112 2315
rect 146 1339 152 2315
rect 106 1327 152 1339
rect 226 2315 272 2327
rect 226 1339 232 2315
rect 266 1339 272 2315
rect 226 1327 272 1339
rect 484 2315 530 2327
rect 484 1339 490 2315
rect 524 1339 530 2315
rect 484 1327 530 1339
rect 604 2315 650 2327
rect 604 1339 610 2315
rect 644 1339 650 2315
rect 604 1327 650 1339
rect 862 2315 908 2327
rect 862 1339 868 2315
rect 902 1339 908 2315
rect 862 1327 908 1339
rect 982 2315 1028 2327
rect 982 1339 988 2315
rect 1022 1339 1028 2315
rect 982 1327 1028 1339
rect 1240 2315 1286 2327
rect 1240 1339 1246 2315
rect 1280 1339 1286 2315
rect 1240 1327 1286 1339
rect 1360 2315 1406 2327
rect 1360 1339 1366 2315
rect 1400 1339 1406 2315
rect 1360 1327 1406 1339
rect 1618 2315 1664 2327
rect 1618 1339 1624 2315
rect 1658 1339 1664 2315
rect 1618 1327 1664 1339
rect 1738 2315 1784 2327
rect 1738 1339 1744 2315
rect 1778 1339 1784 2315
rect 1738 1327 1784 1339
rect 1996 2315 2042 2327
rect 1996 1339 2002 2315
rect 2036 1339 2042 2315
rect 1996 1327 2042 1339
rect 2116 2315 2162 2327
rect 2116 1339 2122 2315
rect 2156 1339 2162 2315
rect 2116 1327 2162 1339
rect 2374 2315 2420 2327
rect 2374 1339 2380 2315
rect 2414 1339 2420 2315
rect 2374 1327 2420 1339
rect 2494 2315 2540 2327
rect 2494 1339 2500 2315
rect 2534 1339 2540 2315
rect 2494 1327 2540 1339
rect 2752 2315 2798 2327
rect 2752 1339 2758 2315
rect 2792 1339 2798 2315
rect 2752 1327 2798 1339
rect 2872 2315 2918 2327
rect 2872 1339 2878 2315
rect 2912 1339 2918 2315
rect 2872 1327 2918 1339
rect 3130 2315 3176 2327
rect 3130 1339 3136 2315
rect 3170 1339 3176 2315
rect 3130 1327 3176 1339
rect 3250 2315 3296 2327
rect 3250 1339 3256 2315
rect 3290 1339 3296 2315
rect 3250 1327 3296 1339
rect 3508 2315 3554 2327
rect 3508 1339 3514 2315
rect 3548 1339 3554 2315
rect 3508 1327 3554 1339
rect 3628 2315 3674 2327
rect 3628 1339 3634 2315
rect 3668 1339 3674 2315
rect 3628 1327 3674 1339
rect 3886 2315 3932 2327
rect 3886 1339 3892 2315
rect 3926 1339 3932 2315
rect 3886 1327 3932 1339
rect 4006 2315 4052 2327
rect 4006 1339 4012 2315
rect 4046 1339 4052 2315
rect 4006 1327 4052 1339
rect 4264 2315 4310 2327
rect 4264 1339 4270 2315
rect 4304 1339 4310 2315
rect 4264 1327 4310 1339
rect 4384 2315 4430 2327
rect 4384 1339 4390 2315
rect 4424 1339 4430 2315
rect 4384 1327 4430 1339
rect 4642 2315 4688 2327
rect 4642 1339 4648 2315
rect 4682 1339 4688 2315
rect 4642 1327 4688 1339
rect -4632 1289 -4440 1295
rect -4632 1255 -4620 1289
rect -4452 1255 -4440 1289
rect -4632 1249 -4440 1255
rect -4254 1289 -4062 1295
rect -4254 1255 -4242 1289
rect -4074 1255 -4062 1289
rect -4254 1249 -4062 1255
rect -3876 1289 -3684 1295
rect -3876 1255 -3864 1289
rect -3696 1255 -3684 1289
rect -3876 1249 -3684 1255
rect -3498 1289 -3306 1295
rect -3498 1255 -3486 1289
rect -3318 1255 -3306 1289
rect -3498 1249 -3306 1255
rect -3120 1289 -2928 1295
rect -3120 1255 -3108 1289
rect -2940 1255 -2928 1289
rect -3120 1249 -2928 1255
rect -2742 1289 -2550 1295
rect -2742 1255 -2730 1289
rect -2562 1255 -2550 1289
rect -2742 1249 -2550 1255
rect -2364 1289 -2172 1295
rect -2364 1255 -2352 1289
rect -2184 1255 -2172 1289
rect -2364 1249 -2172 1255
rect -1986 1289 -1794 1295
rect -1986 1255 -1974 1289
rect -1806 1255 -1794 1289
rect -1986 1249 -1794 1255
rect -1608 1289 -1416 1295
rect -1608 1255 -1596 1289
rect -1428 1255 -1416 1289
rect -1608 1249 -1416 1255
rect -1230 1289 -1038 1295
rect -1230 1255 -1218 1289
rect -1050 1255 -1038 1289
rect -1230 1249 -1038 1255
rect -852 1289 -660 1295
rect -852 1255 -840 1289
rect -672 1255 -660 1289
rect -852 1249 -660 1255
rect -474 1289 -282 1295
rect -474 1255 -462 1289
rect -294 1255 -282 1289
rect -474 1249 -282 1255
rect -96 1289 96 1295
rect -96 1255 -84 1289
rect 84 1255 96 1289
rect -96 1249 96 1255
rect 282 1289 474 1295
rect 282 1255 294 1289
rect 462 1255 474 1289
rect 282 1249 474 1255
rect 660 1289 852 1295
rect 660 1255 672 1289
rect 840 1255 852 1289
rect 660 1249 852 1255
rect 1038 1289 1230 1295
rect 1038 1255 1050 1289
rect 1218 1255 1230 1289
rect 1038 1249 1230 1255
rect 1416 1289 1608 1295
rect 1416 1255 1428 1289
rect 1596 1255 1608 1289
rect 1416 1249 1608 1255
rect 1794 1289 1986 1295
rect 1794 1255 1806 1289
rect 1974 1255 1986 1289
rect 1794 1249 1986 1255
rect 2172 1289 2364 1295
rect 2172 1255 2184 1289
rect 2352 1255 2364 1289
rect 2172 1249 2364 1255
rect 2550 1289 2742 1295
rect 2550 1255 2562 1289
rect 2730 1255 2742 1289
rect 2550 1249 2742 1255
rect 2928 1289 3120 1295
rect 2928 1255 2940 1289
rect 3108 1255 3120 1289
rect 2928 1249 3120 1255
rect 3306 1289 3498 1295
rect 3306 1255 3318 1289
rect 3486 1255 3498 1289
rect 3306 1249 3498 1255
rect 3684 1289 3876 1295
rect 3684 1255 3696 1289
rect 3864 1255 3876 1289
rect 3684 1249 3876 1255
rect 4062 1289 4254 1295
rect 4062 1255 4074 1289
rect 4242 1255 4254 1289
rect 4062 1249 4254 1255
rect 4440 1289 4632 1295
rect 4440 1255 4452 1289
rect 4620 1255 4632 1289
rect 4440 1249 4632 1255
rect -4632 1181 -4440 1187
rect -4632 1147 -4620 1181
rect -4452 1147 -4440 1181
rect -4632 1141 -4440 1147
rect -4254 1181 -4062 1187
rect -4254 1147 -4242 1181
rect -4074 1147 -4062 1181
rect -4254 1141 -4062 1147
rect -3876 1181 -3684 1187
rect -3876 1147 -3864 1181
rect -3696 1147 -3684 1181
rect -3876 1141 -3684 1147
rect -3498 1181 -3306 1187
rect -3498 1147 -3486 1181
rect -3318 1147 -3306 1181
rect -3498 1141 -3306 1147
rect -3120 1181 -2928 1187
rect -3120 1147 -3108 1181
rect -2940 1147 -2928 1181
rect -3120 1141 -2928 1147
rect -2742 1181 -2550 1187
rect -2742 1147 -2730 1181
rect -2562 1147 -2550 1181
rect -2742 1141 -2550 1147
rect -2364 1181 -2172 1187
rect -2364 1147 -2352 1181
rect -2184 1147 -2172 1181
rect -2364 1141 -2172 1147
rect -1986 1181 -1794 1187
rect -1986 1147 -1974 1181
rect -1806 1147 -1794 1181
rect -1986 1141 -1794 1147
rect -1608 1181 -1416 1187
rect -1608 1147 -1596 1181
rect -1428 1147 -1416 1181
rect -1608 1141 -1416 1147
rect -1230 1181 -1038 1187
rect -1230 1147 -1218 1181
rect -1050 1147 -1038 1181
rect -1230 1141 -1038 1147
rect -852 1181 -660 1187
rect -852 1147 -840 1181
rect -672 1147 -660 1181
rect -852 1141 -660 1147
rect -474 1181 -282 1187
rect -474 1147 -462 1181
rect -294 1147 -282 1181
rect -474 1141 -282 1147
rect -96 1181 96 1187
rect -96 1147 -84 1181
rect 84 1147 96 1181
rect -96 1141 96 1147
rect 282 1181 474 1187
rect 282 1147 294 1181
rect 462 1147 474 1181
rect 282 1141 474 1147
rect 660 1181 852 1187
rect 660 1147 672 1181
rect 840 1147 852 1181
rect 660 1141 852 1147
rect 1038 1181 1230 1187
rect 1038 1147 1050 1181
rect 1218 1147 1230 1181
rect 1038 1141 1230 1147
rect 1416 1181 1608 1187
rect 1416 1147 1428 1181
rect 1596 1147 1608 1181
rect 1416 1141 1608 1147
rect 1794 1181 1986 1187
rect 1794 1147 1806 1181
rect 1974 1147 1986 1181
rect 1794 1141 1986 1147
rect 2172 1181 2364 1187
rect 2172 1147 2184 1181
rect 2352 1147 2364 1181
rect 2172 1141 2364 1147
rect 2550 1181 2742 1187
rect 2550 1147 2562 1181
rect 2730 1147 2742 1181
rect 2550 1141 2742 1147
rect 2928 1181 3120 1187
rect 2928 1147 2940 1181
rect 3108 1147 3120 1181
rect 2928 1141 3120 1147
rect 3306 1181 3498 1187
rect 3306 1147 3318 1181
rect 3486 1147 3498 1181
rect 3306 1141 3498 1147
rect 3684 1181 3876 1187
rect 3684 1147 3696 1181
rect 3864 1147 3876 1181
rect 3684 1141 3876 1147
rect 4062 1181 4254 1187
rect 4062 1147 4074 1181
rect 4242 1147 4254 1181
rect 4062 1141 4254 1147
rect 4440 1181 4632 1187
rect 4440 1147 4452 1181
rect 4620 1147 4632 1181
rect 4440 1141 4632 1147
rect -4688 1097 -4642 1109
rect -4688 121 -4682 1097
rect -4648 121 -4642 1097
rect -4688 109 -4642 121
rect -4430 1097 -4384 1109
rect -4430 121 -4424 1097
rect -4390 121 -4384 1097
rect -4430 109 -4384 121
rect -4310 1097 -4264 1109
rect -4310 121 -4304 1097
rect -4270 121 -4264 1097
rect -4310 109 -4264 121
rect -4052 1097 -4006 1109
rect -4052 121 -4046 1097
rect -4012 121 -4006 1097
rect -4052 109 -4006 121
rect -3932 1097 -3886 1109
rect -3932 121 -3926 1097
rect -3892 121 -3886 1097
rect -3932 109 -3886 121
rect -3674 1097 -3628 1109
rect -3674 121 -3668 1097
rect -3634 121 -3628 1097
rect -3674 109 -3628 121
rect -3554 1097 -3508 1109
rect -3554 121 -3548 1097
rect -3514 121 -3508 1097
rect -3554 109 -3508 121
rect -3296 1097 -3250 1109
rect -3296 121 -3290 1097
rect -3256 121 -3250 1097
rect -3296 109 -3250 121
rect -3176 1097 -3130 1109
rect -3176 121 -3170 1097
rect -3136 121 -3130 1097
rect -3176 109 -3130 121
rect -2918 1097 -2872 1109
rect -2918 121 -2912 1097
rect -2878 121 -2872 1097
rect -2918 109 -2872 121
rect -2798 1097 -2752 1109
rect -2798 121 -2792 1097
rect -2758 121 -2752 1097
rect -2798 109 -2752 121
rect -2540 1097 -2494 1109
rect -2540 121 -2534 1097
rect -2500 121 -2494 1097
rect -2540 109 -2494 121
rect -2420 1097 -2374 1109
rect -2420 121 -2414 1097
rect -2380 121 -2374 1097
rect -2420 109 -2374 121
rect -2162 1097 -2116 1109
rect -2162 121 -2156 1097
rect -2122 121 -2116 1097
rect -2162 109 -2116 121
rect -2042 1097 -1996 1109
rect -2042 121 -2036 1097
rect -2002 121 -1996 1097
rect -2042 109 -1996 121
rect -1784 1097 -1738 1109
rect -1784 121 -1778 1097
rect -1744 121 -1738 1097
rect -1784 109 -1738 121
rect -1664 1097 -1618 1109
rect -1664 121 -1658 1097
rect -1624 121 -1618 1097
rect -1664 109 -1618 121
rect -1406 1097 -1360 1109
rect -1406 121 -1400 1097
rect -1366 121 -1360 1097
rect -1406 109 -1360 121
rect -1286 1097 -1240 1109
rect -1286 121 -1280 1097
rect -1246 121 -1240 1097
rect -1286 109 -1240 121
rect -1028 1097 -982 1109
rect -1028 121 -1022 1097
rect -988 121 -982 1097
rect -1028 109 -982 121
rect -908 1097 -862 1109
rect -908 121 -902 1097
rect -868 121 -862 1097
rect -908 109 -862 121
rect -650 1097 -604 1109
rect -650 121 -644 1097
rect -610 121 -604 1097
rect -650 109 -604 121
rect -530 1097 -484 1109
rect -530 121 -524 1097
rect -490 121 -484 1097
rect -530 109 -484 121
rect -272 1097 -226 1109
rect -272 121 -266 1097
rect -232 121 -226 1097
rect -272 109 -226 121
rect -152 1097 -106 1109
rect -152 121 -146 1097
rect -112 121 -106 1097
rect -152 109 -106 121
rect 106 1097 152 1109
rect 106 121 112 1097
rect 146 121 152 1097
rect 106 109 152 121
rect 226 1097 272 1109
rect 226 121 232 1097
rect 266 121 272 1097
rect 226 109 272 121
rect 484 1097 530 1109
rect 484 121 490 1097
rect 524 121 530 1097
rect 484 109 530 121
rect 604 1097 650 1109
rect 604 121 610 1097
rect 644 121 650 1097
rect 604 109 650 121
rect 862 1097 908 1109
rect 862 121 868 1097
rect 902 121 908 1097
rect 862 109 908 121
rect 982 1097 1028 1109
rect 982 121 988 1097
rect 1022 121 1028 1097
rect 982 109 1028 121
rect 1240 1097 1286 1109
rect 1240 121 1246 1097
rect 1280 121 1286 1097
rect 1240 109 1286 121
rect 1360 1097 1406 1109
rect 1360 121 1366 1097
rect 1400 121 1406 1097
rect 1360 109 1406 121
rect 1618 1097 1664 1109
rect 1618 121 1624 1097
rect 1658 121 1664 1097
rect 1618 109 1664 121
rect 1738 1097 1784 1109
rect 1738 121 1744 1097
rect 1778 121 1784 1097
rect 1738 109 1784 121
rect 1996 1097 2042 1109
rect 1996 121 2002 1097
rect 2036 121 2042 1097
rect 1996 109 2042 121
rect 2116 1097 2162 1109
rect 2116 121 2122 1097
rect 2156 121 2162 1097
rect 2116 109 2162 121
rect 2374 1097 2420 1109
rect 2374 121 2380 1097
rect 2414 121 2420 1097
rect 2374 109 2420 121
rect 2494 1097 2540 1109
rect 2494 121 2500 1097
rect 2534 121 2540 1097
rect 2494 109 2540 121
rect 2752 1097 2798 1109
rect 2752 121 2758 1097
rect 2792 121 2798 1097
rect 2752 109 2798 121
rect 2872 1097 2918 1109
rect 2872 121 2878 1097
rect 2912 121 2918 1097
rect 2872 109 2918 121
rect 3130 1097 3176 1109
rect 3130 121 3136 1097
rect 3170 121 3176 1097
rect 3130 109 3176 121
rect 3250 1097 3296 1109
rect 3250 121 3256 1097
rect 3290 121 3296 1097
rect 3250 109 3296 121
rect 3508 1097 3554 1109
rect 3508 121 3514 1097
rect 3548 121 3554 1097
rect 3508 109 3554 121
rect 3628 1097 3674 1109
rect 3628 121 3634 1097
rect 3668 121 3674 1097
rect 3628 109 3674 121
rect 3886 1097 3932 1109
rect 3886 121 3892 1097
rect 3926 121 3932 1097
rect 3886 109 3932 121
rect 4006 1097 4052 1109
rect 4006 121 4012 1097
rect 4046 121 4052 1097
rect 4006 109 4052 121
rect 4264 1097 4310 1109
rect 4264 121 4270 1097
rect 4304 121 4310 1097
rect 4264 109 4310 121
rect 4384 1097 4430 1109
rect 4384 121 4390 1097
rect 4424 121 4430 1097
rect 4384 109 4430 121
rect 4642 1097 4688 1109
rect 4642 121 4648 1097
rect 4682 121 4688 1097
rect 4642 109 4688 121
rect -4632 71 -4440 77
rect -4632 37 -4620 71
rect -4452 37 -4440 71
rect -4632 31 -4440 37
rect -4254 71 -4062 77
rect -4254 37 -4242 71
rect -4074 37 -4062 71
rect -4254 31 -4062 37
rect -3876 71 -3684 77
rect -3876 37 -3864 71
rect -3696 37 -3684 71
rect -3876 31 -3684 37
rect -3498 71 -3306 77
rect -3498 37 -3486 71
rect -3318 37 -3306 71
rect -3498 31 -3306 37
rect -3120 71 -2928 77
rect -3120 37 -3108 71
rect -2940 37 -2928 71
rect -3120 31 -2928 37
rect -2742 71 -2550 77
rect -2742 37 -2730 71
rect -2562 37 -2550 71
rect -2742 31 -2550 37
rect -2364 71 -2172 77
rect -2364 37 -2352 71
rect -2184 37 -2172 71
rect -2364 31 -2172 37
rect -1986 71 -1794 77
rect -1986 37 -1974 71
rect -1806 37 -1794 71
rect -1986 31 -1794 37
rect -1608 71 -1416 77
rect -1608 37 -1596 71
rect -1428 37 -1416 71
rect -1608 31 -1416 37
rect -1230 71 -1038 77
rect -1230 37 -1218 71
rect -1050 37 -1038 71
rect -1230 31 -1038 37
rect -852 71 -660 77
rect -852 37 -840 71
rect -672 37 -660 71
rect -852 31 -660 37
rect -474 71 -282 77
rect -474 37 -462 71
rect -294 37 -282 71
rect -474 31 -282 37
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect 282 71 474 77
rect 282 37 294 71
rect 462 37 474 71
rect 282 31 474 37
rect 660 71 852 77
rect 660 37 672 71
rect 840 37 852 71
rect 660 31 852 37
rect 1038 71 1230 77
rect 1038 37 1050 71
rect 1218 37 1230 71
rect 1038 31 1230 37
rect 1416 71 1608 77
rect 1416 37 1428 71
rect 1596 37 1608 71
rect 1416 31 1608 37
rect 1794 71 1986 77
rect 1794 37 1806 71
rect 1974 37 1986 71
rect 1794 31 1986 37
rect 2172 71 2364 77
rect 2172 37 2184 71
rect 2352 37 2364 71
rect 2172 31 2364 37
rect 2550 71 2742 77
rect 2550 37 2562 71
rect 2730 37 2742 71
rect 2550 31 2742 37
rect 2928 71 3120 77
rect 2928 37 2940 71
rect 3108 37 3120 71
rect 2928 31 3120 37
rect 3306 71 3498 77
rect 3306 37 3318 71
rect 3486 37 3498 71
rect 3306 31 3498 37
rect 3684 71 3876 77
rect 3684 37 3696 71
rect 3864 37 3876 71
rect 3684 31 3876 37
rect 4062 71 4254 77
rect 4062 37 4074 71
rect 4242 37 4254 71
rect 4062 31 4254 37
rect 4440 71 4632 77
rect 4440 37 4452 71
rect 4620 37 4632 71
rect 4440 31 4632 37
rect -4632 -37 -4440 -31
rect -4632 -71 -4620 -37
rect -4452 -71 -4440 -37
rect -4632 -77 -4440 -71
rect -4254 -37 -4062 -31
rect -4254 -71 -4242 -37
rect -4074 -71 -4062 -37
rect -4254 -77 -4062 -71
rect -3876 -37 -3684 -31
rect -3876 -71 -3864 -37
rect -3696 -71 -3684 -37
rect -3876 -77 -3684 -71
rect -3498 -37 -3306 -31
rect -3498 -71 -3486 -37
rect -3318 -71 -3306 -37
rect -3498 -77 -3306 -71
rect -3120 -37 -2928 -31
rect -3120 -71 -3108 -37
rect -2940 -71 -2928 -37
rect -3120 -77 -2928 -71
rect -2742 -37 -2550 -31
rect -2742 -71 -2730 -37
rect -2562 -71 -2550 -37
rect -2742 -77 -2550 -71
rect -2364 -37 -2172 -31
rect -2364 -71 -2352 -37
rect -2184 -71 -2172 -37
rect -2364 -77 -2172 -71
rect -1986 -37 -1794 -31
rect -1986 -71 -1974 -37
rect -1806 -71 -1794 -37
rect -1986 -77 -1794 -71
rect -1608 -37 -1416 -31
rect -1608 -71 -1596 -37
rect -1428 -71 -1416 -37
rect -1608 -77 -1416 -71
rect -1230 -37 -1038 -31
rect -1230 -71 -1218 -37
rect -1050 -71 -1038 -37
rect -1230 -77 -1038 -71
rect -852 -37 -660 -31
rect -852 -71 -840 -37
rect -672 -71 -660 -37
rect -852 -77 -660 -71
rect -474 -37 -282 -31
rect -474 -71 -462 -37
rect -294 -71 -282 -37
rect -474 -77 -282 -71
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect 282 -37 474 -31
rect 282 -71 294 -37
rect 462 -71 474 -37
rect 282 -77 474 -71
rect 660 -37 852 -31
rect 660 -71 672 -37
rect 840 -71 852 -37
rect 660 -77 852 -71
rect 1038 -37 1230 -31
rect 1038 -71 1050 -37
rect 1218 -71 1230 -37
rect 1038 -77 1230 -71
rect 1416 -37 1608 -31
rect 1416 -71 1428 -37
rect 1596 -71 1608 -37
rect 1416 -77 1608 -71
rect 1794 -37 1986 -31
rect 1794 -71 1806 -37
rect 1974 -71 1986 -37
rect 1794 -77 1986 -71
rect 2172 -37 2364 -31
rect 2172 -71 2184 -37
rect 2352 -71 2364 -37
rect 2172 -77 2364 -71
rect 2550 -37 2742 -31
rect 2550 -71 2562 -37
rect 2730 -71 2742 -37
rect 2550 -77 2742 -71
rect 2928 -37 3120 -31
rect 2928 -71 2940 -37
rect 3108 -71 3120 -37
rect 2928 -77 3120 -71
rect 3306 -37 3498 -31
rect 3306 -71 3318 -37
rect 3486 -71 3498 -37
rect 3306 -77 3498 -71
rect 3684 -37 3876 -31
rect 3684 -71 3696 -37
rect 3864 -71 3876 -37
rect 3684 -77 3876 -71
rect 4062 -37 4254 -31
rect 4062 -71 4074 -37
rect 4242 -71 4254 -37
rect 4062 -77 4254 -71
rect 4440 -37 4632 -31
rect 4440 -71 4452 -37
rect 4620 -71 4632 -37
rect 4440 -77 4632 -71
rect -4688 -121 -4642 -109
rect -4688 -1097 -4682 -121
rect -4648 -1097 -4642 -121
rect -4688 -1109 -4642 -1097
rect -4430 -121 -4384 -109
rect -4430 -1097 -4424 -121
rect -4390 -1097 -4384 -121
rect -4430 -1109 -4384 -1097
rect -4310 -121 -4264 -109
rect -4310 -1097 -4304 -121
rect -4270 -1097 -4264 -121
rect -4310 -1109 -4264 -1097
rect -4052 -121 -4006 -109
rect -4052 -1097 -4046 -121
rect -4012 -1097 -4006 -121
rect -4052 -1109 -4006 -1097
rect -3932 -121 -3886 -109
rect -3932 -1097 -3926 -121
rect -3892 -1097 -3886 -121
rect -3932 -1109 -3886 -1097
rect -3674 -121 -3628 -109
rect -3674 -1097 -3668 -121
rect -3634 -1097 -3628 -121
rect -3674 -1109 -3628 -1097
rect -3554 -121 -3508 -109
rect -3554 -1097 -3548 -121
rect -3514 -1097 -3508 -121
rect -3554 -1109 -3508 -1097
rect -3296 -121 -3250 -109
rect -3296 -1097 -3290 -121
rect -3256 -1097 -3250 -121
rect -3296 -1109 -3250 -1097
rect -3176 -121 -3130 -109
rect -3176 -1097 -3170 -121
rect -3136 -1097 -3130 -121
rect -3176 -1109 -3130 -1097
rect -2918 -121 -2872 -109
rect -2918 -1097 -2912 -121
rect -2878 -1097 -2872 -121
rect -2918 -1109 -2872 -1097
rect -2798 -121 -2752 -109
rect -2798 -1097 -2792 -121
rect -2758 -1097 -2752 -121
rect -2798 -1109 -2752 -1097
rect -2540 -121 -2494 -109
rect -2540 -1097 -2534 -121
rect -2500 -1097 -2494 -121
rect -2540 -1109 -2494 -1097
rect -2420 -121 -2374 -109
rect -2420 -1097 -2414 -121
rect -2380 -1097 -2374 -121
rect -2420 -1109 -2374 -1097
rect -2162 -121 -2116 -109
rect -2162 -1097 -2156 -121
rect -2122 -1097 -2116 -121
rect -2162 -1109 -2116 -1097
rect -2042 -121 -1996 -109
rect -2042 -1097 -2036 -121
rect -2002 -1097 -1996 -121
rect -2042 -1109 -1996 -1097
rect -1784 -121 -1738 -109
rect -1784 -1097 -1778 -121
rect -1744 -1097 -1738 -121
rect -1784 -1109 -1738 -1097
rect -1664 -121 -1618 -109
rect -1664 -1097 -1658 -121
rect -1624 -1097 -1618 -121
rect -1664 -1109 -1618 -1097
rect -1406 -121 -1360 -109
rect -1406 -1097 -1400 -121
rect -1366 -1097 -1360 -121
rect -1406 -1109 -1360 -1097
rect -1286 -121 -1240 -109
rect -1286 -1097 -1280 -121
rect -1246 -1097 -1240 -121
rect -1286 -1109 -1240 -1097
rect -1028 -121 -982 -109
rect -1028 -1097 -1022 -121
rect -988 -1097 -982 -121
rect -1028 -1109 -982 -1097
rect -908 -121 -862 -109
rect -908 -1097 -902 -121
rect -868 -1097 -862 -121
rect -908 -1109 -862 -1097
rect -650 -121 -604 -109
rect -650 -1097 -644 -121
rect -610 -1097 -604 -121
rect -650 -1109 -604 -1097
rect -530 -121 -484 -109
rect -530 -1097 -524 -121
rect -490 -1097 -484 -121
rect -530 -1109 -484 -1097
rect -272 -121 -226 -109
rect -272 -1097 -266 -121
rect -232 -1097 -226 -121
rect -272 -1109 -226 -1097
rect -152 -121 -106 -109
rect -152 -1097 -146 -121
rect -112 -1097 -106 -121
rect -152 -1109 -106 -1097
rect 106 -121 152 -109
rect 106 -1097 112 -121
rect 146 -1097 152 -121
rect 106 -1109 152 -1097
rect 226 -121 272 -109
rect 226 -1097 232 -121
rect 266 -1097 272 -121
rect 226 -1109 272 -1097
rect 484 -121 530 -109
rect 484 -1097 490 -121
rect 524 -1097 530 -121
rect 484 -1109 530 -1097
rect 604 -121 650 -109
rect 604 -1097 610 -121
rect 644 -1097 650 -121
rect 604 -1109 650 -1097
rect 862 -121 908 -109
rect 862 -1097 868 -121
rect 902 -1097 908 -121
rect 862 -1109 908 -1097
rect 982 -121 1028 -109
rect 982 -1097 988 -121
rect 1022 -1097 1028 -121
rect 982 -1109 1028 -1097
rect 1240 -121 1286 -109
rect 1240 -1097 1246 -121
rect 1280 -1097 1286 -121
rect 1240 -1109 1286 -1097
rect 1360 -121 1406 -109
rect 1360 -1097 1366 -121
rect 1400 -1097 1406 -121
rect 1360 -1109 1406 -1097
rect 1618 -121 1664 -109
rect 1618 -1097 1624 -121
rect 1658 -1097 1664 -121
rect 1618 -1109 1664 -1097
rect 1738 -121 1784 -109
rect 1738 -1097 1744 -121
rect 1778 -1097 1784 -121
rect 1738 -1109 1784 -1097
rect 1996 -121 2042 -109
rect 1996 -1097 2002 -121
rect 2036 -1097 2042 -121
rect 1996 -1109 2042 -1097
rect 2116 -121 2162 -109
rect 2116 -1097 2122 -121
rect 2156 -1097 2162 -121
rect 2116 -1109 2162 -1097
rect 2374 -121 2420 -109
rect 2374 -1097 2380 -121
rect 2414 -1097 2420 -121
rect 2374 -1109 2420 -1097
rect 2494 -121 2540 -109
rect 2494 -1097 2500 -121
rect 2534 -1097 2540 -121
rect 2494 -1109 2540 -1097
rect 2752 -121 2798 -109
rect 2752 -1097 2758 -121
rect 2792 -1097 2798 -121
rect 2752 -1109 2798 -1097
rect 2872 -121 2918 -109
rect 2872 -1097 2878 -121
rect 2912 -1097 2918 -121
rect 2872 -1109 2918 -1097
rect 3130 -121 3176 -109
rect 3130 -1097 3136 -121
rect 3170 -1097 3176 -121
rect 3130 -1109 3176 -1097
rect 3250 -121 3296 -109
rect 3250 -1097 3256 -121
rect 3290 -1097 3296 -121
rect 3250 -1109 3296 -1097
rect 3508 -121 3554 -109
rect 3508 -1097 3514 -121
rect 3548 -1097 3554 -121
rect 3508 -1109 3554 -1097
rect 3628 -121 3674 -109
rect 3628 -1097 3634 -121
rect 3668 -1097 3674 -121
rect 3628 -1109 3674 -1097
rect 3886 -121 3932 -109
rect 3886 -1097 3892 -121
rect 3926 -1097 3932 -121
rect 3886 -1109 3932 -1097
rect 4006 -121 4052 -109
rect 4006 -1097 4012 -121
rect 4046 -1097 4052 -121
rect 4006 -1109 4052 -1097
rect 4264 -121 4310 -109
rect 4264 -1097 4270 -121
rect 4304 -1097 4310 -121
rect 4264 -1109 4310 -1097
rect 4384 -121 4430 -109
rect 4384 -1097 4390 -121
rect 4424 -1097 4430 -121
rect 4384 -1109 4430 -1097
rect 4642 -121 4688 -109
rect 4642 -1097 4648 -121
rect 4682 -1097 4688 -121
rect 4642 -1109 4688 -1097
rect -4632 -1147 -4440 -1141
rect -4632 -1181 -4620 -1147
rect -4452 -1181 -4440 -1147
rect -4632 -1187 -4440 -1181
rect -4254 -1147 -4062 -1141
rect -4254 -1181 -4242 -1147
rect -4074 -1181 -4062 -1147
rect -4254 -1187 -4062 -1181
rect -3876 -1147 -3684 -1141
rect -3876 -1181 -3864 -1147
rect -3696 -1181 -3684 -1147
rect -3876 -1187 -3684 -1181
rect -3498 -1147 -3306 -1141
rect -3498 -1181 -3486 -1147
rect -3318 -1181 -3306 -1147
rect -3498 -1187 -3306 -1181
rect -3120 -1147 -2928 -1141
rect -3120 -1181 -3108 -1147
rect -2940 -1181 -2928 -1147
rect -3120 -1187 -2928 -1181
rect -2742 -1147 -2550 -1141
rect -2742 -1181 -2730 -1147
rect -2562 -1181 -2550 -1147
rect -2742 -1187 -2550 -1181
rect -2364 -1147 -2172 -1141
rect -2364 -1181 -2352 -1147
rect -2184 -1181 -2172 -1147
rect -2364 -1187 -2172 -1181
rect -1986 -1147 -1794 -1141
rect -1986 -1181 -1974 -1147
rect -1806 -1181 -1794 -1147
rect -1986 -1187 -1794 -1181
rect -1608 -1147 -1416 -1141
rect -1608 -1181 -1596 -1147
rect -1428 -1181 -1416 -1147
rect -1608 -1187 -1416 -1181
rect -1230 -1147 -1038 -1141
rect -1230 -1181 -1218 -1147
rect -1050 -1181 -1038 -1147
rect -1230 -1187 -1038 -1181
rect -852 -1147 -660 -1141
rect -852 -1181 -840 -1147
rect -672 -1181 -660 -1147
rect -852 -1187 -660 -1181
rect -474 -1147 -282 -1141
rect -474 -1181 -462 -1147
rect -294 -1181 -282 -1147
rect -474 -1187 -282 -1181
rect -96 -1147 96 -1141
rect -96 -1181 -84 -1147
rect 84 -1181 96 -1147
rect -96 -1187 96 -1181
rect 282 -1147 474 -1141
rect 282 -1181 294 -1147
rect 462 -1181 474 -1147
rect 282 -1187 474 -1181
rect 660 -1147 852 -1141
rect 660 -1181 672 -1147
rect 840 -1181 852 -1147
rect 660 -1187 852 -1181
rect 1038 -1147 1230 -1141
rect 1038 -1181 1050 -1147
rect 1218 -1181 1230 -1147
rect 1038 -1187 1230 -1181
rect 1416 -1147 1608 -1141
rect 1416 -1181 1428 -1147
rect 1596 -1181 1608 -1147
rect 1416 -1187 1608 -1181
rect 1794 -1147 1986 -1141
rect 1794 -1181 1806 -1147
rect 1974 -1181 1986 -1147
rect 1794 -1187 1986 -1181
rect 2172 -1147 2364 -1141
rect 2172 -1181 2184 -1147
rect 2352 -1181 2364 -1147
rect 2172 -1187 2364 -1181
rect 2550 -1147 2742 -1141
rect 2550 -1181 2562 -1147
rect 2730 -1181 2742 -1147
rect 2550 -1187 2742 -1181
rect 2928 -1147 3120 -1141
rect 2928 -1181 2940 -1147
rect 3108 -1181 3120 -1147
rect 2928 -1187 3120 -1181
rect 3306 -1147 3498 -1141
rect 3306 -1181 3318 -1147
rect 3486 -1181 3498 -1147
rect 3306 -1187 3498 -1181
rect 3684 -1147 3876 -1141
rect 3684 -1181 3696 -1147
rect 3864 -1181 3876 -1147
rect 3684 -1187 3876 -1181
rect 4062 -1147 4254 -1141
rect 4062 -1181 4074 -1147
rect 4242 -1181 4254 -1147
rect 4062 -1187 4254 -1181
rect 4440 -1147 4632 -1141
rect 4440 -1181 4452 -1147
rect 4620 -1181 4632 -1147
rect 4440 -1187 4632 -1181
rect -4632 -1255 -4440 -1249
rect -4632 -1289 -4620 -1255
rect -4452 -1289 -4440 -1255
rect -4632 -1295 -4440 -1289
rect -4254 -1255 -4062 -1249
rect -4254 -1289 -4242 -1255
rect -4074 -1289 -4062 -1255
rect -4254 -1295 -4062 -1289
rect -3876 -1255 -3684 -1249
rect -3876 -1289 -3864 -1255
rect -3696 -1289 -3684 -1255
rect -3876 -1295 -3684 -1289
rect -3498 -1255 -3306 -1249
rect -3498 -1289 -3486 -1255
rect -3318 -1289 -3306 -1255
rect -3498 -1295 -3306 -1289
rect -3120 -1255 -2928 -1249
rect -3120 -1289 -3108 -1255
rect -2940 -1289 -2928 -1255
rect -3120 -1295 -2928 -1289
rect -2742 -1255 -2550 -1249
rect -2742 -1289 -2730 -1255
rect -2562 -1289 -2550 -1255
rect -2742 -1295 -2550 -1289
rect -2364 -1255 -2172 -1249
rect -2364 -1289 -2352 -1255
rect -2184 -1289 -2172 -1255
rect -2364 -1295 -2172 -1289
rect -1986 -1255 -1794 -1249
rect -1986 -1289 -1974 -1255
rect -1806 -1289 -1794 -1255
rect -1986 -1295 -1794 -1289
rect -1608 -1255 -1416 -1249
rect -1608 -1289 -1596 -1255
rect -1428 -1289 -1416 -1255
rect -1608 -1295 -1416 -1289
rect -1230 -1255 -1038 -1249
rect -1230 -1289 -1218 -1255
rect -1050 -1289 -1038 -1255
rect -1230 -1295 -1038 -1289
rect -852 -1255 -660 -1249
rect -852 -1289 -840 -1255
rect -672 -1289 -660 -1255
rect -852 -1295 -660 -1289
rect -474 -1255 -282 -1249
rect -474 -1289 -462 -1255
rect -294 -1289 -282 -1255
rect -474 -1295 -282 -1289
rect -96 -1255 96 -1249
rect -96 -1289 -84 -1255
rect 84 -1289 96 -1255
rect -96 -1295 96 -1289
rect 282 -1255 474 -1249
rect 282 -1289 294 -1255
rect 462 -1289 474 -1255
rect 282 -1295 474 -1289
rect 660 -1255 852 -1249
rect 660 -1289 672 -1255
rect 840 -1289 852 -1255
rect 660 -1295 852 -1289
rect 1038 -1255 1230 -1249
rect 1038 -1289 1050 -1255
rect 1218 -1289 1230 -1255
rect 1038 -1295 1230 -1289
rect 1416 -1255 1608 -1249
rect 1416 -1289 1428 -1255
rect 1596 -1289 1608 -1255
rect 1416 -1295 1608 -1289
rect 1794 -1255 1986 -1249
rect 1794 -1289 1806 -1255
rect 1974 -1289 1986 -1255
rect 1794 -1295 1986 -1289
rect 2172 -1255 2364 -1249
rect 2172 -1289 2184 -1255
rect 2352 -1289 2364 -1255
rect 2172 -1295 2364 -1289
rect 2550 -1255 2742 -1249
rect 2550 -1289 2562 -1255
rect 2730 -1289 2742 -1255
rect 2550 -1295 2742 -1289
rect 2928 -1255 3120 -1249
rect 2928 -1289 2940 -1255
rect 3108 -1289 3120 -1255
rect 2928 -1295 3120 -1289
rect 3306 -1255 3498 -1249
rect 3306 -1289 3318 -1255
rect 3486 -1289 3498 -1255
rect 3306 -1295 3498 -1289
rect 3684 -1255 3876 -1249
rect 3684 -1289 3696 -1255
rect 3864 -1289 3876 -1255
rect 3684 -1295 3876 -1289
rect 4062 -1255 4254 -1249
rect 4062 -1289 4074 -1255
rect 4242 -1289 4254 -1255
rect 4062 -1295 4254 -1289
rect 4440 -1255 4632 -1249
rect 4440 -1289 4452 -1255
rect 4620 -1289 4632 -1255
rect 4440 -1295 4632 -1289
rect -4688 -1339 -4642 -1327
rect -4688 -2315 -4682 -1339
rect -4648 -2315 -4642 -1339
rect -4688 -2327 -4642 -2315
rect -4430 -1339 -4384 -1327
rect -4430 -2315 -4424 -1339
rect -4390 -2315 -4384 -1339
rect -4430 -2327 -4384 -2315
rect -4310 -1339 -4264 -1327
rect -4310 -2315 -4304 -1339
rect -4270 -2315 -4264 -1339
rect -4310 -2327 -4264 -2315
rect -4052 -1339 -4006 -1327
rect -4052 -2315 -4046 -1339
rect -4012 -2315 -4006 -1339
rect -4052 -2327 -4006 -2315
rect -3932 -1339 -3886 -1327
rect -3932 -2315 -3926 -1339
rect -3892 -2315 -3886 -1339
rect -3932 -2327 -3886 -2315
rect -3674 -1339 -3628 -1327
rect -3674 -2315 -3668 -1339
rect -3634 -2315 -3628 -1339
rect -3674 -2327 -3628 -2315
rect -3554 -1339 -3508 -1327
rect -3554 -2315 -3548 -1339
rect -3514 -2315 -3508 -1339
rect -3554 -2327 -3508 -2315
rect -3296 -1339 -3250 -1327
rect -3296 -2315 -3290 -1339
rect -3256 -2315 -3250 -1339
rect -3296 -2327 -3250 -2315
rect -3176 -1339 -3130 -1327
rect -3176 -2315 -3170 -1339
rect -3136 -2315 -3130 -1339
rect -3176 -2327 -3130 -2315
rect -2918 -1339 -2872 -1327
rect -2918 -2315 -2912 -1339
rect -2878 -2315 -2872 -1339
rect -2918 -2327 -2872 -2315
rect -2798 -1339 -2752 -1327
rect -2798 -2315 -2792 -1339
rect -2758 -2315 -2752 -1339
rect -2798 -2327 -2752 -2315
rect -2540 -1339 -2494 -1327
rect -2540 -2315 -2534 -1339
rect -2500 -2315 -2494 -1339
rect -2540 -2327 -2494 -2315
rect -2420 -1339 -2374 -1327
rect -2420 -2315 -2414 -1339
rect -2380 -2315 -2374 -1339
rect -2420 -2327 -2374 -2315
rect -2162 -1339 -2116 -1327
rect -2162 -2315 -2156 -1339
rect -2122 -2315 -2116 -1339
rect -2162 -2327 -2116 -2315
rect -2042 -1339 -1996 -1327
rect -2042 -2315 -2036 -1339
rect -2002 -2315 -1996 -1339
rect -2042 -2327 -1996 -2315
rect -1784 -1339 -1738 -1327
rect -1784 -2315 -1778 -1339
rect -1744 -2315 -1738 -1339
rect -1784 -2327 -1738 -2315
rect -1664 -1339 -1618 -1327
rect -1664 -2315 -1658 -1339
rect -1624 -2315 -1618 -1339
rect -1664 -2327 -1618 -2315
rect -1406 -1339 -1360 -1327
rect -1406 -2315 -1400 -1339
rect -1366 -2315 -1360 -1339
rect -1406 -2327 -1360 -2315
rect -1286 -1339 -1240 -1327
rect -1286 -2315 -1280 -1339
rect -1246 -2315 -1240 -1339
rect -1286 -2327 -1240 -2315
rect -1028 -1339 -982 -1327
rect -1028 -2315 -1022 -1339
rect -988 -2315 -982 -1339
rect -1028 -2327 -982 -2315
rect -908 -1339 -862 -1327
rect -908 -2315 -902 -1339
rect -868 -2315 -862 -1339
rect -908 -2327 -862 -2315
rect -650 -1339 -604 -1327
rect -650 -2315 -644 -1339
rect -610 -2315 -604 -1339
rect -650 -2327 -604 -2315
rect -530 -1339 -484 -1327
rect -530 -2315 -524 -1339
rect -490 -2315 -484 -1339
rect -530 -2327 -484 -2315
rect -272 -1339 -226 -1327
rect -272 -2315 -266 -1339
rect -232 -2315 -226 -1339
rect -272 -2327 -226 -2315
rect -152 -1339 -106 -1327
rect -152 -2315 -146 -1339
rect -112 -2315 -106 -1339
rect -152 -2327 -106 -2315
rect 106 -1339 152 -1327
rect 106 -2315 112 -1339
rect 146 -2315 152 -1339
rect 106 -2327 152 -2315
rect 226 -1339 272 -1327
rect 226 -2315 232 -1339
rect 266 -2315 272 -1339
rect 226 -2327 272 -2315
rect 484 -1339 530 -1327
rect 484 -2315 490 -1339
rect 524 -2315 530 -1339
rect 484 -2327 530 -2315
rect 604 -1339 650 -1327
rect 604 -2315 610 -1339
rect 644 -2315 650 -1339
rect 604 -2327 650 -2315
rect 862 -1339 908 -1327
rect 862 -2315 868 -1339
rect 902 -2315 908 -1339
rect 862 -2327 908 -2315
rect 982 -1339 1028 -1327
rect 982 -2315 988 -1339
rect 1022 -2315 1028 -1339
rect 982 -2327 1028 -2315
rect 1240 -1339 1286 -1327
rect 1240 -2315 1246 -1339
rect 1280 -2315 1286 -1339
rect 1240 -2327 1286 -2315
rect 1360 -1339 1406 -1327
rect 1360 -2315 1366 -1339
rect 1400 -2315 1406 -1339
rect 1360 -2327 1406 -2315
rect 1618 -1339 1664 -1327
rect 1618 -2315 1624 -1339
rect 1658 -2315 1664 -1339
rect 1618 -2327 1664 -2315
rect 1738 -1339 1784 -1327
rect 1738 -2315 1744 -1339
rect 1778 -2315 1784 -1339
rect 1738 -2327 1784 -2315
rect 1996 -1339 2042 -1327
rect 1996 -2315 2002 -1339
rect 2036 -2315 2042 -1339
rect 1996 -2327 2042 -2315
rect 2116 -1339 2162 -1327
rect 2116 -2315 2122 -1339
rect 2156 -2315 2162 -1339
rect 2116 -2327 2162 -2315
rect 2374 -1339 2420 -1327
rect 2374 -2315 2380 -1339
rect 2414 -2315 2420 -1339
rect 2374 -2327 2420 -2315
rect 2494 -1339 2540 -1327
rect 2494 -2315 2500 -1339
rect 2534 -2315 2540 -1339
rect 2494 -2327 2540 -2315
rect 2752 -1339 2798 -1327
rect 2752 -2315 2758 -1339
rect 2792 -2315 2798 -1339
rect 2752 -2327 2798 -2315
rect 2872 -1339 2918 -1327
rect 2872 -2315 2878 -1339
rect 2912 -2315 2918 -1339
rect 2872 -2327 2918 -2315
rect 3130 -1339 3176 -1327
rect 3130 -2315 3136 -1339
rect 3170 -2315 3176 -1339
rect 3130 -2327 3176 -2315
rect 3250 -1339 3296 -1327
rect 3250 -2315 3256 -1339
rect 3290 -2315 3296 -1339
rect 3250 -2327 3296 -2315
rect 3508 -1339 3554 -1327
rect 3508 -2315 3514 -1339
rect 3548 -2315 3554 -1339
rect 3508 -2327 3554 -2315
rect 3628 -1339 3674 -1327
rect 3628 -2315 3634 -1339
rect 3668 -2315 3674 -1339
rect 3628 -2327 3674 -2315
rect 3886 -1339 3932 -1327
rect 3886 -2315 3892 -1339
rect 3926 -2315 3932 -1339
rect 3886 -2327 3932 -2315
rect 4006 -1339 4052 -1327
rect 4006 -2315 4012 -1339
rect 4046 -2315 4052 -1339
rect 4006 -2327 4052 -2315
rect 4264 -1339 4310 -1327
rect 4264 -2315 4270 -1339
rect 4304 -2315 4310 -1339
rect 4264 -2327 4310 -2315
rect 4384 -1339 4430 -1327
rect 4384 -2315 4390 -1339
rect 4424 -2315 4430 -1339
rect 4384 -2327 4430 -2315
rect 4642 -1339 4688 -1327
rect 4642 -2315 4648 -1339
rect 4682 -2315 4688 -1339
rect 4642 -2327 4688 -2315
rect -4632 -2365 -4440 -2359
rect -4632 -2399 -4620 -2365
rect -4452 -2399 -4440 -2365
rect -4632 -2405 -4440 -2399
rect -4254 -2365 -4062 -2359
rect -4254 -2399 -4242 -2365
rect -4074 -2399 -4062 -2365
rect -4254 -2405 -4062 -2399
rect -3876 -2365 -3684 -2359
rect -3876 -2399 -3864 -2365
rect -3696 -2399 -3684 -2365
rect -3876 -2405 -3684 -2399
rect -3498 -2365 -3306 -2359
rect -3498 -2399 -3486 -2365
rect -3318 -2399 -3306 -2365
rect -3498 -2405 -3306 -2399
rect -3120 -2365 -2928 -2359
rect -3120 -2399 -3108 -2365
rect -2940 -2399 -2928 -2365
rect -3120 -2405 -2928 -2399
rect -2742 -2365 -2550 -2359
rect -2742 -2399 -2730 -2365
rect -2562 -2399 -2550 -2365
rect -2742 -2405 -2550 -2399
rect -2364 -2365 -2172 -2359
rect -2364 -2399 -2352 -2365
rect -2184 -2399 -2172 -2365
rect -2364 -2405 -2172 -2399
rect -1986 -2365 -1794 -2359
rect -1986 -2399 -1974 -2365
rect -1806 -2399 -1794 -2365
rect -1986 -2405 -1794 -2399
rect -1608 -2365 -1416 -2359
rect -1608 -2399 -1596 -2365
rect -1428 -2399 -1416 -2365
rect -1608 -2405 -1416 -2399
rect -1230 -2365 -1038 -2359
rect -1230 -2399 -1218 -2365
rect -1050 -2399 -1038 -2365
rect -1230 -2405 -1038 -2399
rect -852 -2365 -660 -2359
rect -852 -2399 -840 -2365
rect -672 -2399 -660 -2365
rect -852 -2405 -660 -2399
rect -474 -2365 -282 -2359
rect -474 -2399 -462 -2365
rect -294 -2399 -282 -2365
rect -474 -2405 -282 -2399
rect -96 -2365 96 -2359
rect -96 -2399 -84 -2365
rect 84 -2399 96 -2365
rect -96 -2405 96 -2399
rect 282 -2365 474 -2359
rect 282 -2399 294 -2365
rect 462 -2399 474 -2365
rect 282 -2405 474 -2399
rect 660 -2365 852 -2359
rect 660 -2399 672 -2365
rect 840 -2399 852 -2365
rect 660 -2405 852 -2399
rect 1038 -2365 1230 -2359
rect 1038 -2399 1050 -2365
rect 1218 -2399 1230 -2365
rect 1038 -2405 1230 -2399
rect 1416 -2365 1608 -2359
rect 1416 -2399 1428 -2365
rect 1596 -2399 1608 -2365
rect 1416 -2405 1608 -2399
rect 1794 -2365 1986 -2359
rect 1794 -2399 1806 -2365
rect 1974 -2399 1986 -2365
rect 1794 -2405 1986 -2399
rect 2172 -2365 2364 -2359
rect 2172 -2399 2184 -2365
rect 2352 -2399 2364 -2365
rect 2172 -2405 2364 -2399
rect 2550 -2365 2742 -2359
rect 2550 -2399 2562 -2365
rect 2730 -2399 2742 -2365
rect 2550 -2405 2742 -2399
rect 2928 -2365 3120 -2359
rect 2928 -2399 2940 -2365
rect 3108 -2399 3120 -2365
rect 2928 -2405 3120 -2399
rect 3306 -2365 3498 -2359
rect 3306 -2399 3318 -2365
rect 3486 -2399 3498 -2365
rect 3306 -2405 3498 -2399
rect 3684 -2365 3876 -2359
rect 3684 -2399 3696 -2365
rect 3864 -2399 3876 -2365
rect 3684 -2405 3876 -2399
rect 4062 -2365 4254 -2359
rect 4062 -2399 4074 -2365
rect 4242 -2399 4254 -2365
rect 4062 -2405 4254 -2399
rect 4440 -2365 4632 -2359
rect 4440 -2399 4452 -2365
rect 4620 -2399 4632 -2365
rect 4440 -2405 4632 -2399
<< properties >>
string FIXED_BBOX -4799 -2520 4799 2520
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 1.0 m 4 nf 25 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
