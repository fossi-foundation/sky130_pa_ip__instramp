magic
tech sky130A
timestamp 1729620069
<< pwell >>
rect -3670 -179 3670 179
<< mvnnmos >>
rect -3556 -50 -3356 50
rect -3268 -50 -3068 50
rect -2980 -50 -2780 50
rect -2692 -50 -2492 50
rect -2404 -50 -2204 50
rect -2116 -50 -1916 50
rect -1828 -50 -1628 50
rect -1540 -50 -1340 50
rect -1252 -50 -1052 50
rect -964 -50 -764 50
rect -676 -50 -476 50
rect -388 -50 -188 50
rect -100 -50 100 50
rect 188 -50 388 50
rect 476 -50 676 50
rect 764 -50 964 50
rect 1052 -50 1252 50
rect 1340 -50 1540 50
rect 1628 -50 1828 50
rect 1916 -50 2116 50
rect 2204 -50 2404 50
rect 2492 -50 2692 50
rect 2780 -50 2980 50
rect 3068 -50 3268 50
rect 3356 -50 3556 50
<< mvndiff >>
rect -3585 44 -3556 50
rect -3585 -44 -3579 44
rect -3562 -44 -3556 44
rect -3585 -50 -3556 -44
rect -3356 44 -3327 50
rect -3356 -44 -3350 44
rect -3333 -44 -3327 44
rect -3356 -50 -3327 -44
rect -3297 44 -3268 50
rect -3297 -44 -3291 44
rect -3274 -44 -3268 44
rect -3297 -50 -3268 -44
rect -3068 44 -3039 50
rect -3068 -44 -3062 44
rect -3045 -44 -3039 44
rect -3068 -50 -3039 -44
rect -3009 44 -2980 50
rect -3009 -44 -3003 44
rect -2986 -44 -2980 44
rect -3009 -50 -2980 -44
rect -2780 44 -2751 50
rect -2780 -44 -2774 44
rect -2757 -44 -2751 44
rect -2780 -50 -2751 -44
rect -2721 44 -2692 50
rect -2721 -44 -2715 44
rect -2698 -44 -2692 44
rect -2721 -50 -2692 -44
rect -2492 44 -2463 50
rect -2492 -44 -2486 44
rect -2469 -44 -2463 44
rect -2492 -50 -2463 -44
rect -2433 44 -2404 50
rect -2433 -44 -2427 44
rect -2410 -44 -2404 44
rect -2433 -50 -2404 -44
rect -2204 44 -2175 50
rect -2204 -44 -2198 44
rect -2181 -44 -2175 44
rect -2204 -50 -2175 -44
rect -2145 44 -2116 50
rect -2145 -44 -2139 44
rect -2122 -44 -2116 44
rect -2145 -50 -2116 -44
rect -1916 44 -1887 50
rect -1916 -44 -1910 44
rect -1893 -44 -1887 44
rect -1916 -50 -1887 -44
rect -1857 44 -1828 50
rect -1857 -44 -1851 44
rect -1834 -44 -1828 44
rect -1857 -50 -1828 -44
rect -1628 44 -1599 50
rect -1628 -44 -1622 44
rect -1605 -44 -1599 44
rect -1628 -50 -1599 -44
rect -1569 44 -1540 50
rect -1569 -44 -1563 44
rect -1546 -44 -1540 44
rect -1569 -50 -1540 -44
rect -1340 44 -1311 50
rect -1340 -44 -1334 44
rect -1317 -44 -1311 44
rect -1340 -50 -1311 -44
rect -1281 44 -1252 50
rect -1281 -44 -1275 44
rect -1258 -44 -1252 44
rect -1281 -50 -1252 -44
rect -1052 44 -1023 50
rect -1052 -44 -1046 44
rect -1029 -44 -1023 44
rect -1052 -50 -1023 -44
rect -993 44 -964 50
rect -993 -44 -987 44
rect -970 -44 -964 44
rect -993 -50 -964 -44
rect -764 44 -735 50
rect -764 -44 -758 44
rect -741 -44 -735 44
rect -764 -50 -735 -44
rect -705 44 -676 50
rect -705 -44 -699 44
rect -682 -44 -676 44
rect -705 -50 -676 -44
rect -476 44 -447 50
rect -476 -44 -470 44
rect -453 -44 -447 44
rect -476 -50 -447 -44
rect -417 44 -388 50
rect -417 -44 -411 44
rect -394 -44 -388 44
rect -417 -50 -388 -44
rect -188 44 -159 50
rect -188 -44 -182 44
rect -165 -44 -159 44
rect -188 -50 -159 -44
rect -129 44 -100 50
rect -129 -44 -123 44
rect -106 -44 -100 44
rect -129 -50 -100 -44
rect 100 44 129 50
rect 100 -44 106 44
rect 123 -44 129 44
rect 100 -50 129 -44
rect 159 44 188 50
rect 159 -44 165 44
rect 182 -44 188 44
rect 159 -50 188 -44
rect 388 44 417 50
rect 388 -44 394 44
rect 411 -44 417 44
rect 388 -50 417 -44
rect 447 44 476 50
rect 447 -44 453 44
rect 470 -44 476 44
rect 447 -50 476 -44
rect 676 44 705 50
rect 676 -44 682 44
rect 699 -44 705 44
rect 676 -50 705 -44
rect 735 44 764 50
rect 735 -44 741 44
rect 758 -44 764 44
rect 735 -50 764 -44
rect 964 44 993 50
rect 964 -44 970 44
rect 987 -44 993 44
rect 964 -50 993 -44
rect 1023 44 1052 50
rect 1023 -44 1029 44
rect 1046 -44 1052 44
rect 1023 -50 1052 -44
rect 1252 44 1281 50
rect 1252 -44 1258 44
rect 1275 -44 1281 44
rect 1252 -50 1281 -44
rect 1311 44 1340 50
rect 1311 -44 1317 44
rect 1334 -44 1340 44
rect 1311 -50 1340 -44
rect 1540 44 1569 50
rect 1540 -44 1546 44
rect 1563 -44 1569 44
rect 1540 -50 1569 -44
rect 1599 44 1628 50
rect 1599 -44 1605 44
rect 1622 -44 1628 44
rect 1599 -50 1628 -44
rect 1828 44 1857 50
rect 1828 -44 1834 44
rect 1851 -44 1857 44
rect 1828 -50 1857 -44
rect 1887 44 1916 50
rect 1887 -44 1893 44
rect 1910 -44 1916 44
rect 1887 -50 1916 -44
rect 2116 44 2145 50
rect 2116 -44 2122 44
rect 2139 -44 2145 44
rect 2116 -50 2145 -44
rect 2175 44 2204 50
rect 2175 -44 2181 44
rect 2198 -44 2204 44
rect 2175 -50 2204 -44
rect 2404 44 2433 50
rect 2404 -44 2410 44
rect 2427 -44 2433 44
rect 2404 -50 2433 -44
rect 2463 44 2492 50
rect 2463 -44 2469 44
rect 2486 -44 2492 44
rect 2463 -50 2492 -44
rect 2692 44 2721 50
rect 2692 -44 2698 44
rect 2715 -44 2721 44
rect 2692 -50 2721 -44
rect 2751 44 2780 50
rect 2751 -44 2757 44
rect 2774 -44 2780 44
rect 2751 -50 2780 -44
rect 2980 44 3009 50
rect 2980 -44 2986 44
rect 3003 -44 3009 44
rect 2980 -50 3009 -44
rect 3039 44 3068 50
rect 3039 -44 3045 44
rect 3062 -44 3068 44
rect 3039 -50 3068 -44
rect 3268 44 3297 50
rect 3268 -44 3274 44
rect 3291 -44 3297 44
rect 3268 -50 3297 -44
rect 3327 44 3356 50
rect 3327 -44 3333 44
rect 3350 -44 3356 44
rect 3327 -50 3356 -44
rect 3556 44 3585 50
rect 3556 -44 3562 44
rect 3579 -44 3585 44
rect 3556 -50 3585 -44
<< mvndiffc >>
rect -3579 -44 -3562 44
rect -3350 -44 -3333 44
rect -3291 -44 -3274 44
rect -3062 -44 -3045 44
rect -3003 -44 -2986 44
rect -2774 -44 -2757 44
rect -2715 -44 -2698 44
rect -2486 -44 -2469 44
rect -2427 -44 -2410 44
rect -2198 -44 -2181 44
rect -2139 -44 -2122 44
rect -1910 -44 -1893 44
rect -1851 -44 -1834 44
rect -1622 -44 -1605 44
rect -1563 -44 -1546 44
rect -1334 -44 -1317 44
rect -1275 -44 -1258 44
rect -1046 -44 -1029 44
rect -987 -44 -970 44
rect -758 -44 -741 44
rect -699 -44 -682 44
rect -470 -44 -453 44
rect -411 -44 -394 44
rect -182 -44 -165 44
rect -123 -44 -106 44
rect 106 -44 123 44
rect 165 -44 182 44
rect 394 -44 411 44
rect 453 -44 470 44
rect 682 -44 699 44
rect 741 -44 758 44
rect 970 -44 987 44
rect 1029 -44 1046 44
rect 1258 -44 1275 44
rect 1317 -44 1334 44
rect 1546 -44 1563 44
rect 1605 -44 1622 44
rect 1834 -44 1851 44
rect 1893 -44 1910 44
rect 2122 -44 2139 44
rect 2181 -44 2198 44
rect 2410 -44 2427 44
rect 2469 -44 2486 44
rect 2698 -44 2715 44
rect 2757 -44 2774 44
rect 2986 -44 3003 44
rect 3045 -44 3062 44
rect 3274 -44 3291 44
rect 3333 -44 3350 44
rect 3562 -44 3579 44
<< mvpsubdiff >>
rect -3652 155 3652 161
rect -3652 138 -3598 155
rect 3598 138 3652 155
rect -3652 132 3652 138
rect -3652 107 -3623 132
rect -3652 -107 -3646 107
rect -3629 -107 -3623 107
rect 3623 107 3652 132
rect -3652 -132 -3623 -107
rect 3623 -107 3629 107
rect 3646 -107 3652 107
rect 3623 -132 3652 -107
rect -3652 -138 3652 -132
rect -3652 -155 -3598 -138
rect 3598 -155 3652 -138
rect -3652 -161 3652 -155
<< mvpsubdiffcont >>
rect -3598 138 3598 155
rect -3646 -107 -3629 107
rect 3629 -107 3646 107
rect -3598 -155 3598 -138
<< poly >>
rect -3556 86 -3356 94
rect -3556 69 -3548 86
rect -3364 69 -3356 86
rect -3556 50 -3356 69
rect -3268 86 -3068 94
rect -3268 69 -3260 86
rect -3076 69 -3068 86
rect -3268 50 -3068 69
rect -2980 86 -2780 94
rect -2980 69 -2972 86
rect -2788 69 -2780 86
rect -2980 50 -2780 69
rect -2692 86 -2492 94
rect -2692 69 -2684 86
rect -2500 69 -2492 86
rect -2692 50 -2492 69
rect -2404 86 -2204 94
rect -2404 69 -2396 86
rect -2212 69 -2204 86
rect -2404 50 -2204 69
rect -2116 86 -1916 94
rect -2116 69 -2108 86
rect -1924 69 -1916 86
rect -2116 50 -1916 69
rect -1828 86 -1628 94
rect -1828 69 -1820 86
rect -1636 69 -1628 86
rect -1828 50 -1628 69
rect -1540 86 -1340 94
rect -1540 69 -1532 86
rect -1348 69 -1340 86
rect -1540 50 -1340 69
rect -1252 86 -1052 94
rect -1252 69 -1244 86
rect -1060 69 -1052 86
rect -1252 50 -1052 69
rect -964 86 -764 94
rect -964 69 -956 86
rect -772 69 -764 86
rect -964 50 -764 69
rect -676 86 -476 94
rect -676 69 -668 86
rect -484 69 -476 86
rect -676 50 -476 69
rect -388 86 -188 94
rect -388 69 -380 86
rect -196 69 -188 86
rect -388 50 -188 69
rect -100 86 100 94
rect -100 69 -92 86
rect 92 69 100 86
rect -100 50 100 69
rect 188 86 388 94
rect 188 69 196 86
rect 380 69 388 86
rect 188 50 388 69
rect 476 86 676 94
rect 476 69 484 86
rect 668 69 676 86
rect 476 50 676 69
rect 764 86 964 94
rect 764 69 772 86
rect 956 69 964 86
rect 764 50 964 69
rect 1052 86 1252 94
rect 1052 69 1060 86
rect 1244 69 1252 86
rect 1052 50 1252 69
rect 1340 86 1540 94
rect 1340 69 1348 86
rect 1532 69 1540 86
rect 1340 50 1540 69
rect 1628 86 1828 94
rect 1628 69 1636 86
rect 1820 69 1828 86
rect 1628 50 1828 69
rect 1916 86 2116 94
rect 1916 69 1924 86
rect 2108 69 2116 86
rect 1916 50 2116 69
rect 2204 86 2404 94
rect 2204 69 2212 86
rect 2396 69 2404 86
rect 2204 50 2404 69
rect 2492 86 2692 94
rect 2492 69 2500 86
rect 2684 69 2692 86
rect 2492 50 2692 69
rect 2780 86 2980 94
rect 2780 69 2788 86
rect 2972 69 2980 86
rect 2780 50 2980 69
rect 3068 86 3268 94
rect 3068 69 3076 86
rect 3260 69 3268 86
rect 3068 50 3268 69
rect 3356 86 3556 94
rect 3356 69 3364 86
rect 3548 69 3556 86
rect 3356 50 3556 69
rect -3556 -69 -3356 -50
rect -3556 -86 -3548 -69
rect -3364 -86 -3356 -69
rect -3556 -94 -3356 -86
rect -3268 -69 -3068 -50
rect -3268 -86 -3260 -69
rect -3076 -86 -3068 -69
rect -3268 -94 -3068 -86
rect -2980 -69 -2780 -50
rect -2980 -86 -2972 -69
rect -2788 -86 -2780 -69
rect -2980 -94 -2780 -86
rect -2692 -69 -2492 -50
rect -2692 -86 -2684 -69
rect -2500 -86 -2492 -69
rect -2692 -94 -2492 -86
rect -2404 -69 -2204 -50
rect -2404 -86 -2396 -69
rect -2212 -86 -2204 -69
rect -2404 -94 -2204 -86
rect -2116 -69 -1916 -50
rect -2116 -86 -2108 -69
rect -1924 -86 -1916 -69
rect -2116 -94 -1916 -86
rect -1828 -69 -1628 -50
rect -1828 -86 -1820 -69
rect -1636 -86 -1628 -69
rect -1828 -94 -1628 -86
rect -1540 -69 -1340 -50
rect -1540 -86 -1532 -69
rect -1348 -86 -1340 -69
rect -1540 -94 -1340 -86
rect -1252 -69 -1052 -50
rect -1252 -86 -1244 -69
rect -1060 -86 -1052 -69
rect -1252 -94 -1052 -86
rect -964 -69 -764 -50
rect -964 -86 -956 -69
rect -772 -86 -764 -69
rect -964 -94 -764 -86
rect -676 -69 -476 -50
rect -676 -86 -668 -69
rect -484 -86 -476 -69
rect -676 -94 -476 -86
rect -388 -69 -188 -50
rect -388 -86 -380 -69
rect -196 -86 -188 -69
rect -388 -94 -188 -86
rect -100 -69 100 -50
rect -100 -86 -92 -69
rect 92 -86 100 -69
rect -100 -94 100 -86
rect 188 -69 388 -50
rect 188 -86 196 -69
rect 380 -86 388 -69
rect 188 -94 388 -86
rect 476 -69 676 -50
rect 476 -86 484 -69
rect 668 -86 676 -69
rect 476 -94 676 -86
rect 764 -69 964 -50
rect 764 -86 772 -69
rect 956 -86 964 -69
rect 764 -94 964 -86
rect 1052 -69 1252 -50
rect 1052 -86 1060 -69
rect 1244 -86 1252 -69
rect 1052 -94 1252 -86
rect 1340 -69 1540 -50
rect 1340 -86 1348 -69
rect 1532 -86 1540 -69
rect 1340 -94 1540 -86
rect 1628 -69 1828 -50
rect 1628 -86 1636 -69
rect 1820 -86 1828 -69
rect 1628 -94 1828 -86
rect 1916 -69 2116 -50
rect 1916 -86 1924 -69
rect 2108 -86 2116 -69
rect 1916 -94 2116 -86
rect 2204 -69 2404 -50
rect 2204 -86 2212 -69
rect 2396 -86 2404 -69
rect 2204 -94 2404 -86
rect 2492 -69 2692 -50
rect 2492 -86 2500 -69
rect 2684 -86 2692 -69
rect 2492 -94 2692 -86
rect 2780 -69 2980 -50
rect 2780 -86 2788 -69
rect 2972 -86 2980 -69
rect 2780 -94 2980 -86
rect 3068 -69 3268 -50
rect 3068 -86 3076 -69
rect 3260 -86 3268 -69
rect 3068 -94 3268 -86
rect 3356 -69 3556 -50
rect 3356 -86 3364 -69
rect 3548 -86 3556 -69
rect 3356 -94 3556 -86
<< polycont >>
rect -3548 69 -3364 86
rect -3260 69 -3076 86
rect -2972 69 -2788 86
rect -2684 69 -2500 86
rect -2396 69 -2212 86
rect -2108 69 -1924 86
rect -1820 69 -1636 86
rect -1532 69 -1348 86
rect -1244 69 -1060 86
rect -956 69 -772 86
rect -668 69 -484 86
rect -380 69 -196 86
rect -92 69 92 86
rect 196 69 380 86
rect 484 69 668 86
rect 772 69 956 86
rect 1060 69 1244 86
rect 1348 69 1532 86
rect 1636 69 1820 86
rect 1924 69 2108 86
rect 2212 69 2396 86
rect 2500 69 2684 86
rect 2788 69 2972 86
rect 3076 69 3260 86
rect 3364 69 3548 86
rect -3548 -86 -3364 -69
rect -3260 -86 -3076 -69
rect -2972 -86 -2788 -69
rect -2684 -86 -2500 -69
rect -2396 -86 -2212 -69
rect -2108 -86 -1924 -69
rect -1820 -86 -1636 -69
rect -1532 -86 -1348 -69
rect -1244 -86 -1060 -69
rect -956 -86 -772 -69
rect -668 -86 -484 -69
rect -380 -86 -196 -69
rect -92 -86 92 -69
rect 196 -86 380 -69
rect 484 -86 668 -69
rect 772 -86 956 -69
rect 1060 -86 1244 -69
rect 1348 -86 1532 -69
rect 1636 -86 1820 -69
rect 1924 -86 2108 -69
rect 2212 -86 2396 -69
rect 2500 -86 2684 -69
rect 2788 -86 2972 -69
rect 3076 -86 3260 -69
rect 3364 -86 3548 -69
<< locali >>
rect -3646 138 -3598 155
rect 3598 138 3646 155
rect -3646 107 -3629 138
rect 3629 107 3646 138
rect -3556 69 -3548 86
rect -3364 69 -3356 86
rect -3268 69 -3260 86
rect -3076 69 -3068 86
rect -2980 69 -2972 86
rect -2788 69 -2780 86
rect -2692 69 -2684 86
rect -2500 69 -2492 86
rect -2404 69 -2396 86
rect -2212 69 -2204 86
rect -2116 69 -2108 86
rect -1924 69 -1916 86
rect -1828 69 -1820 86
rect -1636 69 -1628 86
rect -1540 69 -1532 86
rect -1348 69 -1340 86
rect -1252 69 -1244 86
rect -1060 69 -1052 86
rect -964 69 -956 86
rect -772 69 -764 86
rect -676 69 -668 86
rect -484 69 -476 86
rect -388 69 -380 86
rect -196 69 -188 86
rect -100 69 -92 86
rect 92 69 100 86
rect 188 69 196 86
rect 380 69 388 86
rect 476 69 484 86
rect 668 69 676 86
rect 764 69 772 86
rect 956 69 964 86
rect 1052 69 1060 86
rect 1244 69 1252 86
rect 1340 69 1348 86
rect 1532 69 1540 86
rect 1628 69 1636 86
rect 1820 69 1828 86
rect 1916 69 1924 86
rect 2108 69 2116 86
rect 2204 69 2212 86
rect 2396 69 2404 86
rect 2492 69 2500 86
rect 2684 69 2692 86
rect 2780 69 2788 86
rect 2972 69 2980 86
rect 3068 69 3076 86
rect 3260 69 3268 86
rect 3356 69 3364 86
rect 3548 69 3556 86
rect -3579 44 -3562 52
rect -3579 -52 -3562 -44
rect -3350 44 -3333 52
rect -3350 -52 -3333 -44
rect -3291 44 -3274 52
rect -3291 -52 -3274 -44
rect -3062 44 -3045 52
rect -3062 -52 -3045 -44
rect -3003 44 -2986 52
rect -3003 -52 -2986 -44
rect -2774 44 -2757 52
rect -2774 -52 -2757 -44
rect -2715 44 -2698 52
rect -2715 -52 -2698 -44
rect -2486 44 -2469 52
rect -2486 -52 -2469 -44
rect -2427 44 -2410 52
rect -2427 -52 -2410 -44
rect -2198 44 -2181 52
rect -2198 -52 -2181 -44
rect -2139 44 -2122 52
rect -2139 -52 -2122 -44
rect -1910 44 -1893 52
rect -1910 -52 -1893 -44
rect -1851 44 -1834 52
rect -1851 -52 -1834 -44
rect -1622 44 -1605 52
rect -1622 -52 -1605 -44
rect -1563 44 -1546 52
rect -1563 -52 -1546 -44
rect -1334 44 -1317 52
rect -1334 -52 -1317 -44
rect -1275 44 -1258 52
rect -1275 -52 -1258 -44
rect -1046 44 -1029 52
rect -1046 -52 -1029 -44
rect -987 44 -970 52
rect -987 -52 -970 -44
rect -758 44 -741 52
rect -758 -52 -741 -44
rect -699 44 -682 52
rect -699 -52 -682 -44
rect -470 44 -453 52
rect -470 -52 -453 -44
rect -411 44 -394 52
rect -411 -52 -394 -44
rect -182 44 -165 52
rect -182 -52 -165 -44
rect -123 44 -106 52
rect -123 -52 -106 -44
rect 106 44 123 52
rect 106 -52 123 -44
rect 165 44 182 52
rect 165 -52 182 -44
rect 394 44 411 52
rect 394 -52 411 -44
rect 453 44 470 52
rect 453 -52 470 -44
rect 682 44 699 52
rect 682 -52 699 -44
rect 741 44 758 52
rect 741 -52 758 -44
rect 970 44 987 52
rect 970 -52 987 -44
rect 1029 44 1046 52
rect 1029 -52 1046 -44
rect 1258 44 1275 52
rect 1258 -52 1275 -44
rect 1317 44 1334 52
rect 1317 -52 1334 -44
rect 1546 44 1563 52
rect 1546 -52 1563 -44
rect 1605 44 1622 52
rect 1605 -52 1622 -44
rect 1834 44 1851 52
rect 1834 -52 1851 -44
rect 1893 44 1910 52
rect 1893 -52 1910 -44
rect 2122 44 2139 52
rect 2122 -52 2139 -44
rect 2181 44 2198 52
rect 2181 -52 2198 -44
rect 2410 44 2427 52
rect 2410 -52 2427 -44
rect 2469 44 2486 52
rect 2469 -52 2486 -44
rect 2698 44 2715 52
rect 2698 -52 2715 -44
rect 2757 44 2774 52
rect 2757 -52 2774 -44
rect 2986 44 3003 52
rect 2986 -52 3003 -44
rect 3045 44 3062 52
rect 3045 -52 3062 -44
rect 3274 44 3291 52
rect 3274 -52 3291 -44
rect 3333 44 3350 52
rect 3333 -52 3350 -44
rect 3562 44 3579 52
rect 3562 -52 3579 -44
rect -3556 -86 -3548 -69
rect -3364 -86 -3356 -69
rect -3268 -86 -3260 -69
rect -3076 -86 -3068 -69
rect -2980 -86 -2972 -69
rect -2788 -86 -2780 -69
rect -2692 -86 -2684 -69
rect -2500 -86 -2492 -69
rect -2404 -86 -2396 -69
rect -2212 -86 -2204 -69
rect -2116 -86 -2108 -69
rect -1924 -86 -1916 -69
rect -1828 -86 -1820 -69
rect -1636 -86 -1628 -69
rect -1540 -86 -1532 -69
rect -1348 -86 -1340 -69
rect -1252 -86 -1244 -69
rect -1060 -86 -1052 -69
rect -964 -86 -956 -69
rect -772 -86 -764 -69
rect -676 -86 -668 -69
rect -484 -86 -476 -69
rect -388 -86 -380 -69
rect -196 -86 -188 -69
rect -100 -86 -92 -69
rect 92 -86 100 -69
rect 188 -86 196 -69
rect 380 -86 388 -69
rect 476 -86 484 -69
rect 668 -86 676 -69
rect 764 -86 772 -69
rect 956 -86 964 -69
rect 1052 -86 1060 -69
rect 1244 -86 1252 -69
rect 1340 -86 1348 -69
rect 1532 -86 1540 -69
rect 1628 -86 1636 -69
rect 1820 -86 1828 -69
rect 1916 -86 1924 -69
rect 2108 -86 2116 -69
rect 2204 -86 2212 -69
rect 2396 -86 2404 -69
rect 2492 -86 2500 -69
rect 2684 -86 2692 -69
rect 2780 -86 2788 -69
rect 2972 -86 2980 -69
rect 3068 -86 3076 -69
rect 3260 -86 3268 -69
rect 3356 -86 3364 -69
rect 3548 -86 3556 -69
rect -3646 -138 -3629 -107
rect 3629 -138 3646 -107
rect -3646 -155 -3598 -138
rect 3598 -155 3646 -138
<< viali >>
rect -3548 69 -3364 86
rect -3260 69 -3076 86
rect -2972 69 -2788 86
rect -2684 69 -2500 86
rect -2396 69 -2212 86
rect -2108 69 -1924 86
rect -1820 69 -1636 86
rect -1532 69 -1348 86
rect -1244 69 -1060 86
rect -956 69 -772 86
rect -668 69 -484 86
rect -380 69 -196 86
rect -92 69 92 86
rect 196 69 380 86
rect 484 69 668 86
rect 772 69 956 86
rect 1060 69 1244 86
rect 1348 69 1532 86
rect 1636 69 1820 86
rect 1924 69 2108 86
rect 2212 69 2396 86
rect 2500 69 2684 86
rect 2788 69 2972 86
rect 3076 69 3260 86
rect 3364 69 3548 86
rect -3579 -44 -3562 44
rect -3350 -44 -3333 44
rect -3291 -44 -3274 44
rect -3062 -44 -3045 44
rect -3003 -44 -2986 44
rect -2774 -44 -2757 44
rect -2715 -44 -2698 44
rect -2486 -44 -2469 44
rect -2427 -44 -2410 44
rect -2198 -44 -2181 44
rect -2139 -44 -2122 44
rect -1910 -44 -1893 44
rect -1851 -44 -1834 44
rect -1622 -44 -1605 44
rect -1563 -44 -1546 44
rect -1334 -44 -1317 44
rect -1275 -44 -1258 44
rect -1046 -44 -1029 44
rect -987 -44 -970 44
rect -758 -44 -741 44
rect -699 -44 -682 44
rect -470 -44 -453 44
rect -411 -44 -394 44
rect -182 -44 -165 44
rect -123 -44 -106 44
rect 106 -44 123 44
rect 165 -44 182 44
rect 394 -44 411 44
rect 453 -44 470 44
rect 682 -44 699 44
rect 741 -44 758 44
rect 970 -44 987 44
rect 1029 -44 1046 44
rect 1258 -44 1275 44
rect 1317 -44 1334 44
rect 1546 -44 1563 44
rect 1605 -44 1622 44
rect 1834 -44 1851 44
rect 1893 -44 1910 44
rect 2122 -44 2139 44
rect 2181 -44 2198 44
rect 2410 -44 2427 44
rect 2469 -44 2486 44
rect 2698 -44 2715 44
rect 2757 -44 2774 44
rect 2986 -44 3003 44
rect 3045 -44 3062 44
rect 3274 -44 3291 44
rect 3333 -44 3350 44
rect 3562 -44 3579 44
rect -3548 -86 -3364 -69
rect -3260 -86 -3076 -69
rect -2972 -86 -2788 -69
rect -2684 -86 -2500 -69
rect -2396 -86 -2212 -69
rect -2108 -86 -1924 -69
rect -1820 -86 -1636 -69
rect -1532 -86 -1348 -69
rect -1244 -86 -1060 -69
rect -956 -86 -772 -69
rect -668 -86 -484 -69
rect -380 -86 -196 -69
rect -92 -86 92 -69
rect 196 -86 380 -69
rect 484 -86 668 -69
rect 772 -86 956 -69
rect 1060 -86 1244 -69
rect 1348 -86 1532 -69
rect 1636 -86 1820 -69
rect 1924 -86 2108 -69
rect 2212 -86 2396 -69
rect 2500 -86 2684 -69
rect 2788 -86 2972 -69
rect 3076 -86 3260 -69
rect 3364 -86 3548 -69
<< metal1 >>
rect -3554 86 -3358 89
rect -3554 69 -3548 86
rect -3364 69 -3358 86
rect -3554 66 -3358 69
rect -3266 86 -3070 89
rect -3266 69 -3260 86
rect -3076 69 -3070 86
rect -3266 66 -3070 69
rect -2978 86 -2782 89
rect -2978 69 -2972 86
rect -2788 69 -2782 86
rect -2978 66 -2782 69
rect -2690 86 -2494 89
rect -2690 69 -2684 86
rect -2500 69 -2494 86
rect -2690 66 -2494 69
rect -2402 86 -2206 89
rect -2402 69 -2396 86
rect -2212 69 -2206 86
rect -2402 66 -2206 69
rect -2114 86 -1918 89
rect -2114 69 -2108 86
rect -1924 69 -1918 86
rect -2114 66 -1918 69
rect -1826 86 -1630 89
rect -1826 69 -1820 86
rect -1636 69 -1630 86
rect -1826 66 -1630 69
rect -1538 86 -1342 89
rect -1538 69 -1532 86
rect -1348 69 -1342 86
rect -1538 66 -1342 69
rect -1250 86 -1054 89
rect -1250 69 -1244 86
rect -1060 69 -1054 86
rect -1250 66 -1054 69
rect -962 86 -766 89
rect -962 69 -956 86
rect -772 69 -766 86
rect -962 66 -766 69
rect -674 86 -478 89
rect -674 69 -668 86
rect -484 69 -478 86
rect -674 66 -478 69
rect -386 86 -190 89
rect -386 69 -380 86
rect -196 69 -190 86
rect -386 66 -190 69
rect -98 86 98 89
rect -98 69 -92 86
rect 92 69 98 86
rect -98 66 98 69
rect 190 86 386 89
rect 190 69 196 86
rect 380 69 386 86
rect 190 66 386 69
rect 478 86 674 89
rect 478 69 484 86
rect 668 69 674 86
rect 478 66 674 69
rect 766 86 962 89
rect 766 69 772 86
rect 956 69 962 86
rect 766 66 962 69
rect 1054 86 1250 89
rect 1054 69 1060 86
rect 1244 69 1250 86
rect 1054 66 1250 69
rect 1342 86 1538 89
rect 1342 69 1348 86
rect 1532 69 1538 86
rect 1342 66 1538 69
rect 1630 86 1826 89
rect 1630 69 1636 86
rect 1820 69 1826 86
rect 1630 66 1826 69
rect 1918 86 2114 89
rect 1918 69 1924 86
rect 2108 69 2114 86
rect 1918 66 2114 69
rect 2206 86 2402 89
rect 2206 69 2212 86
rect 2396 69 2402 86
rect 2206 66 2402 69
rect 2494 86 2690 89
rect 2494 69 2500 86
rect 2684 69 2690 86
rect 2494 66 2690 69
rect 2782 86 2978 89
rect 2782 69 2788 86
rect 2972 69 2978 86
rect 2782 66 2978 69
rect 3070 86 3266 89
rect 3070 69 3076 86
rect 3260 69 3266 86
rect 3070 66 3266 69
rect 3358 86 3554 89
rect 3358 69 3364 86
rect 3548 69 3554 86
rect 3358 66 3554 69
rect -3582 44 -3559 50
rect -3582 -44 -3579 44
rect -3562 -44 -3559 44
rect -3582 -50 -3559 -44
rect -3353 44 -3330 50
rect -3353 -44 -3350 44
rect -3333 -44 -3330 44
rect -3353 -50 -3330 -44
rect -3294 44 -3271 50
rect -3294 -44 -3291 44
rect -3274 -44 -3271 44
rect -3294 -50 -3271 -44
rect -3065 44 -3042 50
rect -3065 -44 -3062 44
rect -3045 -44 -3042 44
rect -3065 -50 -3042 -44
rect -3006 44 -2983 50
rect -3006 -44 -3003 44
rect -2986 -44 -2983 44
rect -3006 -50 -2983 -44
rect -2777 44 -2754 50
rect -2777 -44 -2774 44
rect -2757 -44 -2754 44
rect -2777 -50 -2754 -44
rect -2718 44 -2695 50
rect -2718 -44 -2715 44
rect -2698 -44 -2695 44
rect -2718 -50 -2695 -44
rect -2489 44 -2466 50
rect -2489 -44 -2486 44
rect -2469 -44 -2466 44
rect -2489 -50 -2466 -44
rect -2430 44 -2407 50
rect -2430 -44 -2427 44
rect -2410 -44 -2407 44
rect -2430 -50 -2407 -44
rect -2201 44 -2178 50
rect -2201 -44 -2198 44
rect -2181 -44 -2178 44
rect -2201 -50 -2178 -44
rect -2142 44 -2119 50
rect -2142 -44 -2139 44
rect -2122 -44 -2119 44
rect -2142 -50 -2119 -44
rect -1913 44 -1890 50
rect -1913 -44 -1910 44
rect -1893 -44 -1890 44
rect -1913 -50 -1890 -44
rect -1854 44 -1831 50
rect -1854 -44 -1851 44
rect -1834 -44 -1831 44
rect -1854 -50 -1831 -44
rect -1625 44 -1602 50
rect -1625 -44 -1622 44
rect -1605 -44 -1602 44
rect -1625 -50 -1602 -44
rect -1566 44 -1543 50
rect -1566 -44 -1563 44
rect -1546 -44 -1543 44
rect -1566 -50 -1543 -44
rect -1337 44 -1314 50
rect -1337 -44 -1334 44
rect -1317 -44 -1314 44
rect -1337 -50 -1314 -44
rect -1278 44 -1255 50
rect -1278 -44 -1275 44
rect -1258 -44 -1255 44
rect -1278 -50 -1255 -44
rect -1049 44 -1026 50
rect -1049 -44 -1046 44
rect -1029 -44 -1026 44
rect -1049 -50 -1026 -44
rect -990 44 -967 50
rect -990 -44 -987 44
rect -970 -44 -967 44
rect -990 -50 -967 -44
rect -761 44 -738 50
rect -761 -44 -758 44
rect -741 -44 -738 44
rect -761 -50 -738 -44
rect -702 44 -679 50
rect -702 -44 -699 44
rect -682 -44 -679 44
rect -702 -50 -679 -44
rect -473 44 -450 50
rect -473 -44 -470 44
rect -453 -44 -450 44
rect -473 -50 -450 -44
rect -414 44 -391 50
rect -414 -44 -411 44
rect -394 -44 -391 44
rect -414 -50 -391 -44
rect -185 44 -162 50
rect -185 -44 -182 44
rect -165 -44 -162 44
rect -185 -50 -162 -44
rect -126 44 -103 50
rect -126 -44 -123 44
rect -106 -44 -103 44
rect -126 -50 -103 -44
rect 103 44 126 50
rect 103 -44 106 44
rect 123 -44 126 44
rect 103 -50 126 -44
rect 162 44 185 50
rect 162 -44 165 44
rect 182 -44 185 44
rect 162 -50 185 -44
rect 391 44 414 50
rect 391 -44 394 44
rect 411 -44 414 44
rect 391 -50 414 -44
rect 450 44 473 50
rect 450 -44 453 44
rect 470 -44 473 44
rect 450 -50 473 -44
rect 679 44 702 50
rect 679 -44 682 44
rect 699 -44 702 44
rect 679 -50 702 -44
rect 738 44 761 50
rect 738 -44 741 44
rect 758 -44 761 44
rect 738 -50 761 -44
rect 967 44 990 50
rect 967 -44 970 44
rect 987 -44 990 44
rect 967 -50 990 -44
rect 1026 44 1049 50
rect 1026 -44 1029 44
rect 1046 -44 1049 44
rect 1026 -50 1049 -44
rect 1255 44 1278 50
rect 1255 -44 1258 44
rect 1275 -44 1278 44
rect 1255 -50 1278 -44
rect 1314 44 1337 50
rect 1314 -44 1317 44
rect 1334 -44 1337 44
rect 1314 -50 1337 -44
rect 1543 44 1566 50
rect 1543 -44 1546 44
rect 1563 -44 1566 44
rect 1543 -50 1566 -44
rect 1602 44 1625 50
rect 1602 -44 1605 44
rect 1622 -44 1625 44
rect 1602 -50 1625 -44
rect 1831 44 1854 50
rect 1831 -44 1834 44
rect 1851 -44 1854 44
rect 1831 -50 1854 -44
rect 1890 44 1913 50
rect 1890 -44 1893 44
rect 1910 -44 1913 44
rect 1890 -50 1913 -44
rect 2119 44 2142 50
rect 2119 -44 2122 44
rect 2139 -44 2142 44
rect 2119 -50 2142 -44
rect 2178 44 2201 50
rect 2178 -44 2181 44
rect 2198 -44 2201 44
rect 2178 -50 2201 -44
rect 2407 44 2430 50
rect 2407 -44 2410 44
rect 2427 -44 2430 44
rect 2407 -50 2430 -44
rect 2466 44 2489 50
rect 2466 -44 2469 44
rect 2486 -44 2489 44
rect 2466 -50 2489 -44
rect 2695 44 2718 50
rect 2695 -44 2698 44
rect 2715 -44 2718 44
rect 2695 -50 2718 -44
rect 2754 44 2777 50
rect 2754 -44 2757 44
rect 2774 -44 2777 44
rect 2754 -50 2777 -44
rect 2983 44 3006 50
rect 2983 -44 2986 44
rect 3003 -44 3006 44
rect 2983 -50 3006 -44
rect 3042 44 3065 50
rect 3042 -44 3045 44
rect 3062 -44 3065 44
rect 3042 -50 3065 -44
rect 3271 44 3294 50
rect 3271 -44 3274 44
rect 3291 -44 3294 44
rect 3271 -50 3294 -44
rect 3330 44 3353 50
rect 3330 -44 3333 44
rect 3350 -44 3353 44
rect 3330 -50 3353 -44
rect 3559 44 3582 50
rect 3559 -44 3562 44
rect 3579 -44 3582 44
rect 3559 -50 3582 -44
rect -3554 -69 -3358 -66
rect -3554 -86 -3548 -69
rect -3364 -86 -3358 -69
rect -3554 -89 -3358 -86
rect -3266 -69 -3070 -66
rect -3266 -86 -3260 -69
rect -3076 -86 -3070 -69
rect -3266 -89 -3070 -86
rect -2978 -69 -2782 -66
rect -2978 -86 -2972 -69
rect -2788 -86 -2782 -69
rect -2978 -89 -2782 -86
rect -2690 -69 -2494 -66
rect -2690 -86 -2684 -69
rect -2500 -86 -2494 -69
rect -2690 -89 -2494 -86
rect -2402 -69 -2206 -66
rect -2402 -86 -2396 -69
rect -2212 -86 -2206 -69
rect -2402 -89 -2206 -86
rect -2114 -69 -1918 -66
rect -2114 -86 -2108 -69
rect -1924 -86 -1918 -69
rect -2114 -89 -1918 -86
rect -1826 -69 -1630 -66
rect -1826 -86 -1820 -69
rect -1636 -86 -1630 -69
rect -1826 -89 -1630 -86
rect -1538 -69 -1342 -66
rect -1538 -86 -1532 -69
rect -1348 -86 -1342 -69
rect -1538 -89 -1342 -86
rect -1250 -69 -1054 -66
rect -1250 -86 -1244 -69
rect -1060 -86 -1054 -69
rect -1250 -89 -1054 -86
rect -962 -69 -766 -66
rect -962 -86 -956 -69
rect -772 -86 -766 -69
rect -962 -89 -766 -86
rect -674 -69 -478 -66
rect -674 -86 -668 -69
rect -484 -86 -478 -69
rect -674 -89 -478 -86
rect -386 -69 -190 -66
rect -386 -86 -380 -69
rect -196 -86 -190 -69
rect -386 -89 -190 -86
rect -98 -69 98 -66
rect -98 -86 -92 -69
rect 92 -86 98 -69
rect -98 -89 98 -86
rect 190 -69 386 -66
rect 190 -86 196 -69
rect 380 -86 386 -69
rect 190 -89 386 -86
rect 478 -69 674 -66
rect 478 -86 484 -69
rect 668 -86 674 -69
rect 478 -89 674 -86
rect 766 -69 962 -66
rect 766 -86 772 -69
rect 956 -86 962 -69
rect 766 -89 962 -86
rect 1054 -69 1250 -66
rect 1054 -86 1060 -69
rect 1244 -86 1250 -69
rect 1054 -89 1250 -86
rect 1342 -69 1538 -66
rect 1342 -86 1348 -69
rect 1532 -86 1538 -69
rect 1342 -89 1538 -86
rect 1630 -69 1826 -66
rect 1630 -86 1636 -69
rect 1820 -86 1826 -69
rect 1630 -89 1826 -86
rect 1918 -69 2114 -66
rect 1918 -86 1924 -69
rect 2108 -86 2114 -69
rect 1918 -89 2114 -86
rect 2206 -69 2402 -66
rect 2206 -86 2212 -69
rect 2396 -86 2402 -69
rect 2206 -89 2402 -86
rect 2494 -69 2690 -66
rect 2494 -86 2500 -69
rect 2684 -86 2690 -69
rect 2494 -89 2690 -86
rect 2782 -69 2978 -66
rect 2782 -86 2788 -69
rect 2972 -86 2978 -69
rect 2782 -89 2978 -86
rect 3070 -69 3266 -66
rect 3070 -86 3076 -69
rect 3260 -86 3266 -69
rect 3070 -89 3266 -86
rect 3358 -69 3554 -66
rect 3358 -86 3364 -69
rect 3548 -86 3554 -69
rect 3358 -89 3554 -86
<< properties >>
string FIXED_BBOX -3637 -146 3637 146
string gencell sky130_fd_pr__nfet_05v0_nvt
string library sky130
string parameters w 1.0 l 2.0 m 1 nf 25 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.90 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
