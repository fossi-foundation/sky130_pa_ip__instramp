magic
tech sky130A
magscale 1 2
timestamp 1730992657
<< dnwell >>
rect 3906 -2698 7768 -412
<< locali >>
rect 2770 -236 3082 -224
rect 2770 -320 2782 -236
rect 3064 -320 3082 -236
rect 2770 -330 3082 -320
rect 2892 -390 2982 -384
rect 2892 -612 2906 -390
rect 2966 -612 2982 -390
rect 2892 -620 2982 -612
rect 4196 -388 4820 -370
rect 4196 -478 4206 -388
rect 4808 -478 4820 -388
rect 4196 -698 4820 -478
rect 5970 -388 6594 -368
rect 5970 -476 5982 -388
rect 6574 -476 6594 -388
rect 5970 -696 6594 -476
rect 5000 -1226 5650 -1074
rect 5000 -1326 5016 -1226
rect 5334 -1326 5650 -1226
rect 5000 -1340 5650 -1326
rect 6762 -1224 7412 -1076
rect 6762 -1330 6940 -1224
rect 7394 -1330 7412 -1224
rect 6762 -1342 7412 -1330
rect 4176 -1404 7362 -1402
rect 4176 -1408 7390 -1404
rect 4176 -1458 4316 -1408
rect 6704 -1414 7390 -1408
rect 6704 -1458 7334 -1414
rect 4176 -1462 7334 -1458
rect 4176 -1470 4206 -1462
rect 4180 -2562 4206 -1470
rect 4176 -2572 4206 -2562
rect 4276 -1470 7334 -1462
rect 4276 -2562 4292 -1470
rect 7322 -1992 7334 -1470
rect 7382 -1992 7390 -1414
rect 7322 -2562 7390 -1992
rect 4276 -2568 7390 -2562
rect 4276 -2572 4330 -2568
rect 4176 -2618 4330 -2572
rect 7374 -2618 7390 -2568
rect 4176 -2630 7390 -2618
<< viali >>
rect 2782 -320 3064 -236
rect 1958 -496 2116 -420
rect 2906 -612 2966 -390
rect 4206 -478 4808 -388
rect 5982 -476 6574 -388
rect 5016 -1326 5334 -1226
rect 6940 -1330 7394 -1224
rect 4316 -1458 6704 -1408
rect 1966 -2182 2102 -2118
rect 4206 -2572 4276 -1462
rect 7334 -1992 7382 -1414
rect 4330 -2618 7374 -2568
<< metal1 >>
rect 2770 -236 3082 -224
rect 1668 -1594 1736 -264
rect 1944 -420 2128 -406
rect 1944 -496 1958 -420
rect 2116 -496 2128 -420
rect 1944 -508 2128 -496
rect 1668 -2664 1736 -1934
rect 2012 -2092 2054 -508
rect 2376 -1124 2558 -264
rect 2770 -320 2782 -236
rect 3064 -320 3082 -236
rect 3206 -266 3306 -264
rect 2770 -330 3082 -320
rect 2892 -390 2982 -384
rect 2892 -612 2906 -390
rect 2966 -612 2982 -390
rect 2892 -620 2982 -612
rect 1958 -2118 2108 -2092
rect 1958 -2182 1966 -2118
rect 2102 -2182 2108 -2118
rect 1958 -2190 2108 -2182
rect 1958 -2260 1966 -2190
rect 2102 -2260 2108 -2190
rect 1958 -2270 2108 -2260
rect 2120 -2648 2320 -2448
rect 2376 -2464 2558 -1444
rect 3204 -1584 3278 -266
rect 3670 -368 3814 -356
rect 3670 -1578 3814 -490
rect 4198 -388 4818 -368
rect 4198 -478 4206 -388
rect 4808 -478 4818 -388
rect 4198 -492 4818 -478
rect 5968 -388 6588 -362
rect 5968 -476 5982 -388
rect 6574 -476 6588 -388
rect 5968 -486 6588 -476
rect 5324 -554 5420 -534
rect 5324 -814 5420 -628
rect 5692 -778 5892 -772
rect 5692 -864 5892 -838
rect 3908 -938 4122 -930
rect 7462 -938 7670 -928
rect 3908 -1004 4122 -998
rect 5002 -1226 5354 -1208
rect 5002 -1326 5016 -1226
rect 5334 -1326 5354 -1226
rect 5404 -1226 5492 -980
rect 7462 -1008 7670 -998
rect 6792 -1226 6888 -1024
rect 5404 -1314 6888 -1226
rect 5002 -1340 5354 -1326
rect 4162 -1408 6718 -1398
rect 4162 -1430 4316 -1408
rect 3204 -1728 3210 -1584
rect 3204 -2462 3278 -1728
rect 2376 -2664 2588 -2464
rect 3116 -2662 3316 -2462
rect 3164 -2664 3312 -2662
rect 3670 -2760 3814 -1732
rect 4138 -1458 4316 -1430
rect 6704 -1458 6718 -1408
rect 4138 -2564 4162 -1458
rect 4272 -1462 6718 -1458
rect 4276 -1466 6718 -1462
rect 6792 -1462 6888 -1314
rect 6926 -1224 7412 -1208
rect 6926 -1330 6940 -1224
rect 7394 -1330 7412 -1224
rect 6926 -1340 7412 -1330
rect 7322 -1414 7392 -1402
rect 7102 -1462 7190 -1460
rect 4276 -2562 4298 -1466
rect 4392 -1802 4828 -1566
rect 6792 -1636 7228 -1462
rect 4394 -2136 4830 -1900
rect 6792 -1970 7226 -1730
rect 7322 -1992 7334 -1414
rect 7382 -1992 7392 -1414
rect 7322 -2008 7392 -1992
rect 7472 -2064 7672 -1948
rect 6790 -2134 7672 -2064
rect 6790 -2230 7226 -2134
rect 7472 -2148 7672 -2134
rect 4390 -2466 4826 -2230
rect 6790 -2298 7228 -2230
rect 6792 -2300 7228 -2298
rect 7472 -2392 7672 -2378
rect 6792 -2472 7672 -2392
rect 4138 -2572 4206 -2564
rect 4276 -2568 7388 -2562
rect 4276 -2572 4330 -2568
rect 4138 -2598 4330 -2572
rect 4176 -2618 4330 -2598
rect 7374 -2618 7388 -2568
rect 7472 -2578 7672 -2472
rect 4176 -2630 7388 -2618
<< via1 >>
rect 1656 -1934 1762 -1594
rect 2782 -320 3064 -236
rect 2906 -612 2966 -390
rect 2370 -1444 2584 -1124
rect 1966 -2260 2102 -2190
rect 3670 -490 3814 -368
rect 4206 -478 4808 -388
rect 5982 -476 6574 -388
rect 5324 -628 5420 -554
rect 5692 -838 5892 -778
rect 6844 -804 7160 -722
rect 3908 -998 4122 -938
rect 5016 -1326 5334 -1226
rect 7462 -998 7670 -938
rect 3210 -1728 3306 -1584
rect 3670 -1732 3814 -1578
rect 4162 -1462 4272 -1458
rect 4162 -2564 4206 -1462
rect 4206 -2564 4272 -1462
rect 6940 -1330 7394 -1224
<< metal2 >>
rect 2770 -236 3082 -224
rect 2770 -320 2782 -236
rect 3064 -242 3082 -236
rect 3064 -302 3544 -242
rect 3064 -320 3082 -302
rect 2770 -330 3082 -320
rect 2892 -390 2982 -384
rect 2892 -612 2906 -390
rect 2966 -402 2982 -390
rect 2966 -462 3444 -402
rect 2966 -612 2982 -462
rect 2892 -620 2982 -612
rect 3384 -938 3444 -462
rect 3484 -778 3544 -302
rect 3661 -490 3670 -368
rect 3814 -388 6624 -368
rect 3814 -478 4206 -388
rect 4808 -476 5982 -388
rect 6574 -476 6624 -388
rect 4808 -478 6624 -476
rect 3814 -490 6624 -478
rect 7476 -554 7676 -428
rect 5317 -628 5324 -554
rect 5420 -628 7676 -554
rect 7476 -722 7676 -670
rect 3484 -838 5692 -778
rect 5892 -838 5926 -778
rect 6819 -804 6844 -722
rect 7160 -804 7676 -722
rect 7476 -870 7676 -804
rect 3384 -998 3908 -938
rect 4122 -998 7462 -938
rect 7670 -998 7678 -938
rect 2350 -1124 2600 -1110
rect 2350 -1210 2370 -1124
rect 2349 -1340 2370 -1210
rect 2350 -1444 2370 -1340
rect 2584 -1210 2600 -1124
rect 2584 -1224 7408 -1210
rect 2584 -1226 6940 -1224
rect 2584 -1326 5016 -1226
rect 5334 -1326 6940 -1226
rect 2584 -1330 6940 -1326
rect 7394 -1330 7408 -1224
rect 2584 -1340 7408 -1330
rect 2584 -1444 2600 -1340
rect 2350 -1466 2600 -1444
rect 4138 -1458 4298 -1430
rect 1642 -1578 1782 -1564
rect 4138 -1578 4162 -1458
rect 1642 -1584 3318 -1578
rect 1642 -1594 3210 -1584
rect 1642 -1934 1656 -1594
rect 1762 -1728 3210 -1594
rect 3306 -1728 3318 -1584
rect 1762 -1732 3318 -1728
rect 3654 -1732 3670 -1578
rect 3814 -1732 4162 -1578
rect 1762 -1934 1782 -1732
rect 1642 -1954 1782 -1934
rect 1610 -2190 1810 -2172
rect 1610 -2260 1966 -2190
rect 2102 -2260 2114 -2190
rect 1610 -2278 1810 -2260
rect 4138 -2564 4162 -1732
rect 4272 -1578 4298 -1458
rect 4272 -1732 4303 -1578
rect 4272 -2564 4298 -1732
rect 4138 -2598 4298 -2564
use sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP  sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP_0 paramcells
timestamp 1730992408
transform 0 1 5812 -1 0 -2016
box -616 -1582 616 1582
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1729530005
transform 0 1 1661 -1 0 -360
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1729530005
transform 0 1 1661 -1 0 -264
box -66 -43 162 897
use sky130_fd_sc_hvl__lsbuflv2hv_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1729530005
transform 0 1 1661 1 0 -2664
box -66 -43 2178 1671
use sky130_fd_sc_hvl__inv_1  x2 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1729530005
transform 0 -1 3289 1 0 -552
box -66 -43 354 897
use T_Gate_5V  x12
timestamp 1730992408
transform 0 -1 3862 -1 0 -160
box 422 -1926 1038 -134
use T_Gate_5V  x13
timestamp 1730992408
transform 0 -1 5632 -1 0 -160
box 422 -1926 1038 -134
<< labels >>
flabel metal2 7476 -870 7676 -670 0 FreeSans 256 180 0 0 CMOUT
port 3 nsew
flabel metal2 7476 -628 7676 -428 0 FreeSans 256 180 0 0 VIRTOUT
port 2 nsew
flabel metal1 7472 -2148 7672 -1948 0 FreeSans 256 180 0 0 R2ROUT
port 5 nsew
flabel metal1 7472 -2578 7672 -2378 0 FreeSans 256 180 0 0 R2RIN
port 4 nsew
flabel metal2 1610 -2278 1810 -2172 0 FreeSans 256 270 0 0 VD
port 0 nsew
flabel metal1 2120 -2648 2320 -2448 0 FreeSans 256 270 0 0 DVDD
port 1 nsew
flabel metal1 2388 -2664 2588 -2464 0 FreeSans 256 270 0 0 AVDD
port 7 nsew
flabel metal1 3116 -2662 3316 -2462 0 FreeSans 256 270 0 0 DVSS
port 6 nsew
flabel metal2 3372 -274 3372 -274 0 FreeSans 480 0 0 0 VDBAR
flabel metal2 3392 -434 3392 -434 0 FreeSans 480 0 0 0 VDbuf
flabel metal1 3670 -2632 3814 -2462 0 FreeSans 320 90 0 0 AVSS
port 8 nsew
<< end >>
