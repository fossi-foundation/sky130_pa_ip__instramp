magic
tech sky130A
magscale 1 2
timestamp 1730992408
<< pwell >>
rect -2442 -2562 2442 2562
<< psubdiff >>
rect -2406 2492 -2310 2526
rect 2310 2492 2406 2526
rect -2406 2430 -2372 2492
rect 2372 2430 2406 2492
rect -2406 -2492 -2372 -2430
rect 2372 -2492 2406 -2430
rect -2406 -2526 -2310 -2492
rect 2310 -2526 2406 -2492
<< psubdiffcont >>
rect -2310 2492 2310 2526
rect -2406 -2430 -2372 2430
rect 2372 -2430 2406 2430
rect -2310 -2526 2310 -2492
<< xpolycontact >>
rect -2276 1964 -2206 2396
rect -2276 -2396 -2206 -1964
rect -2110 1964 -2040 2396
rect -2110 -2396 -2040 -1964
rect -1944 1964 -1874 2396
rect -1944 -2396 -1874 -1964
rect -1778 1964 -1708 2396
rect -1778 -2396 -1708 -1964
rect -1612 1964 -1542 2396
rect -1612 -2396 -1542 -1964
rect -1446 1964 -1376 2396
rect -1446 -2396 -1376 -1964
rect -1280 1964 -1210 2396
rect -1280 -2396 -1210 -1964
rect -1114 1964 -1044 2396
rect -1114 -2396 -1044 -1964
rect -948 1964 -878 2396
rect -948 -2396 -878 -1964
rect -782 1964 -712 2396
rect -782 -2396 -712 -1964
rect -616 1964 -546 2396
rect -616 -2396 -546 -1964
rect -450 1964 -380 2396
rect -450 -2396 -380 -1964
rect -284 1964 -214 2396
rect -284 -2396 -214 -1964
rect -118 1964 -48 2396
rect -118 -2396 -48 -1964
rect 48 1964 118 2396
rect 48 -2396 118 -1964
rect 214 1964 284 2396
rect 214 -2396 284 -1964
rect 380 1964 450 2396
rect 380 -2396 450 -1964
rect 546 1964 616 2396
rect 546 -2396 616 -1964
rect 712 1964 782 2396
rect 712 -2396 782 -1964
rect 878 1964 948 2396
rect 878 -2396 948 -1964
rect 1044 1964 1114 2396
rect 1044 -2396 1114 -1964
rect 1210 1964 1280 2396
rect 1210 -2396 1280 -1964
rect 1376 1964 1446 2396
rect 1376 -2396 1446 -1964
rect 1542 1964 1612 2396
rect 1542 -2396 1612 -1964
rect 1708 1964 1778 2396
rect 1708 -2396 1778 -1964
rect 1874 1964 1944 2396
rect 1874 -2396 1944 -1964
rect 2040 1964 2110 2396
rect 2040 -2396 2110 -1964
rect 2206 1964 2276 2396
rect 2206 -2396 2276 -1964
<< xpolyres >>
rect -2276 -1964 -2206 1964
rect -2110 -1964 -2040 1964
rect -1944 -1964 -1874 1964
rect -1778 -1964 -1708 1964
rect -1612 -1964 -1542 1964
rect -1446 -1964 -1376 1964
rect -1280 -1964 -1210 1964
rect -1114 -1964 -1044 1964
rect -948 -1964 -878 1964
rect -782 -1964 -712 1964
rect -616 -1964 -546 1964
rect -450 -1964 -380 1964
rect -284 -1964 -214 1964
rect -118 -1964 -48 1964
rect 48 -1964 118 1964
rect 214 -1964 284 1964
rect 380 -1964 450 1964
rect 546 -1964 616 1964
rect 712 -1964 782 1964
rect 878 -1964 948 1964
rect 1044 -1964 1114 1964
rect 1210 -1964 1280 1964
rect 1376 -1964 1446 1964
rect 1542 -1964 1612 1964
rect 1708 -1964 1778 1964
rect 1874 -1964 1944 1964
rect 2040 -1964 2110 1964
rect 2206 -1964 2276 1964
<< locali >>
rect -2406 2492 -2310 2526
rect 2310 2492 2406 2526
rect -2406 2430 -2372 2492
rect 2372 2430 2406 2492
rect -2406 -2492 -2372 -2430
rect 2372 -2492 2406 -2430
rect -2406 -2526 -2310 -2492
rect 2310 -2526 2406 -2492
<< viali >>
rect -2260 1981 -2222 2378
rect -2094 1981 -2056 2378
rect -1928 1981 -1890 2378
rect -1762 1981 -1724 2378
rect -1596 1981 -1558 2378
rect -1430 1981 -1392 2378
rect -1264 1981 -1226 2378
rect -1098 1981 -1060 2378
rect -932 1981 -894 2378
rect -766 1981 -728 2378
rect -600 1981 -562 2378
rect -434 1981 -396 2378
rect -268 1981 -230 2378
rect -102 1981 -64 2378
rect 64 1981 102 2378
rect 230 1981 268 2378
rect 396 1981 434 2378
rect 562 1981 600 2378
rect 728 1981 766 2378
rect 894 1981 932 2378
rect 1060 1981 1098 2378
rect 1226 1981 1264 2378
rect 1392 1981 1430 2378
rect 1558 1981 1596 2378
rect 1724 1981 1762 2378
rect 1890 1981 1928 2378
rect 2056 1981 2094 2378
rect 2222 1981 2260 2378
rect -2260 -2378 -2222 -1981
rect -2094 -2378 -2056 -1981
rect -1928 -2378 -1890 -1981
rect -1762 -2378 -1724 -1981
rect -1596 -2378 -1558 -1981
rect -1430 -2378 -1392 -1981
rect -1264 -2378 -1226 -1981
rect -1098 -2378 -1060 -1981
rect -932 -2378 -894 -1981
rect -766 -2378 -728 -1981
rect -600 -2378 -562 -1981
rect -434 -2378 -396 -1981
rect -268 -2378 -230 -1981
rect -102 -2378 -64 -1981
rect 64 -2378 102 -1981
rect 230 -2378 268 -1981
rect 396 -2378 434 -1981
rect 562 -2378 600 -1981
rect 728 -2378 766 -1981
rect 894 -2378 932 -1981
rect 1060 -2378 1098 -1981
rect 1226 -2378 1264 -1981
rect 1392 -2378 1430 -1981
rect 1558 -2378 1596 -1981
rect 1724 -2378 1762 -1981
rect 1890 -2378 1928 -1981
rect 2056 -2378 2094 -1981
rect 2222 -2378 2260 -1981
<< metal1 >>
rect -2266 2378 -2216 2390
rect -2266 1981 -2260 2378
rect -2222 1981 -2216 2378
rect -2266 1969 -2216 1981
rect -2100 2378 -2050 2390
rect -2100 1981 -2094 2378
rect -2056 1981 -2050 2378
rect -2100 1969 -2050 1981
rect -1934 2378 -1884 2390
rect -1934 1981 -1928 2378
rect -1890 1981 -1884 2378
rect -1934 1969 -1884 1981
rect -1768 2378 -1718 2390
rect -1768 1981 -1762 2378
rect -1724 1981 -1718 2378
rect -1768 1969 -1718 1981
rect -1602 2378 -1552 2390
rect -1602 1981 -1596 2378
rect -1558 1981 -1552 2378
rect -1602 1969 -1552 1981
rect -1436 2378 -1386 2390
rect -1436 1981 -1430 2378
rect -1392 1981 -1386 2378
rect -1436 1969 -1386 1981
rect -1270 2378 -1220 2390
rect -1270 1981 -1264 2378
rect -1226 1981 -1220 2378
rect -1270 1969 -1220 1981
rect -1104 2378 -1054 2390
rect -1104 1981 -1098 2378
rect -1060 1981 -1054 2378
rect -1104 1969 -1054 1981
rect -938 2378 -888 2390
rect -938 1981 -932 2378
rect -894 1981 -888 2378
rect -938 1969 -888 1981
rect -772 2378 -722 2390
rect -772 1981 -766 2378
rect -728 1981 -722 2378
rect -772 1969 -722 1981
rect -606 2378 -556 2390
rect -606 1981 -600 2378
rect -562 1981 -556 2378
rect -606 1969 -556 1981
rect -440 2378 -390 2390
rect -440 1981 -434 2378
rect -396 1981 -390 2378
rect -440 1969 -390 1981
rect -274 2378 -224 2390
rect -274 1981 -268 2378
rect -230 1981 -224 2378
rect -274 1969 -224 1981
rect -108 2378 -58 2390
rect -108 1981 -102 2378
rect -64 1981 -58 2378
rect -108 1969 -58 1981
rect 58 2378 108 2390
rect 58 1981 64 2378
rect 102 1981 108 2378
rect 58 1969 108 1981
rect 224 2378 274 2390
rect 224 1981 230 2378
rect 268 1981 274 2378
rect 224 1969 274 1981
rect 390 2378 440 2390
rect 390 1981 396 2378
rect 434 1981 440 2378
rect 390 1969 440 1981
rect 556 2378 606 2390
rect 556 1981 562 2378
rect 600 1981 606 2378
rect 556 1969 606 1981
rect 722 2378 772 2390
rect 722 1981 728 2378
rect 766 1981 772 2378
rect 722 1969 772 1981
rect 888 2378 938 2390
rect 888 1981 894 2378
rect 932 1981 938 2378
rect 888 1969 938 1981
rect 1054 2378 1104 2390
rect 1054 1981 1060 2378
rect 1098 1981 1104 2378
rect 1054 1969 1104 1981
rect 1220 2378 1270 2390
rect 1220 1981 1226 2378
rect 1264 1981 1270 2378
rect 1220 1969 1270 1981
rect 1386 2378 1436 2390
rect 1386 1981 1392 2378
rect 1430 1981 1436 2378
rect 1386 1969 1436 1981
rect 1552 2378 1602 2390
rect 1552 1981 1558 2378
rect 1596 1981 1602 2378
rect 1552 1969 1602 1981
rect 1718 2378 1768 2390
rect 1718 1981 1724 2378
rect 1762 1981 1768 2378
rect 1718 1969 1768 1981
rect 1884 2378 1934 2390
rect 1884 1981 1890 2378
rect 1928 1981 1934 2378
rect 1884 1969 1934 1981
rect 2050 2378 2100 2390
rect 2050 1981 2056 2378
rect 2094 1981 2100 2378
rect 2050 1969 2100 1981
rect 2216 2378 2266 2390
rect 2216 1981 2222 2378
rect 2260 1981 2266 2378
rect 2216 1969 2266 1981
rect -2266 -1981 -2216 -1969
rect -2266 -2378 -2260 -1981
rect -2222 -2378 -2216 -1981
rect -2266 -2390 -2216 -2378
rect -2100 -1981 -2050 -1969
rect -2100 -2378 -2094 -1981
rect -2056 -2378 -2050 -1981
rect -2100 -2390 -2050 -2378
rect -1934 -1981 -1884 -1969
rect -1934 -2378 -1928 -1981
rect -1890 -2378 -1884 -1981
rect -1934 -2390 -1884 -2378
rect -1768 -1981 -1718 -1969
rect -1768 -2378 -1762 -1981
rect -1724 -2378 -1718 -1981
rect -1768 -2390 -1718 -2378
rect -1602 -1981 -1552 -1969
rect -1602 -2378 -1596 -1981
rect -1558 -2378 -1552 -1981
rect -1602 -2390 -1552 -2378
rect -1436 -1981 -1386 -1969
rect -1436 -2378 -1430 -1981
rect -1392 -2378 -1386 -1981
rect -1436 -2390 -1386 -2378
rect -1270 -1981 -1220 -1969
rect -1270 -2378 -1264 -1981
rect -1226 -2378 -1220 -1981
rect -1270 -2390 -1220 -2378
rect -1104 -1981 -1054 -1969
rect -1104 -2378 -1098 -1981
rect -1060 -2378 -1054 -1981
rect -1104 -2390 -1054 -2378
rect -938 -1981 -888 -1969
rect -938 -2378 -932 -1981
rect -894 -2378 -888 -1981
rect -938 -2390 -888 -2378
rect -772 -1981 -722 -1969
rect -772 -2378 -766 -1981
rect -728 -2378 -722 -1981
rect -772 -2390 -722 -2378
rect -606 -1981 -556 -1969
rect -606 -2378 -600 -1981
rect -562 -2378 -556 -1981
rect -606 -2390 -556 -2378
rect -440 -1981 -390 -1969
rect -440 -2378 -434 -1981
rect -396 -2378 -390 -1981
rect -440 -2390 -390 -2378
rect -274 -1981 -224 -1969
rect -274 -2378 -268 -1981
rect -230 -2378 -224 -1981
rect -274 -2390 -224 -2378
rect -108 -1981 -58 -1969
rect -108 -2378 -102 -1981
rect -64 -2378 -58 -1981
rect -108 -2390 -58 -2378
rect 58 -1981 108 -1969
rect 58 -2378 64 -1981
rect 102 -2378 108 -1981
rect 58 -2390 108 -2378
rect 224 -1981 274 -1969
rect 224 -2378 230 -1981
rect 268 -2378 274 -1981
rect 224 -2390 274 -2378
rect 390 -1981 440 -1969
rect 390 -2378 396 -1981
rect 434 -2378 440 -1981
rect 390 -2390 440 -2378
rect 556 -1981 606 -1969
rect 556 -2378 562 -1981
rect 600 -2378 606 -1981
rect 556 -2390 606 -2378
rect 722 -1981 772 -1969
rect 722 -2378 728 -1981
rect 766 -2378 772 -1981
rect 722 -2390 772 -2378
rect 888 -1981 938 -1969
rect 888 -2378 894 -1981
rect 932 -2378 938 -1981
rect 888 -2390 938 -2378
rect 1054 -1981 1104 -1969
rect 1054 -2378 1060 -1981
rect 1098 -2378 1104 -1981
rect 1054 -2390 1104 -2378
rect 1220 -1981 1270 -1969
rect 1220 -2378 1226 -1981
rect 1264 -2378 1270 -1981
rect 1220 -2390 1270 -2378
rect 1386 -1981 1436 -1969
rect 1386 -2378 1392 -1981
rect 1430 -2378 1436 -1981
rect 1386 -2390 1436 -2378
rect 1552 -1981 1602 -1969
rect 1552 -2378 1558 -1981
rect 1596 -2378 1602 -1981
rect 1552 -2390 1602 -2378
rect 1718 -1981 1768 -1969
rect 1718 -2378 1724 -1981
rect 1762 -2378 1768 -1981
rect 1718 -2390 1768 -2378
rect 1884 -1981 1934 -1969
rect 1884 -2378 1890 -1981
rect 1928 -2378 1934 -1981
rect 1884 -2390 1934 -2378
rect 2050 -1981 2100 -1969
rect 2050 -2378 2056 -1981
rect 2094 -2378 2100 -1981
rect 2050 -2390 2100 -2378
rect 2216 -1981 2266 -1969
rect 2216 -2378 2222 -1981
rect 2260 -2378 2266 -1981
rect 2216 -2390 2266 -2378
<< properties >>
string FIXED_BBOX -2389 -2509 2389 2509
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 19.8 m 1 nx 28 wmin 0.350 lmin 0.50 class resistor rho 2000 val 114.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
