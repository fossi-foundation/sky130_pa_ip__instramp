magic
tech sky130A
magscale 1 2
timestamp 1730948043
<< pwell >>
rect -14394 -2052 14394 2052
<< psubdiff >>
rect -14358 1982 -14262 2016
rect 14262 1982 14358 2016
rect -14358 1920 -14324 1982
rect 14324 1920 14358 1982
rect -14358 -1982 -14324 -1920
rect 14324 -1982 14358 -1920
rect -14358 -2016 -14262 -1982
rect 14262 -2016 14358 -1982
<< psubdiffcont >>
rect -14262 1982 14262 2016
rect -14358 -1920 -14324 1920
rect 14324 -1920 14358 1920
rect -14262 -2016 14262 -1982
<< xpolycontact >>
rect -14228 1454 -14158 1886
rect -14228 -1886 -14158 -1454
rect -14062 1454 -13992 1886
rect -14062 -1886 -13992 -1454
rect -13896 1454 -13826 1886
rect -13896 -1886 -13826 -1454
rect -13730 1454 -13660 1886
rect -13730 -1886 -13660 -1454
rect -13564 1454 -13494 1886
rect -13564 -1886 -13494 -1454
rect -13398 1454 -13328 1886
rect -13398 -1886 -13328 -1454
rect -13232 1454 -13162 1886
rect -13232 -1886 -13162 -1454
rect -13066 1454 -12996 1886
rect -13066 -1886 -12996 -1454
rect -12900 1454 -12830 1886
rect -12900 -1886 -12830 -1454
rect -12734 1454 -12664 1886
rect -12734 -1886 -12664 -1454
rect -12568 1454 -12498 1886
rect -12568 -1886 -12498 -1454
rect -12402 1454 -12332 1886
rect -12402 -1886 -12332 -1454
rect -12236 1454 -12166 1886
rect -12236 -1886 -12166 -1454
rect -12070 1454 -12000 1886
rect -12070 -1886 -12000 -1454
rect -11904 1454 -11834 1886
rect -11904 -1886 -11834 -1454
rect -11738 1454 -11668 1886
rect -11738 -1886 -11668 -1454
rect -11572 1454 -11502 1886
rect -11572 -1886 -11502 -1454
rect -11406 1454 -11336 1886
rect -11406 -1886 -11336 -1454
rect -11240 1454 -11170 1886
rect -11240 -1886 -11170 -1454
rect -11074 1454 -11004 1886
rect -11074 -1886 -11004 -1454
rect -10908 1454 -10838 1886
rect -10908 -1886 -10838 -1454
rect -10742 1454 -10672 1886
rect -10742 -1886 -10672 -1454
rect -10576 1454 -10506 1886
rect -10576 -1886 -10506 -1454
rect -10410 1454 -10340 1886
rect -10410 -1886 -10340 -1454
rect -10244 1454 -10174 1886
rect -10244 -1886 -10174 -1454
rect -10078 1454 -10008 1886
rect -10078 -1886 -10008 -1454
rect -9912 1454 -9842 1886
rect -9912 -1886 -9842 -1454
rect -9746 1454 -9676 1886
rect -9746 -1886 -9676 -1454
rect -9580 1454 -9510 1886
rect -9580 -1886 -9510 -1454
rect -9414 1454 -9344 1886
rect -9414 -1886 -9344 -1454
rect -9248 1454 -9178 1886
rect -9248 -1886 -9178 -1454
rect -9082 1454 -9012 1886
rect -9082 -1886 -9012 -1454
rect -8916 1454 -8846 1886
rect -8916 -1886 -8846 -1454
rect -8750 1454 -8680 1886
rect -8750 -1886 -8680 -1454
rect -8584 1454 -8514 1886
rect -8584 -1886 -8514 -1454
rect -8418 1454 -8348 1886
rect -8418 -1886 -8348 -1454
rect -8252 1454 -8182 1886
rect -8252 -1886 -8182 -1454
rect -8086 1454 -8016 1886
rect -8086 -1886 -8016 -1454
rect -7920 1454 -7850 1886
rect -7920 -1886 -7850 -1454
rect -7754 1454 -7684 1886
rect -7754 -1886 -7684 -1454
rect -7588 1454 -7518 1886
rect -7588 -1886 -7518 -1454
rect -7422 1454 -7352 1886
rect -7422 -1886 -7352 -1454
rect -7256 1454 -7186 1886
rect -7256 -1886 -7186 -1454
rect -7090 1454 -7020 1886
rect -7090 -1886 -7020 -1454
rect -6924 1454 -6854 1886
rect -6924 -1886 -6854 -1454
rect -6758 1454 -6688 1886
rect -6758 -1886 -6688 -1454
rect -6592 1454 -6522 1886
rect -6592 -1886 -6522 -1454
rect -6426 1454 -6356 1886
rect -6426 -1886 -6356 -1454
rect -6260 1454 -6190 1886
rect -6260 -1886 -6190 -1454
rect -6094 1454 -6024 1886
rect -6094 -1886 -6024 -1454
rect -5928 1454 -5858 1886
rect -5928 -1886 -5858 -1454
rect -5762 1454 -5692 1886
rect -5762 -1886 -5692 -1454
rect -5596 1454 -5526 1886
rect -5596 -1886 -5526 -1454
rect -5430 1454 -5360 1886
rect -5430 -1886 -5360 -1454
rect -5264 1454 -5194 1886
rect -5264 -1886 -5194 -1454
rect -5098 1454 -5028 1886
rect -5098 -1886 -5028 -1454
rect -4932 1454 -4862 1886
rect -4932 -1886 -4862 -1454
rect -4766 1454 -4696 1886
rect -4766 -1886 -4696 -1454
rect -4600 1454 -4530 1886
rect -4600 -1886 -4530 -1454
rect -4434 1454 -4364 1886
rect -4434 -1886 -4364 -1454
rect -4268 1454 -4198 1886
rect -4268 -1886 -4198 -1454
rect -4102 1454 -4032 1886
rect -4102 -1886 -4032 -1454
rect -3936 1454 -3866 1886
rect -3936 -1886 -3866 -1454
rect -3770 1454 -3700 1886
rect -3770 -1886 -3700 -1454
rect -3604 1454 -3534 1886
rect -3604 -1886 -3534 -1454
rect -3438 1454 -3368 1886
rect -3438 -1886 -3368 -1454
rect -3272 1454 -3202 1886
rect -3272 -1886 -3202 -1454
rect -3106 1454 -3036 1886
rect -3106 -1886 -3036 -1454
rect -2940 1454 -2870 1886
rect -2940 -1886 -2870 -1454
rect -2774 1454 -2704 1886
rect -2774 -1886 -2704 -1454
rect -2608 1454 -2538 1886
rect -2608 -1886 -2538 -1454
rect -2442 1454 -2372 1886
rect -2442 -1886 -2372 -1454
rect -2276 1454 -2206 1886
rect -2276 -1886 -2206 -1454
rect -2110 1454 -2040 1886
rect -2110 -1886 -2040 -1454
rect -1944 1454 -1874 1886
rect -1944 -1886 -1874 -1454
rect -1778 1454 -1708 1886
rect -1778 -1886 -1708 -1454
rect -1612 1454 -1542 1886
rect -1612 -1886 -1542 -1454
rect -1446 1454 -1376 1886
rect -1446 -1886 -1376 -1454
rect -1280 1454 -1210 1886
rect -1280 -1886 -1210 -1454
rect -1114 1454 -1044 1886
rect -1114 -1886 -1044 -1454
rect -948 1454 -878 1886
rect -948 -1886 -878 -1454
rect -782 1454 -712 1886
rect -782 -1886 -712 -1454
rect -616 1454 -546 1886
rect -616 -1886 -546 -1454
rect -450 1454 -380 1886
rect -450 -1886 -380 -1454
rect -284 1454 -214 1886
rect -284 -1886 -214 -1454
rect -118 1454 -48 1886
rect -118 -1886 -48 -1454
rect 48 1454 118 1886
rect 48 -1886 118 -1454
rect 214 1454 284 1886
rect 214 -1886 284 -1454
rect 380 1454 450 1886
rect 380 -1886 450 -1454
rect 546 1454 616 1886
rect 546 -1886 616 -1454
rect 712 1454 782 1886
rect 712 -1886 782 -1454
rect 878 1454 948 1886
rect 878 -1886 948 -1454
rect 1044 1454 1114 1886
rect 1044 -1886 1114 -1454
rect 1210 1454 1280 1886
rect 1210 -1886 1280 -1454
rect 1376 1454 1446 1886
rect 1376 -1886 1446 -1454
rect 1542 1454 1612 1886
rect 1542 -1886 1612 -1454
rect 1708 1454 1778 1886
rect 1708 -1886 1778 -1454
rect 1874 1454 1944 1886
rect 1874 -1886 1944 -1454
rect 2040 1454 2110 1886
rect 2040 -1886 2110 -1454
rect 2206 1454 2276 1886
rect 2206 -1886 2276 -1454
rect 2372 1454 2442 1886
rect 2372 -1886 2442 -1454
rect 2538 1454 2608 1886
rect 2538 -1886 2608 -1454
rect 2704 1454 2774 1886
rect 2704 -1886 2774 -1454
rect 2870 1454 2940 1886
rect 2870 -1886 2940 -1454
rect 3036 1454 3106 1886
rect 3036 -1886 3106 -1454
rect 3202 1454 3272 1886
rect 3202 -1886 3272 -1454
rect 3368 1454 3438 1886
rect 3368 -1886 3438 -1454
rect 3534 1454 3604 1886
rect 3534 -1886 3604 -1454
rect 3700 1454 3770 1886
rect 3700 -1886 3770 -1454
rect 3866 1454 3936 1886
rect 3866 -1886 3936 -1454
rect 4032 1454 4102 1886
rect 4032 -1886 4102 -1454
rect 4198 1454 4268 1886
rect 4198 -1886 4268 -1454
rect 4364 1454 4434 1886
rect 4364 -1886 4434 -1454
rect 4530 1454 4600 1886
rect 4530 -1886 4600 -1454
rect 4696 1454 4766 1886
rect 4696 -1886 4766 -1454
rect 4862 1454 4932 1886
rect 4862 -1886 4932 -1454
rect 5028 1454 5098 1886
rect 5028 -1886 5098 -1454
rect 5194 1454 5264 1886
rect 5194 -1886 5264 -1454
rect 5360 1454 5430 1886
rect 5360 -1886 5430 -1454
rect 5526 1454 5596 1886
rect 5526 -1886 5596 -1454
rect 5692 1454 5762 1886
rect 5692 -1886 5762 -1454
rect 5858 1454 5928 1886
rect 5858 -1886 5928 -1454
rect 6024 1454 6094 1886
rect 6024 -1886 6094 -1454
rect 6190 1454 6260 1886
rect 6190 -1886 6260 -1454
rect 6356 1454 6426 1886
rect 6356 -1886 6426 -1454
rect 6522 1454 6592 1886
rect 6522 -1886 6592 -1454
rect 6688 1454 6758 1886
rect 6688 -1886 6758 -1454
rect 6854 1454 6924 1886
rect 6854 -1886 6924 -1454
rect 7020 1454 7090 1886
rect 7020 -1886 7090 -1454
rect 7186 1454 7256 1886
rect 7186 -1886 7256 -1454
rect 7352 1454 7422 1886
rect 7352 -1886 7422 -1454
rect 7518 1454 7588 1886
rect 7518 -1886 7588 -1454
rect 7684 1454 7754 1886
rect 7684 -1886 7754 -1454
rect 7850 1454 7920 1886
rect 7850 -1886 7920 -1454
rect 8016 1454 8086 1886
rect 8016 -1886 8086 -1454
rect 8182 1454 8252 1886
rect 8182 -1886 8252 -1454
rect 8348 1454 8418 1886
rect 8348 -1886 8418 -1454
rect 8514 1454 8584 1886
rect 8514 -1886 8584 -1454
rect 8680 1454 8750 1886
rect 8680 -1886 8750 -1454
rect 8846 1454 8916 1886
rect 8846 -1886 8916 -1454
rect 9012 1454 9082 1886
rect 9012 -1886 9082 -1454
rect 9178 1454 9248 1886
rect 9178 -1886 9248 -1454
rect 9344 1454 9414 1886
rect 9344 -1886 9414 -1454
rect 9510 1454 9580 1886
rect 9510 -1886 9580 -1454
rect 9676 1454 9746 1886
rect 9676 -1886 9746 -1454
rect 9842 1454 9912 1886
rect 9842 -1886 9912 -1454
rect 10008 1454 10078 1886
rect 10008 -1886 10078 -1454
rect 10174 1454 10244 1886
rect 10174 -1886 10244 -1454
rect 10340 1454 10410 1886
rect 10340 -1886 10410 -1454
rect 10506 1454 10576 1886
rect 10506 -1886 10576 -1454
rect 10672 1454 10742 1886
rect 10672 -1886 10742 -1454
rect 10838 1454 10908 1886
rect 10838 -1886 10908 -1454
rect 11004 1454 11074 1886
rect 11004 -1886 11074 -1454
rect 11170 1454 11240 1886
rect 11170 -1886 11240 -1454
rect 11336 1454 11406 1886
rect 11336 -1886 11406 -1454
rect 11502 1454 11572 1886
rect 11502 -1886 11572 -1454
rect 11668 1454 11738 1886
rect 11668 -1886 11738 -1454
rect 11834 1454 11904 1886
rect 11834 -1886 11904 -1454
rect 12000 1454 12070 1886
rect 12000 -1886 12070 -1454
rect 12166 1454 12236 1886
rect 12166 -1886 12236 -1454
rect 12332 1454 12402 1886
rect 12332 -1886 12402 -1454
rect 12498 1454 12568 1886
rect 12498 -1886 12568 -1454
rect 12664 1454 12734 1886
rect 12664 -1886 12734 -1454
rect 12830 1454 12900 1886
rect 12830 -1886 12900 -1454
rect 12996 1454 13066 1886
rect 12996 -1886 13066 -1454
rect 13162 1454 13232 1886
rect 13162 -1886 13232 -1454
rect 13328 1454 13398 1886
rect 13328 -1886 13398 -1454
rect 13494 1454 13564 1886
rect 13494 -1886 13564 -1454
rect 13660 1454 13730 1886
rect 13660 -1886 13730 -1454
rect 13826 1454 13896 1886
rect 13826 -1886 13896 -1454
rect 13992 1454 14062 1886
rect 13992 -1886 14062 -1454
rect 14158 1454 14228 1886
rect 14158 -1886 14228 -1454
<< xpolyres >>
rect -14228 -1454 -14158 1454
rect -14062 -1454 -13992 1454
rect -13896 -1454 -13826 1454
rect -13730 -1454 -13660 1454
rect -13564 -1454 -13494 1454
rect -13398 -1454 -13328 1454
rect -13232 -1454 -13162 1454
rect -13066 -1454 -12996 1454
rect -12900 -1454 -12830 1454
rect -12734 -1454 -12664 1454
rect -12568 -1454 -12498 1454
rect -12402 -1454 -12332 1454
rect -12236 -1454 -12166 1454
rect -12070 -1454 -12000 1454
rect -11904 -1454 -11834 1454
rect -11738 -1454 -11668 1454
rect -11572 -1454 -11502 1454
rect -11406 -1454 -11336 1454
rect -11240 -1454 -11170 1454
rect -11074 -1454 -11004 1454
rect -10908 -1454 -10838 1454
rect -10742 -1454 -10672 1454
rect -10576 -1454 -10506 1454
rect -10410 -1454 -10340 1454
rect -10244 -1454 -10174 1454
rect -10078 -1454 -10008 1454
rect -9912 -1454 -9842 1454
rect -9746 -1454 -9676 1454
rect -9580 -1454 -9510 1454
rect -9414 -1454 -9344 1454
rect -9248 -1454 -9178 1454
rect -9082 -1454 -9012 1454
rect -8916 -1454 -8846 1454
rect -8750 -1454 -8680 1454
rect -8584 -1454 -8514 1454
rect -8418 -1454 -8348 1454
rect -8252 -1454 -8182 1454
rect -8086 -1454 -8016 1454
rect -7920 -1454 -7850 1454
rect -7754 -1454 -7684 1454
rect -7588 -1454 -7518 1454
rect -7422 -1454 -7352 1454
rect -7256 -1454 -7186 1454
rect -7090 -1454 -7020 1454
rect -6924 -1454 -6854 1454
rect -6758 -1454 -6688 1454
rect -6592 -1454 -6522 1454
rect -6426 -1454 -6356 1454
rect -6260 -1454 -6190 1454
rect -6094 -1454 -6024 1454
rect -5928 -1454 -5858 1454
rect -5762 -1454 -5692 1454
rect -5596 -1454 -5526 1454
rect -5430 -1454 -5360 1454
rect -5264 -1454 -5194 1454
rect -5098 -1454 -5028 1454
rect -4932 -1454 -4862 1454
rect -4766 -1454 -4696 1454
rect -4600 -1454 -4530 1454
rect -4434 -1454 -4364 1454
rect -4268 -1454 -4198 1454
rect -4102 -1454 -4032 1454
rect -3936 -1454 -3866 1454
rect -3770 -1454 -3700 1454
rect -3604 -1454 -3534 1454
rect -3438 -1454 -3368 1454
rect -3272 -1454 -3202 1454
rect -3106 -1454 -3036 1454
rect -2940 -1454 -2870 1454
rect -2774 -1454 -2704 1454
rect -2608 -1454 -2538 1454
rect -2442 -1454 -2372 1454
rect -2276 -1454 -2206 1454
rect -2110 -1454 -2040 1454
rect -1944 -1454 -1874 1454
rect -1778 -1454 -1708 1454
rect -1612 -1454 -1542 1454
rect -1446 -1454 -1376 1454
rect -1280 -1454 -1210 1454
rect -1114 -1454 -1044 1454
rect -948 -1454 -878 1454
rect -782 -1454 -712 1454
rect -616 -1454 -546 1454
rect -450 -1454 -380 1454
rect -284 -1454 -214 1454
rect -118 -1454 -48 1454
rect 48 -1454 118 1454
rect 214 -1454 284 1454
rect 380 -1454 450 1454
rect 546 -1454 616 1454
rect 712 -1454 782 1454
rect 878 -1454 948 1454
rect 1044 -1454 1114 1454
rect 1210 -1454 1280 1454
rect 1376 -1454 1446 1454
rect 1542 -1454 1612 1454
rect 1708 -1454 1778 1454
rect 1874 -1454 1944 1454
rect 2040 -1454 2110 1454
rect 2206 -1454 2276 1454
rect 2372 -1454 2442 1454
rect 2538 -1454 2608 1454
rect 2704 -1454 2774 1454
rect 2870 -1454 2940 1454
rect 3036 -1454 3106 1454
rect 3202 -1454 3272 1454
rect 3368 -1454 3438 1454
rect 3534 -1454 3604 1454
rect 3700 -1454 3770 1454
rect 3866 -1454 3936 1454
rect 4032 -1454 4102 1454
rect 4198 -1454 4268 1454
rect 4364 -1454 4434 1454
rect 4530 -1454 4600 1454
rect 4696 -1454 4766 1454
rect 4862 -1454 4932 1454
rect 5028 -1454 5098 1454
rect 5194 -1454 5264 1454
rect 5360 -1454 5430 1454
rect 5526 -1454 5596 1454
rect 5692 -1454 5762 1454
rect 5858 -1454 5928 1454
rect 6024 -1454 6094 1454
rect 6190 -1454 6260 1454
rect 6356 -1454 6426 1454
rect 6522 -1454 6592 1454
rect 6688 -1454 6758 1454
rect 6854 -1454 6924 1454
rect 7020 -1454 7090 1454
rect 7186 -1454 7256 1454
rect 7352 -1454 7422 1454
rect 7518 -1454 7588 1454
rect 7684 -1454 7754 1454
rect 7850 -1454 7920 1454
rect 8016 -1454 8086 1454
rect 8182 -1454 8252 1454
rect 8348 -1454 8418 1454
rect 8514 -1454 8584 1454
rect 8680 -1454 8750 1454
rect 8846 -1454 8916 1454
rect 9012 -1454 9082 1454
rect 9178 -1454 9248 1454
rect 9344 -1454 9414 1454
rect 9510 -1454 9580 1454
rect 9676 -1454 9746 1454
rect 9842 -1454 9912 1454
rect 10008 -1454 10078 1454
rect 10174 -1454 10244 1454
rect 10340 -1454 10410 1454
rect 10506 -1454 10576 1454
rect 10672 -1454 10742 1454
rect 10838 -1454 10908 1454
rect 11004 -1454 11074 1454
rect 11170 -1454 11240 1454
rect 11336 -1454 11406 1454
rect 11502 -1454 11572 1454
rect 11668 -1454 11738 1454
rect 11834 -1454 11904 1454
rect 12000 -1454 12070 1454
rect 12166 -1454 12236 1454
rect 12332 -1454 12402 1454
rect 12498 -1454 12568 1454
rect 12664 -1454 12734 1454
rect 12830 -1454 12900 1454
rect 12996 -1454 13066 1454
rect 13162 -1454 13232 1454
rect 13328 -1454 13398 1454
rect 13494 -1454 13564 1454
rect 13660 -1454 13730 1454
rect 13826 -1454 13896 1454
rect 13992 -1454 14062 1454
rect 14158 -1454 14228 1454
<< locali >>
rect -14358 1982 -14262 2016
rect 14262 1982 14358 2016
rect -14358 1920 -14324 1982
rect 14324 1920 14358 1982
rect -14358 -1982 -14324 -1920
rect 14324 -1982 14358 -1920
rect -14358 -2016 -14262 -1982
rect 14262 -2016 14358 -1982
<< viali >>
rect -14212 1471 -14174 1868
rect -14046 1471 -14008 1868
rect -13880 1471 -13842 1868
rect -13714 1471 -13676 1868
rect -13548 1471 -13510 1868
rect -13382 1471 -13344 1868
rect -13216 1471 -13178 1868
rect -13050 1471 -13012 1868
rect -12884 1471 -12846 1868
rect -12718 1471 -12680 1868
rect -12552 1471 -12514 1868
rect -12386 1471 -12348 1868
rect -12220 1471 -12182 1868
rect -12054 1471 -12016 1868
rect -11888 1471 -11850 1868
rect -11722 1471 -11684 1868
rect -11556 1471 -11518 1868
rect -11390 1471 -11352 1868
rect -11224 1471 -11186 1868
rect -11058 1471 -11020 1868
rect -10892 1471 -10854 1868
rect -10726 1471 -10688 1868
rect -10560 1471 -10522 1868
rect -10394 1471 -10356 1868
rect -10228 1471 -10190 1868
rect -10062 1471 -10024 1868
rect -9896 1471 -9858 1868
rect -9730 1471 -9692 1868
rect -9564 1471 -9526 1868
rect -9398 1471 -9360 1868
rect -9232 1471 -9194 1868
rect -9066 1471 -9028 1868
rect -8900 1471 -8862 1868
rect -8734 1471 -8696 1868
rect -8568 1471 -8530 1868
rect -8402 1471 -8364 1868
rect -8236 1471 -8198 1868
rect -8070 1471 -8032 1868
rect -7904 1471 -7866 1868
rect -7738 1471 -7700 1868
rect -7572 1471 -7534 1868
rect -7406 1471 -7368 1868
rect -7240 1471 -7202 1868
rect -7074 1471 -7036 1868
rect -6908 1471 -6870 1868
rect -6742 1471 -6704 1868
rect -6576 1471 -6538 1868
rect -6410 1471 -6372 1868
rect -6244 1471 -6206 1868
rect -6078 1471 -6040 1868
rect -5912 1471 -5874 1868
rect -5746 1471 -5708 1868
rect -5580 1471 -5542 1868
rect -5414 1471 -5376 1868
rect -5248 1471 -5210 1868
rect -5082 1471 -5044 1868
rect -4916 1471 -4878 1868
rect -4750 1471 -4712 1868
rect -4584 1471 -4546 1868
rect -4418 1471 -4380 1868
rect -4252 1471 -4214 1868
rect -4086 1471 -4048 1868
rect -3920 1471 -3882 1868
rect -3754 1471 -3716 1868
rect -3588 1471 -3550 1868
rect -3422 1471 -3384 1868
rect -3256 1471 -3218 1868
rect -3090 1471 -3052 1868
rect -2924 1471 -2886 1868
rect -2758 1471 -2720 1868
rect -2592 1471 -2554 1868
rect -2426 1471 -2388 1868
rect -2260 1471 -2222 1868
rect -2094 1471 -2056 1868
rect -1928 1471 -1890 1868
rect -1762 1471 -1724 1868
rect -1596 1471 -1558 1868
rect -1430 1471 -1392 1868
rect -1264 1471 -1226 1868
rect -1098 1471 -1060 1868
rect -932 1471 -894 1868
rect -766 1471 -728 1868
rect -600 1471 -562 1868
rect -434 1471 -396 1868
rect -268 1471 -230 1868
rect -102 1471 -64 1868
rect 64 1471 102 1868
rect 230 1471 268 1868
rect 396 1471 434 1868
rect 562 1471 600 1868
rect 728 1471 766 1868
rect 894 1471 932 1868
rect 1060 1471 1098 1868
rect 1226 1471 1264 1868
rect 1392 1471 1430 1868
rect 1558 1471 1596 1868
rect 1724 1471 1762 1868
rect 1890 1471 1928 1868
rect 2056 1471 2094 1868
rect 2222 1471 2260 1868
rect 2388 1471 2426 1868
rect 2554 1471 2592 1868
rect 2720 1471 2758 1868
rect 2886 1471 2924 1868
rect 3052 1471 3090 1868
rect 3218 1471 3256 1868
rect 3384 1471 3422 1868
rect 3550 1471 3588 1868
rect 3716 1471 3754 1868
rect 3882 1471 3920 1868
rect 4048 1471 4086 1868
rect 4214 1471 4252 1868
rect 4380 1471 4418 1868
rect 4546 1471 4584 1868
rect 4712 1471 4750 1868
rect 4878 1471 4916 1868
rect 5044 1471 5082 1868
rect 5210 1471 5248 1868
rect 5376 1471 5414 1868
rect 5542 1471 5580 1868
rect 5708 1471 5746 1868
rect 5874 1471 5912 1868
rect 6040 1471 6078 1868
rect 6206 1471 6244 1868
rect 6372 1471 6410 1868
rect 6538 1471 6576 1868
rect 6704 1471 6742 1868
rect 6870 1471 6908 1868
rect 7036 1471 7074 1868
rect 7202 1471 7240 1868
rect 7368 1471 7406 1868
rect 7534 1471 7572 1868
rect 7700 1471 7738 1868
rect 7866 1471 7904 1868
rect 8032 1471 8070 1868
rect 8198 1471 8236 1868
rect 8364 1471 8402 1868
rect 8530 1471 8568 1868
rect 8696 1471 8734 1868
rect 8862 1471 8900 1868
rect 9028 1471 9066 1868
rect 9194 1471 9232 1868
rect 9360 1471 9398 1868
rect 9526 1471 9564 1868
rect 9692 1471 9730 1868
rect 9858 1471 9896 1868
rect 10024 1471 10062 1868
rect 10190 1471 10228 1868
rect 10356 1471 10394 1868
rect 10522 1471 10560 1868
rect 10688 1471 10726 1868
rect 10854 1471 10892 1868
rect 11020 1471 11058 1868
rect 11186 1471 11224 1868
rect 11352 1471 11390 1868
rect 11518 1471 11556 1868
rect 11684 1471 11722 1868
rect 11850 1471 11888 1868
rect 12016 1471 12054 1868
rect 12182 1471 12220 1868
rect 12348 1471 12386 1868
rect 12514 1471 12552 1868
rect 12680 1471 12718 1868
rect 12846 1471 12884 1868
rect 13012 1471 13050 1868
rect 13178 1471 13216 1868
rect 13344 1471 13382 1868
rect 13510 1471 13548 1868
rect 13676 1471 13714 1868
rect 13842 1471 13880 1868
rect 14008 1471 14046 1868
rect 14174 1471 14212 1868
rect -14212 -1868 -14174 -1471
rect -14046 -1868 -14008 -1471
rect -13880 -1868 -13842 -1471
rect -13714 -1868 -13676 -1471
rect -13548 -1868 -13510 -1471
rect -13382 -1868 -13344 -1471
rect -13216 -1868 -13178 -1471
rect -13050 -1868 -13012 -1471
rect -12884 -1868 -12846 -1471
rect -12718 -1868 -12680 -1471
rect -12552 -1868 -12514 -1471
rect -12386 -1868 -12348 -1471
rect -12220 -1868 -12182 -1471
rect -12054 -1868 -12016 -1471
rect -11888 -1868 -11850 -1471
rect -11722 -1868 -11684 -1471
rect -11556 -1868 -11518 -1471
rect -11390 -1868 -11352 -1471
rect -11224 -1868 -11186 -1471
rect -11058 -1868 -11020 -1471
rect -10892 -1868 -10854 -1471
rect -10726 -1868 -10688 -1471
rect -10560 -1868 -10522 -1471
rect -10394 -1868 -10356 -1471
rect -10228 -1868 -10190 -1471
rect -10062 -1868 -10024 -1471
rect -9896 -1868 -9858 -1471
rect -9730 -1868 -9692 -1471
rect -9564 -1868 -9526 -1471
rect -9398 -1868 -9360 -1471
rect -9232 -1868 -9194 -1471
rect -9066 -1868 -9028 -1471
rect -8900 -1868 -8862 -1471
rect -8734 -1868 -8696 -1471
rect -8568 -1868 -8530 -1471
rect -8402 -1868 -8364 -1471
rect -8236 -1868 -8198 -1471
rect -8070 -1868 -8032 -1471
rect -7904 -1868 -7866 -1471
rect -7738 -1868 -7700 -1471
rect -7572 -1868 -7534 -1471
rect -7406 -1868 -7368 -1471
rect -7240 -1868 -7202 -1471
rect -7074 -1868 -7036 -1471
rect -6908 -1868 -6870 -1471
rect -6742 -1868 -6704 -1471
rect -6576 -1868 -6538 -1471
rect -6410 -1868 -6372 -1471
rect -6244 -1868 -6206 -1471
rect -6078 -1868 -6040 -1471
rect -5912 -1868 -5874 -1471
rect -5746 -1868 -5708 -1471
rect -5580 -1868 -5542 -1471
rect -5414 -1868 -5376 -1471
rect -5248 -1868 -5210 -1471
rect -5082 -1868 -5044 -1471
rect -4916 -1868 -4878 -1471
rect -4750 -1868 -4712 -1471
rect -4584 -1868 -4546 -1471
rect -4418 -1868 -4380 -1471
rect -4252 -1868 -4214 -1471
rect -4086 -1868 -4048 -1471
rect -3920 -1868 -3882 -1471
rect -3754 -1868 -3716 -1471
rect -3588 -1868 -3550 -1471
rect -3422 -1868 -3384 -1471
rect -3256 -1868 -3218 -1471
rect -3090 -1868 -3052 -1471
rect -2924 -1868 -2886 -1471
rect -2758 -1868 -2720 -1471
rect -2592 -1868 -2554 -1471
rect -2426 -1868 -2388 -1471
rect -2260 -1868 -2222 -1471
rect -2094 -1868 -2056 -1471
rect -1928 -1868 -1890 -1471
rect -1762 -1868 -1724 -1471
rect -1596 -1868 -1558 -1471
rect -1430 -1868 -1392 -1471
rect -1264 -1868 -1226 -1471
rect -1098 -1868 -1060 -1471
rect -932 -1868 -894 -1471
rect -766 -1868 -728 -1471
rect -600 -1868 -562 -1471
rect -434 -1868 -396 -1471
rect -268 -1868 -230 -1471
rect -102 -1868 -64 -1471
rect 64 -1868 102 -1471
rect 230 -1868 268 -1471
rect 396 -1868 434 -1471
rect 562 -1868 600 -1471
rect 728 -1868 766 -1471
rect 894 -1868 932 -1471
rect 1060 -1868 1098 -1471
rect 1226 -1868 1264 -1471
rect 1392 -1868 1430 -1471
rect 1558 -1868 1596 -1471
rect 1724 -1868 1762 -1471
rect 1890 -1868 1928 -1471
rect 2056 -1868 2094 -1471
rect 2222 -1868 2260 -1471
rect 2388 -1868 2426 -1471
rect 2554 -1868 2592 -1471
rect 2720 -1868 2758 -1471
rect 2886 -1868 2924 -1471
rect 3052 -1868 3090 -1471
rect 3218 -1868 3256 -1471
rect 3384 -1868 3422 -1471
rect 3550 -1868 3588 -1471
rect 3716 -1868 3754 -1471
rect 3882 -1868 3920 -1471
rect 4048 -1868 4086 -1471
rect 4214 -1868 4252 -1471
rect 4380 -1868 4418 -1471
rect 4546 -1868 4584 -1471
rect 4712 -1868 4750 -1471
rect 4878 -1868 4916 -1471
rect 5044 -1868 5082 -1471
rect 5210 -1868 5248 -1471
rect 5376 -1868 5414 -1471
rect 5542 -1868 5580 -1471
rect 5708 -1868 5746 -1471
rect 5874 -1868 5912 -1471
rect 6040 -1868 6078 -1471
rect 6206 -1868 6244 -1471
rect 6372 -1868 6410 -1471
rect 6538 -1868 6576 -1471
rect 6704 -1868 6742 -1471
rect 6870 -1868 6908 -1471
rect 7036 -1868 7074 -1471
rect 7202 -1868 7240 -1471
rect 7368 -1868 7406 -1471
rect 7534 -1868 7572 -1471
rect 7700 -1868 7738 -1471
rect 7866 -1868 7904 -1471
rect 8032 -1868 8070 -1471
rect 8198 -1868 8236 -1471
rect 8364 -1868 8402 -1471
rect 8530 -1868 8568 -1471
rect 8696 -1868 8734 -1471
rect 8862 -1868 8900 -1471
rect 9028 -1868 9066 -1471
rect 9194 -1868 9232 -1471
rect 9360 -1868 9398 -1471
rect 9526 -1868 9564 -1471
rect 9692 -1868 9730 -1471
rect 9858 -1868 9896 -1471
rect 10024 -1868 10062 -1471
rect 10190 -1868 10228 -1471
rect 10356 -1868 10394 -1471
rect 10522 -1868 10560 -1471
rect 10688 -1868 10726 -1471
rect 10854 -1868 10892 -1471
rect 11020 -1868 11058 -1471
rect 11186 -1868 11224 -1471
rect 11352 -1868 11390 -1471
rect 11518 -1868 11556 -1471
rect 11684 -1868 11722 -1471
rect 11850 -1868 11888 -1471
rect 12016 -1868 12054 -1471
rect 12182 -1868 12220 -1471
rect 12348 -1868 12386 -1471
rect 12514 -1868 12552 -1471
rect 12680 -1868 12718 -1471
rect 12846 -1868 12884 -1471
rect 13012 -1868 13050 -1471
rect 13178 -1868 13216 -1471
rect 13344 -1868 13382 -1471
rect 13510 -1868 13548 -1471
rect 13676 -1868 13714 -1471
rect 13842 -1868 13880 -1471
rect 14008 -1868 14046 -1471
rect 14174 -1868 14212 -1471
<< metal1 >>
rect -14218 1868 -14168 1880
rect -14218 1471 -14212 1868
rect -14174 1471 -14168 1868
rect -14218 1459 -14168 1471
rect -14052 1868 -14002 1880
rect -14052 1471 -14046 1868
rect -14008 1471 -14002 1868
rect -14052 1459 -14002 1471
rect -13886 1868 -13836 1880
rect -13886 1471 -13880 1868
rect -13842 1471 -13836 1868
rect -13886 1459 -13836 1471
rect -13720 1868 -13670 1880
rect -13720 1471 -13714 1868
rect -13676 1471 -13670 1868
rect -13720 1459 -13670 1471
rect -13554 1868 -13504 1880
rect -13554 1471 -13548 1868
rect -13510 1471 -13504 1868
rect -13554 1459 -13504 1471
rect -13388 1868 -13338 1880
rect -13388 1471 -13382 1868
rect -13344 1471 -13338 1868
rect -13388 1459 -13338 1471
rect -13222 1868 -13172 1880
rect -13222 1471 -13216 1868
rect -13178 1471 -13172 1868
rect -13222 1459 -13172 1471
rect -13056 1868 -13006 1880
rect -13056 1471 -13050 1868
rect -13012 1471 -13006 1868
rect -13056 1459 -13006 1471
rect -12890 1868 -12840 1880
rect -12890 1471 -12884 1868
rect -12846 1471 -12840 1868
rect -12890 1459 -12840 1471
rect -12724 1868 -12674 1880
rect -12724 1471 -12718 1868
rect -12680 1471 -12674 1868
rect -12724 1459 -12674 1471
rect -12558 1868 -12508 1880
rect -12558 1471 -12552 1868
rect -12514 1471 -12508 1868
rect -12558 1459 -12508 1471
rect -12392 1868 -12342 1880
rect -12392 1471 -12386 1868
rect -12348 1471 -12342 1868
rect -12392 1459 -12342 1471
rect -12226 1868 -12176 1880
rect -12226 1471 -12220 1868
rect -12182 1471 -12176 1868
rect -12226 1459 -12176 1471
rect -12060 1868 -12010 1880
rect -12060 1471 -12054 1868
rect -12016 1471 -12010 1868
rect -12060 1459 -12010 1471
rect -11894 1868 -11844 1880
rect -11894 1471 -11888 1868
rect -11850 1471 -11844 1868
rect -11894 1459 -11844 1471
rect -11728 1868 -11678 1880
rect -11728 1471 -11722 1868
rect -11684 1471 -11678 1868
rect -11728 1459 -11678 1471
rect -11562 1868 -11512 1880
rect -11562 1471 -11556 1868
rect -11518 1471 -11512 1868
rect -11562 1459 -11512 1471
rect -11396 1868 -11346 1880
rect -11396 1471 -11390 1868
rect -11352 1471 -11346 1868
rect -11396 1459 -11346 1471
rect -11230 1868 -11180 1880
rect -11230 1471 -11224 1868
rect -11186 1471 -11180 1868
rect -11230 1459 -11180 1471
rect -11064 1868 -11014 1880
rect -11064 1471 -11058 1868
rect -11020 1471 -11014 1868
rect -11064 1459 -11014 1471
rect -10898 1868 -10848 1880
rect -10898 1471 -10892 1868
rect -10854 1471 -10848 1868
rect -10898 1459 -10848 1471
rect -10732 1868 -10682 1880
rect -10732 1471 -10726 1868
rect -10688 1471 -10682 1868
rect -10732 1459 -10682 1471
rect -10566 1868 -10516 1880
rect -10566 1471 -10560 1868
rect -10522 1471 -10516 1868
rect -10566 1459 -10516 1471
rect -10400 1868 -10350 1880
rect -10400 1471 -10394 1868
rect -10356 1471 -10350 1868
rect -10400 1459 -10350 1471
rect -10234 1868 -10184 1880
rect -10234 1471 -10228 1868
rect -10190 1471 -10184 1868
rect -10234 1459 -10184 1471
rect -10068 1868 -10018 1880
rect -10068 1471 -10062 1868
rect -10024 1471 -10018 1868
rect -10068 1459 -10018 1471
rect -9902 1868 -9852 1880
rect -9902 1471 -9896 1868
rect -9858 1471 -9852 1868
rect -9902 1459 -9852 1471
rect -9736 1868 -9686 1880
rect -9736 1471 -9730 1868
rect -9692 1471 -9686 1868
rect -9736 1459 -9686 1471
rect -9570 1868 -9520 1880
rect -9570 1471 -9564 1868
rect -9526 1471 -9520 1868
rect -9570 1459 -9520 1471
rect -9404 1868 -9354 1880
rect -9404 1471 -9398 1868
rect -9360 1471 -9354 1868
rect -9404 1459 -9354 1471
rect -9238 1868 -9188 1880
rect -9238 1471 -9232 1868
rect -9194 1471 -9188 1868
rect -9238 1459 -9188 1471
rect -9072 1868 -9022 1880
rect -9072 1471 -9066 1868
rect -9028 1471 -9022 1868
rect -9072 1459 -9022 1471
rect -8906 1868 -8856 1880
rect -8906 1471 -8900 1868
rect -8862 1471 -8856 1868
rect -8906 1459 -8856 1471
rect -8740 1868 -8690 1880
rect -8740 1471 -8734 1868
rect -8696 1471 -8690 1868
rect -8740 1459 -8690 1471
rect -8574 1868 -8524 1880
rect -8574 1471 -8568 1868
rect -8530 1471 -8524 1868
rect -8574 1459 -8524 1471
rect -8408 1868 -8358 1880
rect -8408 1471 -8402 1868
rect -8364 1471 -8358 1868
rect -8408 1459 -8358 1471
rect -8242 1868 -8192 1880
rect -8242 1471 -8236 1868
rect -8198 1471 -8192 1868
rect -8242 1459 -8192 1471
rect -8076 1868 -8026 1880
rect -8076 1471 -8070 1868
rect -8032 1471 -8026 1868
rect -8076 1459 -8026 1471
rect -7910 1868 -7860 1880
rect -7910 1471 -7904 1868
rect -7866 1471 -7860 1868
rect -7910 1459 -7860 1471
rect -7744 1868 -7694 1880
rect -7744 1471 -7738 1868
rect -7700 1471 -7694 1868
rect -7744 1459 -7694 1471
rect -7578 1868 -7528 1880
rect -7578 1471 -7572 1868
rect -7534 1471 -7528 1868
rect -7578 1459 -7528 1471
rect -7412 1868 -7362 1880
rect -7412 1471 -7406 1868
rect -7368 1471 -7362 1868
rect -7412 1459 -7362 1471
rect -7246 1868 -7196 1880
rect -7246 1471 -7240 1868
rect -7202 1471 -7196 1868
rect -7246 1459 -7196 1471
rect -7080 1868 -7030 1880
rect -7080 1471 -7074 1868
rect -7036 1471 -7030 1868
rect -7080 1459 -7030 1471
rect -6914 1868 -6864 1880
rect -6914 1471 -6908 1868
rect -6870 1471 -6864 1868
rect -6914 1459 -6864 1471
rect -6748 1868 -6698 1880
rect -6748 1471 -6742 1868
rect -6704 1471 -6698 1868
rect -6748 1459 -6698 1471
rect -6582 1868 -6532 1880
rect -6582 1471 -6576 1868
rect -6538 1471 -6532 1868
rect -6582 1459 -6532 1471
rect -6416 1868 -6366 1880
rect -6416 1471 -6410 1868
rect -6372 1471 -6366 1868
rect -6416 1459 -6366 1471
rect -6250 1868 -6200 1880
rect -6250 1471 -6244 1868
rect -6206 1471 -6200 1868
rect -6250 1459 -6200 1471
rect -6084 1868 -6034 1880
rect -6084 1471 -6078 1868
rect -6040 1471 -6034 1868
rect -6084 1459 -6034 1471
rect -5918 1868 -5868 1880
rect -5918 1471 -5912 1868
rect -5874 1471 -5868 1868
rect -5918 1459 -5868 1471
rect -5752 1868 -5702 1880
rect -5752 1471 -5746 1868
rect -5708 1471 -5702 1868
rect -5752 1459 -5702 1471
rect -5586 1868 -5536 1880
rect -5586 1471 -5580 1868
rect -5542 1471 -5536 1868
rect -5586 1459 -5536 1471
rect -5420 1868 -5370 1880
rect -5420 1471 -5414 1868
rect -5376 1471 -5370 1868
rect -5420 1459 -5370 1471
rect -5254 1868 -5204 1880
rect -5254 1471 -5248 1868
rect -5210 1471 -5204 1868
rect -5254 1459 -5204 1471
rect -5088 1868 -5038 1880
rect -5088 1471 -5082 1868
rect -5044 1471 -5038 1868
rect -5088 1459 -5038 1471
rect -4922 1868 -4872 1880
rect -4922 1471 -4916 1868
rect -4878 1471 -4872 1868
rect -4922 1459 -4872 1471
rect -4756 1868 -4706 1880
rect -4756 1471 -4750 1868
rect -4712 1471 -4706 1868
rect -4756 1459 -4706 1471
rect -4590 1868 -4540 1880
rect -4590 1471 -4584 1868
rect -4546 1471 -4540 1868
rect -4590 1459 -4540 1471
rect -4424 1868 -4374 1880
rect -4424 1471 -4418 1868
rect -4380 1471 -4374 1868
rect -4424 1459 -4374 1471
rect -4258 1868 -4208 1880
rect -4258 1471 -4252 1868
rect -4214 1471 -4208 1868
rect -4258 1459 -4208 1471
rect -4092 1868 -4042 1880
rect -4092 1471 -4086 1868
rect -4048 1471 -4042 1868
rect -4092 1459 -4042 1471
rect -3926 1868 -3876 1880
rect -3926 1471 -3920 1868
rect -3882 1471 -3876 1868
rect -3926 1459 -3876 1471
rect -3760 1868 -3710 1880
rect -3760 1471 -3754 1868
rect -3716 1471 -3710 1868
rect -3760 1459 -3710 1471
rect -3594 1868 -3544 1880
rect -3594 1471 -3588 1868
rect -3550 1471 -3544 1868
rect -3594 1459 -3544 1471
rect -3428 1868 -3378 1880
rect -3428 1471 -3422 1868
rect -3384 1471 -3378 1868
rect -3428 1459 -3378 1471
rect -3262 1868 -3212 1880
rect -3262 1471 -3256 1868
rect -3218 1471 -3212 1868
rect -3262 1459 -3212 1471
rect -3096 1868 -3046 1880
rect -3096 1471 -3090 1868
rect -3052 1471 -3046 1868
rect -3096 1459 -3046 1471
rect -2930 1868 -2880 1880
rect -2930 1471 -2924 1868
rect -2886 1471 -2880 1868
rect -2930 1459 -2880 1471
rect -2764 1868 -2714 1880
rect -2764 1471 -2758 1868
rect -2720 1471 -2714 1868
rect -2764 1459 -2714 1471
rect -2598 1868 -2548 1880
rect -2598 1471 -2592 1868
rect -2554 1471 -2548 1868
rect -2598 1459 -2548 1471
rect -2432 1868 -2382 1880
rect -2432 1471 -2426 1868
rect -2388 1471 -2382 1868
rect -2432 1459 -2382 1471
rect -2266 1868 -2216 1880
rect -2266 1471 -2260 1868
rect -2222 1471 -2216 1868
rect -2266 1459 -2216 1471
rect -2100 1868 -2050 1880
rect -2100 1471 -2094 1868
rect -2056 1471 -2050 1868
rect -2100 1459 -2050 1471
rect -1934 1868 -1884 1880
rect -1934 1471 -1928 1868
rect -1890 1471 -1884 1868
rect -1934 1459 -1884 1471
rect -1768 1868 -1718 1880
rect -1768 1471 -1762 1868
rect -1724 1471 -1718 1868
rect -1768 1459 -1718 1471
rect -1602 1868 -1552 1880
rect -1602 1471 -1596 1868
rect -1558 1471 -1552 1868
rect -1602 1459 -1552 1471
rect -1436 1868 -1386 1880
rect -1436 1471 -1430 1868
rect -1392 1471 -1386 1868
rect -1436 1459 -1386 1471
rect -1270 1868 -1220 1880
rect -1270 1471 -1264 1868
rect -1226 1471 -1220 1868
rect -1270 1459 -1220 1471
rect -1104 1868 -1054 1880
rect -1104 1471 -1098 1868
rect -1060 1471 -1054 1868
rect -1104 1459 -1054 1471
rect -938 1868 -888 1880
rect -938 1471 -932 1868
rect -894 1471 -888 1868
rect -938 1459 -888 1471
rect -772 1868 -722 1880
rect -772 1471 -766 1868
rect -728 1471 -722 1868
rect -772 1459 -722 1471
rect -606 1868 -556 1880
rect -606 1471 -600 1868
rect -562 1471 -556 1868
rect -606 1459 -556 1471
rect -440 1868 -390 1880
rect -440 1471 -434 1868
rect -396 1471 -390 1868
rect -440 1459 -390 1471
rect -274 1868 -224 1880
rect -274 1471 -268 1868
rect -230 1471 -224 1868
rect -274 1459 -224 1471
rect -108 1868 -58 1880
rect -108 1471 -102 1868
rect -64 1471 -58 1868
rect -108 1459 -58 1471
rect 58 1868 108 1880
rect 58 1471 64 1868
rect 102 1471 108 1868
rect 58 1459 108 1471
rect 224 1868 274 1880
rect 224 1471 230 1868
rect 268 1471 274 1868
rect 224 1459 274 1471
rect 390 1868 440 1880
rect 390 1471 396 1868
rect 434 1471 440 1868
rect 390 1459 440 1471
rect 556 1868 606 1880
rect 556 1471 562 1868
rect 600 1471 606 1868
rect 556 1459 606 1471
rect 722 1868 772 1880
rect 722 1471 728 1868
rect 766 1471 772 1868
rect 722 1459 772 1471
rect 888 1868 938 1880
rect 888 1471 894 1868
rect 932 1471 938 1868
rect 888 1459 938 1471
rect 1054 1868 1104 1880
rect 1054 1471 1060 1868
rect 1098 1471 1104 1868
rect 1054 1459 1104 1471
rect 1220 1868 1270 1880
rect 1220 1471 1226 1868
rect 1264 1471 1270 1868
rect 1220 1459 1270 1471
rect 1386 1868 1436 1880
rect 1386 1471 1392 1868
rect 1430 1471 1436 1868
rect 1386 1459 1436 1471
rect 1552 1868 1602 1880
rect 1552 1471 1558 1868
rect 1596 1471 1602 1868
rect 1552 1459 1602 1471
rect 1718 1868 1768 1880
rect 1718 1471 1724 1868
rect 1762 1471 1768 1868
rect 1718 1459 1768 1471
rect 1884 1868 1934 1880
rect 1884 1471 1890 1868
rect 1928 1471 1934 1868
rect 1884 1459 1934 1471
rect 2050 1868 2100 1880
rect 2050 1471 2056 1868
rect 2094 1471 2100 1868
rect 2050 1459 2100 1471
rect 2216 1868 2266 1880
rect 2216 1471 2222 1868
rect 2260 1471 2266 1868
rect 2216 1459 2266 1471
rect 2382 1868 2432 1880
rect 2382 1471 2388 1868
rect 2426 1471 2432 1868
rect 2382 1459 2432 1471
rect 2548 1868 2598 1880
rect 2548 1471 2554 1868
rect 2592 1471 2598 1868
rect 2548 1459 2598 1471
rect 2714 1868 2764 1880
rect 2714 1471 2720 1868
rect 2758 1471 2764 1868
rect 2714 1459 2764 1471
rect 2880 1868 2930 1880
rect 2880 1471 2886 1868
rect 2924 1471 2930 1868
rect 2880 1459 2930 1471
rect 3046 1868 3096 1880
rect 3046 1471 3052 1868
rect 3090 1471 3096 1868
rect 3046 1459 3096 1471
rect 3212 1868 3262 1880
rect 3212 1471 3218 1868
rect 3256 1471 3262 1868
rect 3212 1459 3262 1471
rect 3378 1868 3428 1880
rect 3378 1471 3384 1868
rect 3422 1471 3428 1868
rect 3378 1459 3428 1471
rect 3544 1868 3594 1880
rect 3544 1471 3550 1868
rect 3588 1471 3594 1868
rect 3544 1459 3594 1471
rect 3710 1868 3760 1880
rect 3710 1471 3716 1868
rect 3754 1471 3760 1868
rect 3710 1459 3760 1471
rect 3876 1868 3926 1880
rect 3876 1471 3882 1868
rect 3920 1471 3926 1868
rect 3876 1459 3926 1471
rect 4042 1868 4092 1880
rect 4042 1471 4048 1868
rect 4086 1471 4092 1868
rect 4042 1459 4092 1471
rect 4208 1868 4258 1880
rect 4208 1471 4214 1868
rect 4252 1471 4258 1868
rect 4208 1459 4258 1471
rect 4374 1868 4424 1880
rect 4374 1471 4380 1868
rect 4418 1471 4424 1868
rect 4374 1459 4424 1471
rect 4540 1868 4590 1880
rect 4540 1471 4546 1868
rect 4584 1471 4590 1868
rect 4540 1459 4590 1471
rect 4706 1868 4756 1880
rect 4706 1471 4712 1868
rect 4750 1471 4756 1868
rect 4706 1459 4756 1471
rect 4872 1868 4922 1880
rect 4872 1471 4878 1868
rect 4916 1471 4922 1868
rect 4872 1459 4922 1471
rect 5038 1868 5088 1880
rect 5038 1471 5044 1868
rect 5082 1471 5088 1868
rect 5038 1459 5088 1471
rect 5204 1868 5254 1880
rect 5204 1471 5210 1868
rect 5248 1471 5254 1868
rect 5204 1459 5254 1471
rect 5370 1868 5420 1880
rect 5370 1471 5376 1868
rect 5414 1471 5420 1868
rect 5370 1459 5420 1471
rect 5536 1868 5586 1880
rect 5536 1471 5542 1868
rect 5580 1471 5586 1868
rect 5536 1459 5586 1471
rect 5702 1868 5752 1880
rect 5702 1471 5708 1868
rect 5746 1471 5752 1868
rect 5702 1459 5752 1471
rect 5868 1868 5918 1880
rect 5868 1471 5874 1868
rect 5912 1471 5918 1868
rect 5868 1459 5918 1471
rect 6034 1868 6084 1880
rect 6034 1471 6040 1868
rect 6078 1471 6084 1868
rect 6034 1459 6084 1471
rect 6200 1868 6250 1880
rect 6200 1471 6206 1868
rect 6244 1471 6250 1868
rect 6200 1459 6250 1471
rect 6366 1868 6416 1880
rect 6366 1471 6372 1868
rect 6410 1471 6416 1868
rect 6366 1459 6416 1471
rect 6532 1868 6582 1880
rect 6532 1471 6538 1868
rect 6576 1471 6582 1868
rect 6532 1459 6582 1471
rect 6698 1868 6748 1880
rect 6698 1471 6704 1868
rect 6742 1471 6748 1868
rect 6698 1459 6748 1471
rect 6864 1868 6914 1880
rect 6864 1471 6870 1868
rect 6908 1471 6914 1868
rect 6864 1459 6914 1471
rect 7030 1868 7080 1880
rect 7030 1471 7036 1868
rect 7074 1471 7080 1868
rect 7030 1459 7080 1471
rect 7196 1868 7246 1880
rect 7196 1471 7202 1868
rect 7240 1471 7246 1868
rect 7196 1459 7246 1471
rect 7362 1868 7412 1880
rect 7362 1471 7368 1868
rect 7406 1471 7412 1868
rect 7362 1459 7412 1471
rect 7528 1868 7578 1880
rect 7528 1471 7534 1868
rect 7572 1471 7578 1868
rect 7528 1459 7578 1471
rect 7694 1868 7744 1880
rect 7694 1471 7700 1868
rect 7738 1471 7744 1868
rect 7694 1459 7744 1471
rect 7860 1868 7910 1880
rect 7860 1471 7866 1868
rect 7904 1471 7910 1868
rect 7860 1459 7910 1471
rect 8026 1868 8076 1880
rect 8026 1471 8032 1868
rect 8070 1471 8076 1868
rect 8026 1459 8076 1471
rect 8192 1868 8242 1880
rect 8192 1471 8198 1868
rect 8236 1471 8242 1868
rect 8192 1459 8242 1471
rect 8358 1868 8408 1880
rect 8358 1471 8364 1868
rect 8402 1471 8408 1868
rect 8358 1459 8408 1471
rect 8524 1868 8574 1880
rect 8524 1471 8530 1868
rect 8568 1471 8574 1868
rect 8524 1459 8574 1471
rect 8690 1868 8740 1880
rect 8690 1471 8696 1868
rect 8734 1471 8740 1868
rect 8690 1459 8740 1471
rect 8856 1868 8906 1880
rect 8856 1471 8862 1868
rect 8900 1471 8906 1868
rect 8856 1459 8906 1471
rect 9022 1868 9072 1880
rect 9022 1471 9028 1868
rect 9066 1471 9072 1868
rect 9022 1459 9072 1471
rect 9188 1868 9238 1880
rect 9188 1471 9194 1868
rect 9232 1471 9238 1868
rect 9188 1459 9238 1471
rect 9354 1868 9404 1880
rect 9354 1471 9360 1868
rect 9398 1471 9404 1868
rect 9354 1459 9404 1471
rect 9520 1868 9570 1880
rect 9520 1471 9526 1868
rect 9564 1471 9570 1868
rect 9520 1459 9570 1471
rect 9686 1868 9736 1880
rect 9686 1471 9692 1868
rect 9730 1471 9736 1868
rect 9686 1459 9736 1471
rect 9852 1868 9902 1880
rect 9852 1471 9858 1868
rect 9896 1471 9902 1868
rect 9852 1459 9902 1471
rect 10018 1868 10068 1880
rect 10018 1471 10024 1868
rect 10062 1471 10068 1868
rect 10018 1459 10068 1471
rect 10184 1868 10234 1880
rect 10184 1471 10190 1868
rect 10228 1471 10234 1868
rect 10184 1459 10234 1471
rect 10350 1868 10400 1880
rect 10350 1471 10356 1868
rect 10394 1471 10400 1868
rect 10350 1459 10400 1471
rect 10516 1868 10566 1880
rect 10516 1471 10522 1868
rect 10560 1471 10566 1868
rect 10516 1459 10566 1471
rect 10682 1868 10732 1880
rect 10682 1471 10688 1868
rect 10726 1471 10732 1868
rect 10682 1459 10732 1471
rect 10848 1868 10898 1880
rect 10848 1471 10854 1868
rect 10892 1471 10898 1868
rect 10848 1459 10898 1471
rect 11014 1868 11064 1880
rect 11014 1471 11020 1868
rect 11058 1471 11064 1868
rect 11014 1459 11064 1471
rect 11180 1868 11230 1880
rect 11180 1471 11186 1868
rect 11224 1471 11230 1868
rect 11180 1459 11230 1471
rect 11346 1868 11396 1880
rect 11346 1471 11352 1868
rect 11390 1471 11396 1868
rect 11346 1459 11396 1471
rect 11512 1868 11562 1880
rect 11512 1471 11518 1868
rect 11556 1471 11562 1868
rect 11512 1459 11562 1471
rect 11678 1868 11728 1880
rect 11678 1471 11684 1868
rect 11722 1471 11728 1868
rect 11678 1459 11728 1471
rect 11844 1868 11894 1880
rect 11844 1471 11850 1868
rect 11888 1471 11894 1868
rect 11844 1459 11894 1471
rect 12010 1868 12060 1880
rect 12010 1471 12016 1868
rect 12054 1471 12060 1868
rect 12010 1459 12060 1471
rect 12176 1868 12226 1880
rect 12176 1471 12182 1868
rect 12220 1471 12226 1868
rect 12176 1459 12226 1471
rect 12342 1868 12392 1880
rect 12342 1471 12348 1868
rect 12386 1471 12392 1868
rect 12342 1459 12392 1471
rect 12508 1868 12558 1880
rect 12508 1471 12514 1868
rect 12552 1471 12558 1868
rect 12508 1459 12558 1471
rect 12674 1868 12724 1880
rect 12674 1471 12680 1868
rect 12718 1471 12724 1868
rect 12674 1459 12724 1471
rect 12840 1868 12890 1880
rect 12840 1471 12846 1868
rect 12884 1471 12890 1868
rect 12840 1459 12890 1471
rect 13006 1868 13056 1880
rect 13006 1471 13012 1868
rect 13050 1471 13056 1868
rect 13006 1459 13056 1471
rect 13172 1868 13222 1880
rect 13172 1471 13178 1868
rect 13216 1471 13222 1868
rect 13172 1459 13222 1471
rect 13338 1868 13388 1880
rect 13338 1471 13344 1868
rect 13382 1471 13388 1868
rect 13338 1459 13388 1471
rect 13504 1868 13554 1880
rect 13504 1471 13510 1868
rect 13548 1471 13554 1868
rect 13504 1459 13554 1471
rect 13670 1868 13720 1880
rect 13670 1471 13676 1868
rect 13714 1471 13720 1868
rect 13670 1459 13720 1471
rect 13836 1868 13886 1880
rect 13836 1471 13842 1868
rect 13880 1471 13886 1868
rect 13836 1459 13886 1471
rect 14002 1868 14052 1880
rect 14002 1471 14008 1868
rect 14046 1471 14052 1868
rect 14002 1459 14052 1471
rect 14168 1868 14218 1880
rect 14168 1471 14174 1868
rect 14212 1471 14218 1868
rect 14168 1459 14218 1471
rect -14218 -1471 -14168 -1459
rect -14218 -1868 -14212 -1471
rect -14174 -1868 -14168 -1471
rect -14218 -1880 -14168 -1868
rect -14052 -1471 -14002 -1459
rect -14052 -1868 -14046 -1471
rect -14008 -1868 -14002 -1471
rect -14052 -1880 -14002 -1868
rect -13886 -1471 -13836 -1459
rect -13886 -1868 -13880 -1471
rect -13842 -1868 -13836 -1471
rect -13886 -1880 -13836 -1868
rect -13720 -1471 -13670 -1459
rect -13720 -1868 -13714 -1471
rect -13676 -1868 -13670 -1471
rect -13720 -1880 -13670 -1868
rect -13554 -1471 -13504 -1459
rect -13554 -1868 -13548 -1471
rect -13510 -1868 -13504 -1471
rect -13554 -1880 -13504 -1868
rect -13388 -1471 -13338 -1459
rect -13388 -1868 -13382 -1471
rect -13344 -1868 -13338 -1471
rect -13388 -1880 -13338 -1868
rect -13222 -1471 -13172 -1459
rect -13222 -1868 -13216 -1471
rect -13178 -1868 -13172 -1471
rect -13222 -1880 -13172 -1868
rect -13056 -1471 -13006 -1459
rect -13056 -1868 -13050 -1471
rect -13012 -1868 -13006 -1471
rect -13056 -1880 -13006 -1868
rect -12890 -1471 -12840 -1459
rect -12890 -1868 -12884 -1471
rect -12846 -1868 -12840 -1471
rect -12890 -1880 -12840 -1868
rect -12724 -1471 -12674 -1459
rect -12724 -1868 -12718 -1471
rect -12680 -1868 -12674 -1471
rect -12724 -1880 -12674 -1868
rect -12558 -1471 -12508 -1459
rect -12558 -1868 -12552 -1471
rect -12514 -1868 -12508 -1471
rect -12558 -1880 -12508 -1868
rect -12392 -1471 -12342 -1459
rect -12392 -1868 -12386 -1471
rect -12348 -1868 -12342 -1471
rect -12392 -1880 -12342 -1868
rect -12226 -1471 -12176 -1459
rect -12226 -1868 -12220 -1471
rect -12182 -1868 -12176 -1471
rect -12226 -1880 -12176 -1868
rect -12060 -1471 -12010 -1459
rect -12060 -1868 -12054 -1471
rect -12016 -1868 -12010 -1471
rect -12060 -1880 -12010 -1868
rect -11894 -1471 -11844 -1459
rect -11894 -1868 -11888 -1471
rect -11850 -1868 -11844 -1471
rect -11894 -1880 -11844 -1868
rect -11728 -1471 -11678 -1459
rect -11728 -1868 -11722 -1471
rect -11684 -1868 -11678 -1471
rect -11728 -1880 -11678 -1868
rect -11562 -1471 -11512 -1459
rect -11562 -1868 -11556 -1471
rect -11518 -1868 -11512 -1471
rect -11562 -1880 -11512 -1868
rect -11396 -1471 -11346 -1459
rect -11396 -1868 -11390 -1471
rect -11352 -1868 -11346 -1471
rect -11396 -1880 -11346 -1868
rect -11230 -1471 -11180 -1459
rect -11230 -1868 -11224 -1471
rect -11186 -1868 -11180 -1471
rect -11230 -1880 -11180 -1868
rect -11064 -1471 -11014 -1459
rect -11064 -1868 -11058 -1471
rect -11020 -1868 -11014 -1471
rect -11064 -1880 -11014 -1868
rect -10898 -1471 -10848 -1459
rect -10898 -1868 -10892 -1471
rect -10854 -1868 -10848 -1471
rect -10898 -1880 -10848 -1868
rect -10732 -1471 -10682 -1459
rect -10732 -1868 -10726 -1471
rect -10688 -1868 -10682 -1471
rect -10732 -1880 -10682 -1868
rect -10566 -1471 -10516 -1459
rect -10566 -1868 -10560 -1471
rect -10522 -1868 -10516 -1471
rect -10566 -1880 -10516 -1868
rect -10400 -1471 -10350 -1459
rect -10400 -1868 -10394 -1471
rect -10356 -1868 -10350 -1471
rect -10400 -1880 -10350 -1868
rect -10234 -1471 -10184 -1459
rect -10234 -1868 -10228 -1471
rect -10190 -1868 -10184 -1471
rect -10234 -1880 -10184 -1868
rect -10068 -1471 -10018 -1459
rect -10068 -1868 -10062 -1471
rect -10024 -1868 -10018 -1471
rect -10068 -1880 -10018 -1868
rect -9902 -1471 -9852 -1459
rect -9902 -1868 -9896 -1471
rect -9858 -1868 -9852 -1471
rect -9902 -1880 -9852 -1868
rect -9736 -1471 -9686 -1459
rect -9736 -1868 -9730 -1471
rect -9692 -1868 -9686 -1471
rect -9736 -1880 -9686 -1868
rect -9570 -1471 -9520 -1459
rect -9570 -1868 -9564 -1471
rect -9526 -1868 -9520 -1471
rect -9570 -1880 -9520 -1868
rect -9404 -1471 -9354 -1459
rect -9404 -1868 -9398 -1471
rect -9360 -1868 -9354 -1471
rect -9404 -1880 -9354 -1868
rect -9238 -1471 -9188 -1459
rect -9238 -1868 -9232 -1471
rect -9194 -1868 -9188 -1471
rect -9238 -1880 -9188 -1868
rect -9072 -1471 -9022 -1459
rect -9072 -1868 -9066 -1471
rect -9028 -1868 -9022 -1471
rect -9072 -1880 -9022 -1868
rect -8906 -1471 -8856 -1459
rect -8906 -1868 -8900 -1471
rect -8862 -1868 -8856 -1471
rect -8906 -1880 -8856 -1868
rect -8740 -1471 -8690 -1459
rect -8740 -1868 -8734 -1471
rect -8696 -1868 -8690 -1471
rect -8740 -1880 -8690 -1868
rect -8574 -1471 -8524 -1459
rect -8574 -1868 -8568 -1471
rect -8530 -1868 -8524 -1471
rect -8574 -1880 -8524 -1868
rect -8408 -1471 -8358 -1459
rect -8408 -1868 -8402 -1471
rect -8364 -1868 -8358 -1471
rect -8408 -1880 -8358 -1868
rect -8242 -1471 -8192 -1459
rect -8242 -1868 -8236 -1471
rect -8198 -1868 -8192 -1471
rect -8242 -1880 -8192 -1868
rect -8076 -1471 -8026 -1459
rect -8076 -1868 -8070 -1471
rect -8032 -1868 -8026 -1471
rect -8076 -1880 -8026 -1868
rect -7910 -1471 -7860 -1459
rect -7910 -1868 -7904 -1471
rect -7866 -1868 -7860 -1471
rect -7910 -1880 -7860 -1868
rect -7744 -1471 -7694 -1459
rect -7744 -1868 -7738 -1471
rect -7700 -1868 -7694 -1471
rect -7744 -1880 -7694 -1868
rect -7578 -1471 -7528 -1459
rect -7578 -1868 -7572 -1471
rect -7534 -1868 -7528 -1471
rect -7578 -1880 -7528 -1868
rect -7412 -1471 -7362 -1459
rect -7412 -1868 -7406 -1471
rect -7368 -1868 -7362 -1471
rect -7412 -1880 -7362 -1868
rect -7246 -1471 -7196 -1459
rect -7246 -1868 -7240 -1471
rect -7202 -1868 -7196 -1471
rect -7246 -1880 -7196 -1868
rect -7080 -1471 -7030 -1459
rect -7080 -1868 -7074 -1471
rect -7036 -1868 -7030 -1471
rect -7080 -1880 -7030 -1868
rect -6914 -1471 -6864 -1459
rect -6914 -1868 -6908 -1471
rect -6870 -1868 -6864 -1471
rect -6914 -1880 -6864 -1868
rect -6748 -1471 -6698 -1459
rect -6748 -1868 -6742 -1471
rect -6704 -1868 -6698 -1471
rect -6748 -1880 -6698 -1868
rect -6582 -1471 -6532 -1459
rect -6582 -1868 -6576 -1471
rect -6538 -1868 -6532 -1471
rect -6582 -1880 -6532 -1868
rect -6416 -1471 -6366 -1459
rect -6416 -1868 -6410 -1471
rect -6372 -1868 -6366 -1471
rect -6416 -1880 -6366 -1868
rect -6250 -1471 -6200 -1459
rect -6250 -1868 -6244 -1471
rect -6206 -1868 -6200 -1471
rect -6250 -1880 -6200 -1868
rect -6084 -1471 -6034 -1459
rect -6084 -1868 -6078 -1471
rect -6040 -1868 -6034 -1471
rect -6084 -1880 -6034 -1868
rect -5918 -1471 -5868 -1459
rect -5918 -1868 -5912 -1471
rect -5874 -1868 -5868 -1471
rect -5918 -1880 -5868 -1868
rect -5752 -1471 -5702 -1459
rect -5752 -1868 -5746 -1471
rect -5708 -1868 -5702 -1471
rect -5752 -1880 -5702 -1868
rect -5586 -1471 -5536 -1459
rect -5586 -1868 -5580 -1471
rect -5542 -1868 -5536 -1471
rect -5586 -1880 -5536 -1868
rect -5420 -1471 -5370 -1459
rect -5420 -1868 -5414 -1471
rect -5376 -1868 -5370 -1471
rect -5420 -1880 -5370 -1868
rect -5254 -1471 -5204 -1459
rect -5254 -1868 -5248 -1471
rect -5210 -1868 -5204 -1471
rect -5254 -1880 -5204 -1868
rect -5088 -1471 -5038 -1459
rect -5088 -1868 -5082 -1471
rect -5044 -1868 -5038 -1471
rect -5088 -1880 -5038 -1868
rect -4922 -1471 -4872 -1459
rect -4922 -1868 -4916 -1471
rect -4878 -1868 -4872 -1471
rect -4922 -1880 -4872 -1868
rect -4756 -1471 -4706 -1459
rect -4756 -1868 -4750 -1471
rect -4712 -1868 -4706 -1471
rect -4756 -1880 -4706 -1868
rect -4590 -1471 -4540 -1459
rect -4590 -1868 -4584 -1471
rect -4546 -1868 -4540 -1471
rect -4590 -1880 -4540 -1868
rect -4424 -1471 -4374 -1459
rect -4424 -1868 -4418 -1471
rect -4380 -1868 -4374 -1471
rect -4424 -1880 -4374 -1868
rect -4258 -1471 -4208 -1459
rect -4258 -1868 -4252 -1471
rect -4214 -1868 -4208 -1471
rect -4258 -1880 -4208 -1868
rect -4092 -1471 -4042 -1459
rect -4092 -1868 -4086 -1471
rect -4048 -1868 -4042 -1471
rect -4092 -1880 -4042 -1868
rect -3926 -1471 -3876 -1459
rect -3926 -1868 -3920 -1471
rect -3882 -1868 -3876 -1471
rect -3926 -1880 -3876 -1868
rect -3760 -1471 -3710 -1459
rect -3760 -1868 -3754 -1471
rect -3716 -1868 -3710 -1471
rect -3760 -1880 -3710 -1868
rect -3594 -1471 -3544 -1459
rect -3594 -1868 -3588 -1471
rect -3550 -1868 -3544 -1471
rect -3594 -1880 -3544 -1868
rect -3428 -1471 -3378 -1459
rect -3428 -1868 -3422 -1471
rect -3384 -1868 -3378 -1471
rect -3428 -1880 -3378 -1868
rect -3262 -1471 -3212 -1459
rect -3262 -1868 -3256 -1471
rect -3218 -1868 -3212 -1471
rect -3262 -1880 -3212 -1868
rect -3096 -1471 -3046 -1459
rect -3096 -1868 -3090 -1471
rect -3052 -1868 -3046 -1471
rect -3096 -1880 -3046 -1868
rect -2930 -1471 -2880 -1459
rect -2930 -1868 -2924 -1471
rect -2886 -1868 -2880 -1471
rect -2930 -1880 -2880 -1868
rect -2764 -1471 -2714 -1459
rect -2764 -1868 -2758 -1471
rect -2720 -1868 -2714 -1471
rect -2764 -1880 -2714 -1868
rect -2598 -1471 -2548 -1459
rect -2598 -1868 -2592 -1471
rect -2554 -1868 -2548 -1471
rect -2598 -1880 -2548 -1868
rect -2432 -1471 -2382 -1459
rect -2432 -1868 -2426 -1471
rect -2388 -1868 -2382 -1471
rect -2432 -1880 -2382 -1868
rect -2266 -1471 -2216 -1459
rect -2266 -1868 -2260 -1471
rect -2222 -1868 -2216 -1471
rect -2266 -1880 -2216 -1868
rect -2100 -1471 -2050 -1459
rect -2100 -1868 -2094 -1471
rect -2056 -1868 -2050 -1471
rect -2100 -1880 -2050 -1868
rect -1934 -1471 -1884 -1459
rect -1934 -1868 -1928 -1471
rect -1890 -1868 -1884 -1471
rect -1934 -1880 -1884 -1868
rect -1768 -1471 -1718 -1459
rect -1768 -1868 -1762 -1471
rect -1724 -1868 -1718 -1471
rect -1768 -1880 -1718 -1868
rect -1602 -1471 -1552 -1459
rect -1602 -1868 -1596 -1471
rect -1558 -1868 -1552 -1471
rect -1602 -1880 -1552 -1868
rect -1436 -1471 -1386 -1459
rect -1436 -1868 -1430 -1471
rect -1392 -1868 -1386 -1471
rect -1436 -1880 -1386 -1868
rect -1270 -1471 -1220 -1459
rect -1270 -1868 -1264 -1471
rect -1226 -1868 -1220 -1471
rect -1270 -1880 -1220 -1868
rect -1104 -1471 -1054 -1459
rect -1104 -1868 -1098 -1471
rect -1060 -1868 -1054 -1471
rect -1104 -1880 -1054 -1868
rect -938 -1471 -888 -1459
rect -938 -1868 -932 -1471
rect -894 -1868 -888 -1471
rect -938 -1880 -888 -1868
rect -772 -1471 -722 -1459
rect -772 -1868 -766 -1471
rect -728 -1868 -722 -1471
rect -772 -1880 -722 -1868
rect -606 -1471 -556 -1459
rect -606 -1868 -600 -1471
rect -562 -1868 -556 -1471
rect -606 -1880 -556 -1868
rect -440 -1471 -390 -1459
rect -440 -1868 -434 -1471
rect -396 -1868 -390 -1471
rect -440 -1880 -390 -1868
rect -274 -1471 -224 -1459
rect -274 -1868 -268 -1471
rect -230 -1868 -224 -1471
rect -274 -1880 -224 -1868
rect -108 -1471 -58 -1459
rect -108 -1868 -102 -1471
rect -64 -1868 -58 -1471
rect -108 -1880 -58 -1868
rect 58 -1471 108 -1459
rect 58 -1868 64 -1471
rect 102 -1868 108 -1471
rect 58 -1880 108 -1868
rect 224 -1471 274 -1459
rect 224 -1868 230 -1471
rect 268 -1868 274 -1471
rect 224 -1880 274 -1868
rect 390 -1471 440 -1459
rect 390 -1868 396 -1471
rect 434 -1868 440 -1471
rect 390 -1880 440 -1868
rect 556 -1471 606 -1459
rect 556 -1868 562 -1471
rect 600 -1868 606 -1471
rect 556 -1880 606 -1868
rect 722 -1471 772 -1459
rect 722 -1868 728 -1471
rect 766 -1868 772 -1471
rect 722 -1880 772 -1868
rect 888 -1471 938 -1459
rect 888 -1868 894 -1471
rect 932 -1868 938 -1471
rect 888 -1880 938 -1868
rect 1054 -1471 1104 -1459
rect 1054 -1868 1060 -1471
rect 1098 -1868 1104 -1471
rect 1054 -1880 1104 -1868
rect 1220 -1471 1270 -1459
rect 1220 -1868 1226 -1471
rect 1264 -1868 1270 -1471
rect 1220 -1880 1270 -1868
rect 1386 -1471 1436 -1459
rect 1386 -1868 1392 -1471
rect 1430 -1868 1436 -1471
rect 1386 -1880 1436 -1868
rect 1552 -1471 1602 -1459
rect 1552 -1868 1558 -1471
rect 1596 -1868 1602 -1471
rect 1552 -1880 1602 -1868
rect 1718 -1471 1768 -1459
rect 1718 -1868 1724 -1471
rect 1762 -1868 1768 -1471
rect 1718 -1880 1768 -1868
rect 1884 -1471 1934 -1459
rect 1884 -1868 1890 -1471
rect 1928 -1868 1934 -1471
rect 1884 -1880 1934 -1868
rect 2050 -1471 2100 -1459
rect 2050 -1868 2056 -1471
rect 2094 -1868 2100 -1471
rect 2050 -1880 2100 -1868
rect 2216 -1471 2266 -1459
rect 2216 -1868 2222 -1471
rect 2260 -1868 2266 -1471
rect 2216 -1880 2266 -1868
rect 2382 -1471 2432 -1459
rect 2382 -1868 2388 -1471
rect 2426 -1868 2432 -1471
rect 2382 -1880 2432 -1868
rect 2548 -1471 2598 -1459
rect 2548 -1868 2554 -1471
rect 2592 -1868 2598 -1471
rect 2548 -1880 2598 -1868
rect 2714 -1471 2764 -1459
rect 2714 -1868 2720 -1471
rect 2758 -1868 2764 -1471
rect 2714 -1880 2764 -1868
rect 2880 -1471 2930 -1459
rect 2880 -1868 2886 -1471
rect 2924 -1868 2930 -1471
rect 2880 -1880 2930 -1868
rect 3046 -1471 3096 -1459
rect 3046 -1868 3052 -1471
rect 3090 -1868 3096 -1471
rect 3046 -1880 3096 -1868
rect 3212 -1471 3262 -1459
rect 3212 -1868 3218 -1471
rect 3256 -1868 3262 -1471
rect 3212 -1880 3262 -1868
rect 3378 -1471 3428 -1459
rect 3378 -1868 3384 -1471
rect 3422 -1868 3428 -1471
rect 3378 -1880 3428 -1868
rect 3544 -1471 3594 -1459
rect 3544 -1868 3550 -1471
rect 3588 -1868 3594 -1471
rect 3544 -1880 3594 -1868
rect 3710 -1471 3760 -1459
rect 3710 -1868 3716 -1471
rect 3754 -1868 3760 -1471
rect 3710 -1880 3760 -1868
rect 3876 -1471 3926 -1459
rect 3876 -1868 3882 -1471
rect 3920 -1868 3926 -1471
rect 3876 -1880 3926 -1868
rect 4042 -1471 4092 -1459
rect 4042 -1868 4048 -1471
rect 4086 -1868 4092 -1471
rect 4042 -1880 4092 -1868
rect 4208 -1471 4258 -1459
rect 4208 -1868 4214 -1471
rect 4252 -1868 4258 -1471
rect 4208 -1880 4258 -1868
rect 4374 -1471 4424 -1459
rect 4374 -1868 4380 -1471
rect 4418 -1868 4424 -1471
rect 4374 -1880 4424 -1868
rect 4540 -1471 4590 -1459
rect 4540 -1868 4546 -1471
rect 4584 -1868 4590 -1471
rect 4540 -1880 4590 -1868
rect 4706 -1471 4756 -1459
rect 4706 -1868 4712 -1471
rect 4750 -1868 4756 -1471
rect 4706 -1880 4756 -1868
rect 4872 -1471 4922 -1459
rect 4872 -1868 4878 -1471
rect 4916 -1868 4922 -1471
rect 4872 -1880 4922 -1868
rect 5038 -1471 5088 -1459
rect 5038 -1868 5044 -1471
rect 5082 -1868 5088 -1471
rect 5038 -1880 5088 -1868
rect 5204 -1471 5254 -1459
rect 5204 -1868 5210 -1471
rect 5248 -1868 5254 -1471
rect 5204 -1880 5254 -1868
rect 5370 -1471 5420 -1459
rect 5370 -1868 5376 -1471
rect 5414 -1868 5420 -1471
rect 5370 -1880 5420 -1868
rect 5536 -1471 5586 -1459
rect 5536 -1868 5542 -1471
rect 5580 -1868 5586 -1471
rect 5536 -1880 5586 -1868
rect 5702 -1471 5752 -1459
rect 5702 -1868 5708 -1471
rect 5746 -1868 5752 -1471
rect 5702 -1880 5752 -1868
rect 5868 -1471 5918 -1459
rect 5868 -1868 5874 -1471
rect 5912 -1868 5918 -1471
rect 5868 -1880 5918 -1868
rect 6034 -1471 6084 -1459
rect 6034 -1868 6040 -1471
rect 6078 -1868 6084 -1471
rect 6034 -1880 6084 -1868
rect 6200 -1471 6250 -1459
rect 6200 -1868 6206 -1471
rect 6244 -1868 6250 -1471
rect 6200 -1880 6250 -1868
rect 6366 -1471 6416 -1459
rect 6366 -1868 6372 -1471
rect 6410 -1868 6416 -1471
rect 6366 -1880 6416 -1868
rect 6532 -1471 6582 -1459
rect 6532 -1868 6538 -1471
rect 6576 -1868 6582 -1471
rect 6532 -1880 6582 -1868
rect 6698 -1471 6748 -1459
rect 6698 -1868 6704 -1471
rect 6742 -1868 6748 -1471
rect 6698 -1880 6748 -1868
rect 6864 -1471 6914 -1459
rect 6864 -1868 6870 -1471
rect 6908 -1868 6914 -1471
rect 6864 -1880 6914 -1868
rect 7030 -1471 7080 -1459
rect 7030 -1868 7036 -1471
rect 7074 -1868 7080 -1471
rect 7030 -1880 7080 -1868
rect 7196 -1471 7246 -1459
rect 7196 -1868 7202 -1471
rect 7240 -1868 7246 -1471
rect 7196 -1880 7246 -1868
rect 7362 -1471 7412 -1459
rect 7362 -1868 7368 -1471
rect 7406 -1868 7412 -1471
rect 7362 -1880 7412 -1868
rect 7528 -1471 7578 -1459
rect 7528 -1868 7534 -1471
rect 7572 -1868 7578 -1471
rect 7528 -1880 7578 -1868
rect 7694 -1471 7744 -1459
rect 7694 -1868 7700 -1471
rect 7738 -1868 7744 -1471
rect 7694 -1880 7744 -1868
rect 7860 -1471 7910 -1459
rect 7860 -1868 7866 -1471
rect 7904 -1868 7910 -1471
rect 7860 -1880 7910 -1868
rect 8026 -1471 8076 -1459
rect 8026 -1868 8032 -1471
rect 8070 -1868 8076 -1471
rect 8026 -1880 8076 -1868
rect 8192 -1471 8242 -1459
rect 8192 -1868 8198 -1471
rect 8236 -1868 8242 -1471
rect 8192 -1880 8242 -1868
rect 8358 -1471 8408 -1459
rect 8358 -1868 8364 -1471
rect 8402 -1868 8408 -1471
rect 8358 -1880 8408 -1868
rect 8524 -1471 8574 -1459
rect 8524 -1868 8530 -1471
rect 8568 -1868 8574 -1471
rect 8524 -1880 8574 -1868
rect 8690 -1471 8740 -1459
rect 8690 -1868 8696 -1471
rect 8734 -1868 8740 -1471
rect 8690 -1880 8740 -1868
rect 8856 -1471 8906 -1459
rect 8856 -1868 8862 -1471
rect 8900 -1868 8906 -1471
rect 8856 -1880 8906 -1868
rect 9022 -1471 9072 -1459
rect 9022 -1868 9028 -1471
rect 9066 -1868 9072 -1471
rect 9022 -1880 9072 -1868
rect 9188 -1471 9238 -1459
rect 9188 -1868 9194 -1471
rect 9232 -1868 9238 -1471
rect 9188 -1880 9238 -1868
rect 9354 -1471 9404 -1459
rect 9354 -1868 9360 -1471
rect 9398 -1868 9404 -1471
rect 9354 -1880 9404 -1868
rect 9520 -1471 9570 -1459
rect 9520 -1868 9526 -1471
rect 9564 -1868 9570 -1471
rect 9520 -1880 9570 -1868
rect 9686 -1471 9736 -1459
rect 9686 -1868 9692 -1471
rect 9730 -1868 9736 -1471
rect 9686 -1880 9736 -1868
rect 9852 -1471 9902 -1459
rect 9852 -1868 9858 -1471
rect 9896 -1868 9902 -1471
rect 9852 -1880 9902 -1868
rect 10018 -1471 10068 -1459
rect 10018 -1868 10024 -1471
rect 10062 -1868 10068 -1471
rect 10018 -1880 10068 -1868
rect 10184 -1471 10234 -1459
rect 10184 -1868 10190 -1471
rect 10228 -1868 10234 -1471
rect 10184 -1880 10234 -1868
rect 10350 -1471 10400 -1459
rect 10350 -1868 10356 -1471
rect 10394 -1868 10400 -1471
rect 10350 -1880 10400 -1868
rect 10516 -1471 10566 -1459
rect 10516 -1868 10522 -1471
rect 10560 -1868 10566 -1471
rect 10516 -1880 10566 -1868
rect 10682 -1471 10732 -1459
rect 10682 -1868 10688 -1471
rect 10726 -1868 10732 -1471
rect 10682 -1880 10732 -1868
rect 10848 -1471 10898 -1459
rect 10848 -1868 10854 -1471
rect 10892 -1868 10898 -1471
rect 10848 -1880 10898 -1868
rect 11014 -1471 11064 -1459
rect 11014 -1868 11020 -1471
rect 11058 -1868 11064 -1471
rect 11014 -1880 11064 -1868
rect 11180 -1471 11230 -1459
rect 11180 -1868 11186 -1471
rect 11224 -1868 11230 -1471
rect 11180 -1880 11230 -1868
rect 11346 -1471 11396 -1459
rect 11346 -1868 11352 -1471
rect 11390 -1868 11396 -1471
rect 11346 -1880 11396 -1868
rect 11512 -1471 11562 -1459
rect 11512 -1868 11518 -1471
rect 11556 -1868 11562 -1471
rect 11512 -1880 11562 -1868
rect 11678 -1471 11728 -1459
rect 11678 -1868 11684 -1471
rect 11722 -1868 11728 -1471
rect 11678 -1880 11728 -1868
rect 11844 -1471 11894 -1459
rect 11844 -1868 11850 -1471
rect 11888 -1868 11894 -1471
rect 11844 -1880 11894 -1868
rect 12010 -1471 12060 -1459
rect 12010 -1868 12016 -1471
rect 12054 -1868 12060 -1471
rect 12010 -1880 12060 -1868
rect 12176 -1471 12226 -1459
rect 12176 -1868 12182 -1471
rect 12220 -1868 12226 -1471
rect 12176 -1880 12226 -1868
rect 12342 -1471 12392 -1459
rect 12342 -1868 12348 -1471
rect 12386 -1868 12392 -1471
rect 12342 -1880 12392 -1868
rect 12508 -1471 12558 -1459
rect 12508 -1868 12514 -1471
rect 12552 -1868 12558 -1471
rect 12508 -1880 12558 -1868
rect 12674 -1471 12724 -1459
rect 12674 -1868 12680 -1471
rect 12718 -1868 12724 -1471
rect 12674 -1880 12724 -1868
rect 12840 -1471 12890 -1459
rect 12840 -1868 12846 -1471
rect 12884 -1868 12890 -1471
rect 12840 -1880 12890 -1868
rect 13006 -1471 13056 -1459
rect 13006 -1868 13012 -1471
rect 13050 -1868 13056 -1471
rect 13006 -1880 13056 -1868
rect 13172 -1471 13222 -1459
rect 13172 -1868 13178 -1471
rect 13216 -1868 13222 -1471
rect 13172 -1880 13222 -1868
rect 13338 -1471 13388 -1459
rect 13338 -1868 13344 -1471
rect 13382 -1868 13388 -1471
rect 13338 -1880 13388 -1868
rect 13504 -1471 13554 -1459
rect 13504 -1868 13510 -1471
rect 13548 -1868 13554 -1471
rect 13504 -1880 13554 -1868
rect 13670 -1471 13720 -1459
rect 13670 -1868 13676 -1471
rect 13714 -1868 13720 -1471
rect 13670 -1880 13720 -1868
rect 13836 -1471 13886 -1459
rect 13836 -1868 13842 -1471
rect 13880 -1868 13886 -1471
rect 13836 -1880 13886 -1868
rect 14002 -1471 14052 -1459
rect 14002 -1868 14008 -1471
rect 14046 -1868 14052 -1471
rect 14002 -1880 14052 -1868
rect 14168 -1471 14218 -1459
rect 14168 -1868 14174 -1471
rect 14212 -1868 14218 -1471
rect 14168 -1880 14218 -1868
<< properties >>
string FIXED_BBOX -14341 -1999 14341 1999
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 14.7 m 1 nx 172 wmin 0.350 lmin 0.50 class resistor rho 2000 val 85.075k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
