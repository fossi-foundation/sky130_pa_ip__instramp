magic
tech sky130A
magscale 1 2
timestamp 1730858156
<< pwell >>
rect -14062 -2082 14062 2082
<< psubdiff >>
rect -14026 2012 -13930 2046
rect 13930 2012 14026 2046
rect -14026 1950 -13992 2012
rect 13992 1950 14026 2012
rect -14026 -2012 -13992 -1950
rect 13992 -2012 14026 -1950
rect -14026 -2046 -13930 -2012
rect 13930 -2046 14026 -2012
<< psubdiffcont >>
rect -13930 2012 13930 2046
rect -14026 -1950 -13992 1950
rect 13992 -1950 14026 1950
rect -13930 -2046 13930 -2012
<< xpolycontact >>
rect -13896 1484 -13826 1916
rect -13896 -1916 -13826 -1484
rect -13730 1484 -13660 1916
rect -13730 -1916 -13660 -1484
rect -13564 1484 -13494 1916
rect -13564 -1916 -13494 -1484
rect -13398 1484 -13328 1916
rect -13398 -1916 -13328 -1484
rect -13232 1484 -13162 1916
rect -13232 -1916 -13162 -1484
rect -13066 1484 -12996 1916
rect -13066 -1916 -12996 -1484
rect -12900 1484 -12830 1916
rect -12900 -1916 -12830 -1484
rect -12734 1484 -12664 1916
rect -12734 -1916 -12664 -1484
rect -12568 1484 -12498 1916
rect -12568 -1916 -12498 -1484
rect -12402 1484 -12332 1916
rect -12402 -1916 -12332 -1484
rect -12236 1484 -12166 1916
rect -12236 -1916 -12166 -1484
rect -12070 1484 -12000 1916
rect -12070 -1916 -12000 -1484
rect -11904 1484 -11834 1916
rect -11904 -1916 -11834 -1484
rect -11738 1484 -11668 1916
rect -11738 -1916 -11668 -1484
rect -11572 1484 -11502 1916
rect -11572 -1916 -11502 -1484
rect -11406 1484 -11336 1916
rect -11406 -1916 -11336 -1484
rect -11240 1484 -11170 1916
rect -11240 -1916 -11170 -1484
rect -11074 1484 -11004 1916
rect -11074 -1916 -11004 -1484
rect -10908 1484 -10838 1916
rect -10908 -1916 -10838 -1484
rect -10742 1484 -10672 1916
rect -10742 -1916 -10672 -1484
rect -10576 1484 -10506 1916
rect -10576 -1916 -10506 -1484
rect -10410 1484 -10340 1916
rect -10410 -1916 -10340 -1484
rect -10244 1484 -10174 1916
rect -10244 -1916 -10174 -1484
rect -10078 1484 -10008 1916
rect -10078 -1916 -10008 -1484
rect -9912 1484 -9842 1916
rect -9912 -1916 -9842 -1484
rect -9746 1484 -9676 1916
rect -9746 -1916 -9676 -1484
rect -9580 1484 -9510 1916
rect -9580 -1916 -9510 -1484
rect -9414 1484 -9344 1916
rect -9414 -1916 -9344 -1484
rect -9248 1484 -9178 1916
rect -9248 -1916 -9178 -1484
rect -9082 1484 -9012 1916
rect -9082 -1916 -9012 -1484
rect -8916 1484 -8846 1916
rect -8916 -1916 -8846 -1484
rect -8750 1484 -8680 1916
rect -8750 -1916 -8680 -1484
rect -8584 1484 -8514 1916
rect -8584 -1916 -8514 -1484
rect -8418 1484 -8348 1916
rect -8418 -1916 -8348 -1484
rect -8252 1484 -8182 1916
rect -8252 -1916 -8182 -1484
rect -8086 1484 -8016 1916
rect -8086 -1916 -8016 -1484
rect -7920 1484 -7850 1916
rect -7920 -1916 -7850 -1484
rect -7754 1484 -7684 1916
rect -7754 -1916 -7684 -1484
rect -7588 1484 -7518 1916
rect -7588 -1916 -7518 -1484
rect -7422 1484 -7352 1916
rect -7422 -1916 -7352 -1484
rect -7256 1484 -7186 1916
rect -7256 -1916 -7186 -1484
rect -7090 1484 -7020 1916
rect -7090 -1916 -7020 -1484
rect -6924 1484 -6854 1916
rect -6924 -1916 -6854 -1484
rect -6758 1484 -6688 1916
rect -6758 -1916 -6688 -1484
rect -6592 1484 -6522 1916
rect -6592 -1916 -6522 -1484
rect -6426 1484 -6356 1916
rect -6426 -1916 -6356 -1484
rect -6260 1484 -6190 1916
rect -6260 -1916 -6190 -1484
rect -6094 1484 -6024 1916
rect -6094 -1916 -6024 -1484
rect -5928 1484 -5858 1916
rect -5928 -1916 -5858 -1484
rect -5762 1484 -5692 1916
rect -5762 -1916 -5692 -1484
rect -5596 1484 -5526 1916
rect -5596 -1916 -5526 -1484
rect -5430 1484 -5360 1916
rect -5430 -1916 -5360 -1484
rect -5264 1484 -5194 1916
rect -5264 -1916 -5194 -1484
rect -5098 1484 -5028 1916
rect -5098 -1916 -5028 -1484
rect -4932 1484 -4862 1916
rect -4932 -1916 -4862 -1484
rect -4766 1484 -4696 1916
rect -4766 -1916 -4696 -1484
rect -4600 1484 -4530 1916
rect -4600 -1916 -4530 -1484
rect -4434 1484 -4364 1916
rect -4434 -1916 -4364 -1484
rect -4268 1484 -4198 1916
rect -4268 -1916 -4198 -1484
rect -4102 1484 -4032 1916
rect -4102 -1916 -4032 -1484
rect -3936 1484 -3866 1916
rect -3936 -1916 -3866 -1484
rect -3770 1484 -3700 1916
rect -3770 -1916 -3700 -1484
rect -3604 1484 -3534 1916
rect -3604 -1916 -3534 -1484
rect -3438 1484 -3368 1916
rect -3438 -1916 -3368 -1484
rect -3272 1484 -3202 1916
rect -3272 -1916 -3202 -1484
rect -3106 1484 -3036 1916
rect -3106 -1916 -3036 -1484
rect -2940 1484 -2870 1916
rect -2940 -1916 -2870 -1484
rect -2774 1484 -2704 1916
rect -2774 -1916 -2704 -1484
rect -2608 1484 -2538 1916
rect -2608 -1916 -2538 -1484
rect -2442 1484 -2372 1916
rect -2442 -1916 -2372 -1484
rect -2276 1484 -2206 1916
rect -2276 -1916 -2206 -1484
rect -2110 1484 -2040 1916
rect -2110 -1916 -2040 -1484
rect -1944 1484 -1874 1916
rect -1944 -1916 -1874 -1484
rect -1778 1484 -1708 1916
rect -1778 -1916 -1708 -1484
rect -1612 1484 -1542 1916
rect -1612 -1916 -1542 -1484
rect -1446 1484 -1376 1916
rect -1446 -1916 -1376 -1484
rect -1280 1484 -1210 1916
rect -1280 -1916 -1210 -1484
rect -1114 1484 -1044 1916
rect -1114 -1916 -1044 -1484
rect -948 1484 -878 1916
rect -948 -1916 -878 -1484
rect -782 1484 -712 1916
rect -782 -1916 -712 -1484
rect -616 1484 -546 1916
rect -616 -1916 -546 -1484
rect -450 1484 -380 1916
rect -450 -1916 -380 -1484
rect -284 1484 -214 1916
rect -284 -1916 -214 -1484
rect -118 1484 -48 1916
rect -118 -1916 -48 -1484
rect 48 1484 118 1916
rect 48 -1916 118 -1484
rect 214 1484 284 1916
rect 214 -1916 284 -1484
rect 380 1484 450 1916
rect 380 -1916 450 -1484
rect 546 1484 616 1916
rect 546 -1916 616 -1484
rect 712 1484 782 1916
rect 712 -1916 782 -1484
rect 878 1484 948 1916
rect 878 -1916 948 -1484
rect 1044 1484 1114 1916
rect 1044 -1916 1114 -1484
rect 1210 1484 1280 1916
rect 1210 -1916 1280 -1484
rect 1376 1484 1446 1916
rect 1376 -1916 1446 -1484
rect 1542 1484 1612 1916
rect 1542 -1916 1612 -1484
rect 1708 1484 1778 1916
rect 1708 -1916 1778 -1484
rect 1874 1484 1944 1916
rect 1874 -1916 1944 -1484
rect 2040 1484 2110 1916
rect 2040 -1916 2110 -1484
rect 2206 1484 2276 1916
rect 2206 -1916 2276 -1484
rect 2372 1484 2442 1916
rect 2372 -1916 2442 -1484
rect 2538 1484 2608 1916
rect 2538 -1916 2608 -1484
rect 2704 1484 2774 1916
rect 2704 -1916 2774 -1484
rect 2870 1484 2940 1916
rect 2870 -1916 2940 -1484
rect 3036 1484 3106 1916
rect 3036 -1916 3106 -1484
rect 3202 1484 3272 1916
rect 3202 -1916 3272 -1484
rect 3368 1484 3438 1916
rect 3368 -1916 3438 -1484
rect 3534 1484 3604 1916
rect 3534 -1916 3604 -1484
rect 3700 1484 3770 1916
rect 3700 -1916 3770 -1484
rect 3866 1484 3936 1916
rect 3866 -1916 3936 -1484
rect 4032 1484 4102 1916
rect 4032 -1916 4102 -1484
rect 4198 1484 4268 1916
rect 4198 -1916 4268 -1484
rect 4364 1484 4434 1916
rect 4364 -1916 4434 -1484
rect 4530 1484 4600 1916
rect 4530 -1916 4600 -1484
rect 4696 1484 4766 1916
rect 4696 -1916 4766 -1484
rect 4862 1484 4932 1916
rect 4862 -1916 4932 -1484
rect 5028 1484 5098 1916
rect 5028 -1916 5098 -1484
rect 5194 1484 5264 1916
rect 5194 -1916 5264 -1484
rect 5360 1484 5430 1916
rect 5360 -1916 5430 -1484
rect 5526 1484 5596 1916
rect 5526 -1916 5596 -1484
rect 5692 1484 5762 1916
rect 5692 -1916 5762 -1484
rect 5858 1484 5928 1916
rect 5858 -1916 5928 -1484
rect 6024 1484 6094 1916
rect 6024 -1916 6094 -1484
rect 6190 1484 6260 1916
rect 6190 -1916 6260 -1484
rect 6356 1484 6426 1916
rect 6356 -1916 6426 -1484
rect 6522 1484 6592 1916
rect 6522 -1916 6592 -1484
rect 6688 1484 6758 1916
rect 6688 -1916 6758 -1484
rect 6854 1484 6924 1916
rect 6854 -1916 6924 -1484
rect 7020 1484 7090 1916
rect 7020 -1916 7090 -1484
rect 7186 1484 7256 1916
rect 7186 -1916 7256 -1484
rect 7352 1484 7422 1916
rect 7352 -1916 7422 -1484
rect 7518 1484 7588 1916
rect 7518 -1916 7588 -1484
rect 7684 1484 7754 1916
rect 7684 -1916 7754 -1484
rect 7850 1484 7920 1916
rect 7850 -1916 7920 -1484
rect 8016 1484 8086 1916
rect 8016 -1916 8086 -1484
rect 8182 1484 8252 1916
rect 8182 -1916 8252 -1484
rect 8348 1484 8418 1916
rect 8348 -1916 8418 -1484
rect 8514 1484 8584 1916
rect 8514 -1916 8584 -1484
rect 8680 1484 8750 1916
rect 8680 -1916 8750 -1484
rect 8846 1484 8916 1916
rect 8846 -1916 8916 -1484
rect 9012 1484 9082 1916
rect 9012 -1916 9082 -1484
rect 9178 1484 9248 1916
rect 9178 -1916 9248 -1484
rect 9344 1484 9414 1916
rect 9344 -1916 9414 -1484
rect 9510 1484 9580 1916
rect 9510 -1916 9580 -1484
rect 9676 1484 9746 1916
rect 9676 -1916 9746 -1484
rect 9842 1484 9912 1916
rect 9842 -1916 9912 -1484
rect 10008 1484 10078 1916
rect 10008 -1916 10078 -1484
rect 10174 1484 10244 1916
rect 10174 -1916 10244 -1484
rect 10340 1484 10410 1916
rect 10340 -1916 10410 -1484
rect 10506 1484 10576 1916
rect 10506 -1916 10576 -1484
rect 10672 1484 10742 1916
rect 10672 -1916 10742 -1484
rect 10838 1484 10908 1916
rect 10838 -1916 10908 -1484
rect 11004 1484 11074 1916
rect 11004 -1916 11074 -1484
rect 11170 1484 11240 1916
rect 11170 -1916 11240 -1484
rect 11336 1484 11406 1916
rect 11336 -1916 11406 -1484
rect 11502 1484 11572 1916
rect 11502 -1916 11572 -1484
rect 11668 1484 11738 1916
rect 11668 -1916 11738 -1484
rect 11834 1484 11904 1916
rect 11834 -1916 11904 -1484
rect 12000 1484 12070 1916
rect 12000 -1916 12070 -1484
rect 12166 1484 12236 1916
rect 12166 -1916 12236 -1484
rect 12332 1484 12402 1916
rect 12332 -1916 12402 -1484
rect 12498 1484 12568 1916
rect 12498 -1916 12568 -1484
rect 12664 1484 12734 1916
rect 12664 -1916 12734 -1484
rect 12830 1484 12900 1916
rect 12830 -1916 12900 -1484
rect 12996 1484 13066 1916
rect 12996 -1916 13066 -1484
rect 13162 1484 13232 1916
rect 13162 -1916 13232 -1484
rect 13328 1484 13398 1916
rect 13328 -1916 13398 -1484
rect 13494 1484 13564 1916
rect 13494 -1916 13564 -1484
rect 13660 1484 13730 1916
rect 13660 -1916 13730 -1484
rect 13826 1484 13896 1916
rect 13826 -1916 13896 -1484
<< xpolyres >>
rect -13896 -1484 -13826 1484
rect -13730 -1484 -13660 1484
rect -13564 -1484 -13494 1484
rect -13398 -1484 -13328 1484
rect -13232 -1484 -13162 1484
rect -13066 -1484 -12996 1484
rect -12900 -1484 -12830 1484
rect -12734 -1484 -12664 1484
rect -12568 -1484 -12498 1484
rect -12402 -1484 -12332 1484
rect -12236 -1484 -12166 1484
rect -12070 -1484 -12000 1484
rect -11904 -1484 -11834 1484
rect -11738 -1484 -11668 1484
rect -11572 -1484 -11502 1484
rect -11406 -1484 -11336 1484
rect -11240 -1484 -11170 1484
rect -11074 -1484 -11004 1484
rect -10908 -1484 -10838 1484
rect -10742 -1484 -10672 1484
rect -10576 -1484 -10506 1484
rect -10410 -1484 -10340 1484
rect -10244 -1484 -10174 1484
rect -10078 -1484 -10008 1484
rect -9912 -1484 -9842 1484
rect -9746 -1484 -9676 1484
rect -9580 -1484 -9510 1484
rect -9414 -1484 -9344 1484
rect -9248 -1484 -9178 1484
rect -9082 -1484 -9012 1484
rect -8916 -1484 -8846 1484
rect -8750 -1484 -8680 1484
rect -8584 -1484 -8514 1484
rect -8418 -1484 -8348 1484
rect -8252 -1484 -8182 1484
rect -8086 -1484 -8016 1484
rect -7920 -1484 -7850 1484
rect -7754 -1484 -7684 1484
rect -7588 -1484 -7518 1484
rect -7422 -1484 -7352 1484
rect -7256 -1484 -7186 1484
rect -7090 -1484 -7020 1484
rect -6924 -1484 -6854 1484
rect -6758 -1484 -6688 1484
rect -6592 -1484 -6522 1484
rect -6426 -1484 -6356 1484
rect -6260 -1484 -6190 1484
rect -6094 -1484 -6024 1484
rect -5928 -1484 -5858 1484
rect -5762 -1484 -5692 1484
rect -5596 -1484 -5526 1484
rect -5430 -1484 -5360 1484
rect -5264 -1484 -5194 1484
rect -5098 -1484 -5028 1484
rect -4932 -1484 -4862 1484
rect -4766 -1484 -4696 1484
rect -4600 -1484 -4530 1484
rect -4434 -1484 -4364 1484
rect -4268 -1484 -4198 1484
rect -4102 -1484 -4032 1484
rect -3936 -1484 -3866 1484
rect -3770 -1484 -3700 1484
rect -3604 -1484 -3534 1484
rect -3438 -1484 -3368 1484
rect -3272 -1484 -3202 1484
rect -3106 -1484 -3036 1484
rect -2940 -1484 -2870 1484
rect -2774 -1484 -2704 1484
rect -2608 -1484 -2538 1484
rect -2442 -1484 -2372 1484
rect -2276 -1484 -2206 1484
rect -2110 -1484 -2040 1484
rect -1944 -1484 -1874 1484
rect -1778 -1484 -1708 1484
rect -1612 -1484 -1542 1484
rect -1446 -1484 -1376 1484
rect -1280 -1484 -1210 1484
rect -1114 -1484 -1044 1484
rect -948 -1484 -878 1484
rect -782 -1484 -712 1484
rect -616 -1484 -546 1484
rect -450 -1484 -380 1484
rect -284 -1484 -214 1484
rect -118 -1484 -48 1484
rect 48 -1484 118 1484
rect 214 -1484 284 1484
rect 380 -1484 450 1484
rect 546 -1484 616 1484
rect 712 -1484 782 1484
rect 878 -1484 948 1484
rect 1044 -1484 1114 1484
rect 1210 -1484 1280 1484
rect 1376 -1484 1446 1484
rect 1542 -1484 1612 1484
rect 1708 -1484 1778 1484
rect 1874 -1484 1944 1484
rect 2040 -1484 2110 1484
rect 2206 -1484 2276 1484
rect 2372 -1484 2442 1484
rect 2538 -1484 2608 1484
rect 2704 -1484 2774 1484
rect 2870 -1484 2940 1484
rect 3036 -1484 3106 1484
rect 3202 -1484 3272 1484
rect 3368 -1484 3438 1484
rect 3534 -1484 3604 1484
rect 3700 -1484 3770 1484
rect 3866 -1484 3936 1484
rect 4032 -1484 4102 1484
rect 4198 -1484 4268 1484
rect 4364 -1484 4434 1484
rect 4530 -1484 4600 1484
rect 4696 -1484 4766 1484
rect 4862 -1484 4932 1484
rect 5028 -1484 5098 1484
rect 5194 -1484 5264 1484
rect 5360 -1484 5430 1484
rect 5526 -1484 5596 1484
rect 5692 -1484 5762 1484
rect 5858 -1484 5928 1484
rect 6024 -1484 6094 1484
rect 6190 -1484 6260 1484
rect 6356 -1484 6426 1484
rect 6522 -1484 6592 1484
rect 6688 -1484 6758 1484
rect 6854 -1484 6924 1484
rect 7020 -1484 7090 1484
rect 7186 -1484 7256 1484
rect 7352 -1484 7422 1484
rect 7518 -1484 7588 1484
rect 7684 -1484 7754 1484
rect 7850 -1484 7920 1484
rect 8016 -1484 8086 1484
rect 8182 -1484 8252 1484
rect 8348 -1484 8418 1484
rect 8514 -1484 8584 1484
rect 8680 -1484 8750 1484
rect 8846 -1484 8916 1484
rect 9012 -1484 9082 1484
rect 9178 -1484 9248 1484
rect 9344 -1484 9414 1484
rect 9510 -1484 9580 1484
rect 9676 -1484 9746 1484
rect 9842 -1484 9912 1484
rect 10008 -1484 10078 1484
rect 10174 -1484 10244 1484
rect 10340 -1484 10410 1484
rect 10506 -1484 10576 1484
rect 10672 -1484 10742 1484
rect 10838 -1484 10908 1484
rect 11004 -1484 11074 1484
rect 11170 -1484 11240 1484
rect 11336 -1484 11406 1484
rect 11502 -1484 11572 1484
rect 11668 -1484 11738 1484
rect 11834 -1484 11904 1484
rect 12000 -1484 12070 1484
rect 12166 -1484 12236 1484
rect 12332 -1484 12402 1484
rect 12498 -1484 12568 1484
rect 12664 -1484 12734 1484
rect 12830 -1484 12900 1484
rect 12996 -1484 13066 1484
rect 13162 -1484 13232 1484
rect 13328 -1484 13398 1484
rect 13494 -1484 13564 1484
rect 13660 -1484 13730 1484
rect 13826 -1484 13896 1484
<< locali >>
rect -14026 2012 -13930 2046
rect 13930 2012 14026 2046
rect -14026 1950 -13992 2012
rect 13992 1950 14026 2012
rect -14026 -2012 -13992 -1950
rect 13992 -2012 14026 -1950
rect -14026 -2046 -13930 -2012
rect 13930 -2046 14026 -2012
<< viali >>
rect -13880 1501 -13842 1898
rect -13714 1501 -13676 1898
rect -13548 1501 -13510 1898
rect -13382 1501 -13344 1898
rect -13216 1501 -13178 1898
rect -13050 1501 -13012 1898
rect -12884 1501 -12846 1898
rect -12718 1501 -12680 1898
rect -12552 1501 -12514 1898
rect -12386 1501 -12348 1898
rect -12220 1501 -12182 1898
rect -12054 1501 -12016 1898
rect -11888 1501 -11850 1898
rect -11722 1501 -11684 1898
rect -11556 1501 -11518 1898
rect -11390 1501 -11352 1898
rect -11224 1501 -11186 1898
rect -11058 1501 -11020 1898
rect -10892 1501 -10854 1898
rect -10726 1501 -10688 1898
rect -10560 1501 -10522 1898
rect -10394 1501 -10356 1898
rect -10228 1501 -10190 1898
rect -10062 1501 -10024 1898
rect -9896 1501 -9858 1898
rect -9730 1501 -9692 1898
rect -9564 1501 -9526 1898
rect -9398 1501 -9360 1898
rect -9232 1501 -9194 1898
rect -9066 1501 -9028 1898
rect -8900 1501 -8862 1898
rect -8734 1501 -8696 1898
rect -8568 1501 -8530 1898
rect -8402 1501 -8364 1898
rect -8236 1501 -8198 1898
rect -8070 1501 -8032 1898
rect -7904 1501 -7866 1898
rect -7738 1501 -7700 1898
rect -7572 1501 -7534 1898
rect -7406 1501 -7368 1898
rect -7240 1501 -7202 1898
rect -7074 1501 -7036 1898
rect -6908 1501 -6870 1898
rect -6742 1501 -6704 1898
rect -6576 1501 -6538 1898
rect -6410 1501 -6372 1898
rect -6244 1501 -6206 1898
rect -6078 1501 -6040 1898
rect -5912 1501 -5874 1898
rect -5746 1501 -5708 1898
rect -5580 1501 -5542 1898
rect -5414 1501 -5376 1898
rect -5248 1501 -5210 1898
rect -5082 1501 -5044 1898
rect -4916 1501 -4878 1898
rect -4750 1501 -4712 1898
rect -4584 1501 -4546 1898
rect -4418 1501 -4380 1898
rect -4252 1501 -4214 1898
rect -4086 1501 -4048 1898
rect -3920 1501 -3882 1898
rect -3754 1501 -3716 1898
rect -3588 1501 -3550 1898
rect -3422 1501 -3384 1898
rect -3256 1501 -3218 1898
rect -3090 1501 -3052 1898
rect -2924 1501 -2886 1898
rect -2758 1501 -2720 1898
rect -2592 1501 -2554 1898
rect -2426 1501 -2388 1898
rect -2260 1501 -2222 1898
rect -2094 1501 -2056 1898
rect -1928 1501 -1890 1898
rect -1762 1501 -1724 1898
rect -1596 1501 -1558 1898
rect -1430 1501 -1392 1898
rect -1264 1501 -1226 1898
rect -1098 1501 -1060 1898
rect -932 1501 -894 1898
rect -766 1501 -728 1898
rect -600 1501 -562 1898
rect -434 1501 -396 1898
rect -268 1501 -230 1898
rect -102 1501 -64 1898
rect 64 1501 102 1898
rect 230 1501 268 1898
rect 396 1501 434 1898
rect 562 1501 600 1898
rect 728 1501 766 1898
rect 894 1501 932 1898
rect 1060 1501 1098 1898
rect 1226 1501 1264 1898
rect 1392 1501 1430 1898
rect 1558 1501 1596 1898
rect 1724 1501 1762 1898
rect 1890 1501 1928 1898
rect 2056 1501 2094 1898
rect 2222 1501 2260 1898
rect 2388 1501 2426 1898
rect 2554 1501 2592 1898
rect 2720 1501 2758 1898
rect 2886 1501 2924 1898
rect 3052 1501 3090 1898
rect 3218 1501 3256 1898
rect 3384 1501 3422 1898
rect 3550 1501 3588 1898
rect 3716 1501 3754 1898
rect 3882 1501 3920 1898
rect 4048 1501 4086 1898
rect 4214 1501 4252 1898
rect 4380 1501 4418 1898
rect 4546 1501 4584 1898
rect 4712 1501 4750 1898
rect 4878 1501 4916 1898
rect 5044 1501 5082 1898
rect 5210 1501 5248 1898
rect 5376 1501 5414 1898
rect 5542 1501 5580 1898
rect 5708 1501 5746 1898
rect 5874 1501 5912 1898
rect 6040 1501 6078 1898
rect 6206 1501 6244 1898
rect 6372 1501 6410 1898
rect 6538 1501 6576 1898
rect 6704 1501 6742 1898
rect 6870 1501 6908 1898
rect 7036 1501 7074 1898
rect 7202 1501 7240 1898
rect 7368 1501 7406 1898
rect 7534 1501 7572 1898
rect 7700 1501 7738 1898
rect 7866 1501 7904 1898
rect 8032 1501 8070 1898
rect 8198 1501 8236 1898
rect 8364 1501 8402 1898
rect 8530 1501 8568 1898
rect 8696 1501 8734 1898
rect 8862 1501 8900 1898
rect 9028 1501 9066 1898
rect 9194 1501 9232 1898
rect 9360 1501 9398 1898
rect 9526 1501 9564 1898
rect 9692 1501 9730 1898
rect 9858 1501 9896 1898
rect 10024 1501 10062 1898
rect 10190 1501 10228 1898
rect 10356 1501 10394 1898
rect 10522 1501 10560 1898
rect 10688 1501 10726 1898
rect 10854 1501 10892 1898
rect 11020 1501 11058 1898
rect 11186 1501 11224 1898
rect 11352 1501 11390 1898
rect 11518 1501 11556 1898
rect 11684 1501 11722 1898
rect 11850 1501 11888 1898
rect 12016 1501 12054 1898
rect 12182 1501 12220 1898
rect 12348 1501 12386 1898
rect 12514 1501 12552 1898
rect 12680 1501 12718 1898
rect 12846 1501 12884 1898
rect 13012 1501 13050 1898
rect 13178 1501 13216 1898
rect 13344 1501 13382 1898
rect 13510 1501 13548 1898
rect 13676 1501 13714 1898
rect 13842 1501 13880 1898
rect -13880 -1898 -13842 -1501
rect -13714 -1898 -13676 -1501
rect -13548 -1898 -13510 -1501
rect -13382 -1898 -13344 -1501
rect -13216 -1898 -13178 -1501
rect -13050 -1898 -13012 -1501
rect -12884 -1898 -12846 -1501
rect -12718 -1898 -12680 -1501
rect -12552 -1898 -12514 -1501
rect -12386 -1898 -12348 -1501
rect -12220 -1898 -12182 -1501
rect -12054 -1898 -12016 -1501
rect -11888 -1898 -11850 -1501
rect -11722 -1898 -11684 -1501
rect -11556 -1898 -11518 -1501
rect -11390 -1898 -11352 -1501
rect -11224 -1898 -11186 -1501
rect -11058 -1898 -11020 -1501
rect -10892 -1898 -10854 -1501
rect -10726 -1898 -10688 -1501
rect -10560 -1898 -10522 -1501
rect -10394 -1898 -10356 -1501
rect -10228 -1898 -10190 -1501
rect -10062 -1898 -10024 -1501
rect -9896 -1898 -9858 -1501
rect -9730 -1898 -9692 -1501
rect -9564 -1898 -9526 -1501
rect -9398 -1898 -9360 -1501
rect -9232 -1898 -9194 -1501
rect -9066 -1898 -9028 -1501
rect -8900 -1898 -8862 -1501
rect -8734 -1898 -8696 -1501
rect -8568 -1898 -8530 -1501
rect -8402 -1898 -8364 -1501
rect -8236 -1898 -8198 -1501
rect -8070 -1898 -8032 -1501
rect -7904 -1898 -7866 -1501
rect -7738 -1898 -7700 -1501
rect -7572 -1898 -7534 -1501
rect -7406 -1898 -7368 -1501
rect -7240 -1898 -7202 -1501
rect -7074 -1898 -7036 -1501
rect -6908 -1898 -6870 -1501
rect -6742 -1898 -6704 -1501
rect -6576 -1898 -6538 -1501
rect -6410 -1898 -6372 -1501
rect -6244 -1898 -6206 -1501
rect -6078 -1898 -6040 -1501
rect -5912 -1898 -5874 -1501
rect -5746 -1898 -5708 -1501
rect -5580 -1898 -5542 -1501
rect -5414 -1898 -5376 -1501
rect -5248 -1898 -5210 -1501
rect -5082 -1898 -5044 -1501
rect -4916 -1898 -4878 -1501
rect -4750 -1898 -4712 -1501
rect -4584 -1898 -4546 -1501
rect -4418 -1898 -4380 -1501
rect -4252 -1898 -4214 -1501
rect -4086 -1898 -4048 -1501
rect -3920 -1898 -3882 -1501
rect -3754 -1898 -3716 -1501
rect -3588 -1898 -3550 -1501
rect -3422 -1898 -3384 -1501
rect -3256 -1898 -3218 -1501
rect -3090 -1898 -3052 -1501
rect -2924 -1898 -2886 -1501
rect -2758 -1898 -2720 -1501
rect -2592 -1898 -2554 -1501
rect -2426 -1898 -2388 -1501
rect -2260 -1898 -2222 -1501
rect -2094 -1898 -2056 -1501
rect -1928 -1898 -1890 -1501
rect -1762 -1898 -1724 -1501
rect -1596 -1898 -1558 -1501
rect -1430 -1898 -1392 -1501
rect -1264 -1898 -1226 -1501
rect -1098 -1898 -1060 -1501
rect -932 -1898 -894 -1501
rect -766 -1898 -728 -1501
rect -600 -1898 -562 -1501
rect -434 -1898 -396 -1501
rect -268 -1898 -230 -1501
rect -102 -1898 -64 -1501
rect 64 -1898 102 -1501
rect 230 -1898 268 -1501
rect 396 -1898 434 -1501
rect 562 -1898 600 -1501
rect 728 -1898 766 -1501
rect 894 -1898 932 -1501
rect 1060 -1898 1098 -1501
rect 1226 -1898 1264 -1501
rect 1392 -1898 1430 -1501
rect 1558 -1898 1596 -1501
rect 1724 -1898 1762 -1501
rect 1890 -1898 1928 -1501
rect 2056 -1898 2094 -1501
rect 2222 -1898 2260 -1501
rect 2388 -1898 2426 -1501
rect 2554 -1898 2592 -1501
rect 2720 -1898 2758 -1501
rect 2886 -1898 2924 -1501
rect 3052 -1898 3090 -1501
rect 3218 -1898 3256 -1501
rect 3384 -1898 3422 -1501
rect 3550 -1898 3588 -1501
rect 3716 -1898 3754 -1501
rect 3882 -1898 3920 -1501
rect 4048 -1898 4086 -1501
rect 4214 -1898 4252 -1501
rect 4380 -1898 4418 -1501
rect 4546 -1898 4584 -1501
rect 4712 -1898 4750 -1501
rect 4878 -1898 4916 -1501
rect 5044 -1898 5082 -1501
rect 5210 -1898 5248 -1501
rect 5376 -1898 5414 -1501
rect 5542 -1898 5580 -1501
rect 5708 -1898 5746 -1501
rect 5874 -1898 5912 -1501
rect 6040 -1898 6078 -1501
rect 6206 -1898 6244 -1501
rect 6372 -1898 6410 -1501
rect 6538 -1898 6576 -1501
rect 6704 -1898 6742 -1501
rect 6870 -1898 6908 -1501
rect 7036 -1898 7074 -1501
rect 7202 -1898 7240 -1501
rect 7368 -1898 7406 -1501
rect 7534 -1898 7572 -1501
rect 7700 -1898 7738 -1501
rect 7866 -1898 7904 -1501
rect 8032 -1898 8070 -1501
rect 8198 -1898 8236 -1501
rect 8364 -1898 8402 -1501
rect 8530 -1898 8568 -1501
rect 8696 -1898 8734 -1501
rect 8862 -1898 8900 -1501
rect 9028 -1898 9066 -1501
rect 9194 -1898 9232 -1501
rect 9360 -1898 9398 -1501
rect 9526 -1898 9564 -1501
rect 9692 -1898 9730 -1501
rect 9858 -1898 9896 -1501
rect 10024 -1898 10062 -1501
rect 10190 -1898 10228 -1501
rect 10356 -1898 10394 -1501
rect 10522 -1898 10560 -1501
rect 10688 -1898 10726 -1501
rect 10854 -1898 10892 -1501
rect 11020 -1898 11058 -1501
rect 11186 -1898 11224 -1501
rect 11352 -1898 11390 -1501
rect 11518 -1898 11556 -1501
rect 11684 -1898 11722 -1501
rect 11850 -1898 11888 -1501
rect 12016 -1898 12054 -1501
rect 12182 -1898 12220 -1501
rect 12348 -1898 12386 -1501
rect 12514 -1898 12552 -1501
rect 12680 -1898 12718 -1501
rect 12846 -1898 12884 -1501
rect 13012 -1898 13050 -1501
rect 13178 -1898 13216 -1501
rect 13344 -1898 13382 -1501
rect 13510 -1898 13548 -1501
rect 13676 -1898 13714 -1501
rect 13842 -1898 13880 -1501
<< metal1 >>
rect -13886 1898 -13836 1910
rect -13886 1501 -13880 1898
rect -13842 1501 -13836 1898
rect -13886 1489 -13836 1501
rect -13720 1898 -13670 1910
rect -13720 1501 -13714 1898
rect -13676 1501 -13670 1898
rect -13720 1489 -13670 1501
rect -13554 1898 -13504 1910
rect -13554 1501 -13548 1898
rect -13510 1501 -13504 1898
rect -13554 1489 -13504 1501
rect -13388 1898 -13338 1910
rect -13388 1501 -13382 1898
rect -13344 1501 -13338 1898
rect -13388 1489 -13338 1501
rect -13222 1898 -13172 1910
rect -13222 1501 -13216 1898
rect -13178 1501 -13172 1898
rect -13222 1489 -13172 1501
rect -13056 1898 -13006 1910
rect -13056 1501 -13050 1898
rect -13012 1501 -13006 1898
rect -13056 1489 -13006 1501
rect -12890 1898 -12840 1910
rect -12890 1501 -12884 1898
rect -12846 1501 -12840 1898
rect -12890 1489 -12840 1501
rect -12724 1898 -12674 1910
rect -12724 1501 -12718 1898
rect -12680 1501 -12674 1898
rect -12724 1489 -12674 1501
rect -12558 1898 -12508 1910
rect -12558 1501 -12552 1898
rect -12514 1501 -12508 1898
rect -12558 1489 -12508 1501
rect -12392 1898 -12342 1910
rect -12392 1501 -12386 1898
rect -12348 1501 -12342 1898
rect -12392 1489 -12342 1501
rect -12226 1898 -12176 1910
rect -12226 1501 -12220 1898
rect -12182 1501 -12176 1898
rect -12226 1489 -12176 1501
rect -12060 1898 -12010 1910
rect -12060 1501 -12054 1898
rect -12016 1501 -12010 1898
rect -12060 1489 -12010 1501
rect -11894 1898 -11844 1910
rect -11894 1501 -11888 1898
rect -11850 1501 -11844 1898
rect -11894 1489 -11844 1501
rect -11728 1898 -11678 1910
rect -11728 1501 -11722 1898
rect -11684 1501 -11678 1898
rect -11728 1489 -11678 1501
rect -11562 1898 -11512 1910
rect -11562 1501 -11556 1898
rect -11518 1501 -11512 1898
rect -11562 1489 -11512 1501
rect -11396 1898 -11346 1910
rect -11396 1501 -11390 1898
rect -11352 1501 -11346 1898
rect -11396 1489 -11346 1501
rect -11230 1898 -11180 1910
rect -11230 1501 -11224 1898
rect -11186 1501 -11180 1898
rect -11230 1489 -11180 1501
rect -11064 1898 -11014 1910
rect -11064 1501 -11058 1898
rect -11020 1501 -11014 1898
rect -11064 1489 -11014 1501
rect -10898 1898 -10848 1910
rect -10898 1501 -10892 1898
rect -10854 1501 -10848 1898
rect -10898 1489 -10848 1501
rect -10732 1898 -10682 1910
rect -10732 1501 -10726 1898
rect -10688 1501 -10682 1898
rect -10732 1489 -10682 1501
rect -10566 1898 -10516 1910
rect -10566 1501 -10560 1898
rect -10522 1501 -10516 1898
rect -10566 1489 -10516 1501
rect -10400 1898 -10350 1910
rect -10400 1501 -10394 1898
rect -10356 1501 -10350 1898
rect -10400 1489 -10350 1501
rect -10234 1898 -10184 1910
rect -10234 1501 -10228 1898
rect -10190 1501 -10184 1898
rect -10234 1489 -10184 1501
rect -10068 1898 -10018 1910
rect -10068 1501 -10062 1898
rect -10024 1501 -10018 1898
rect -10068 1489 -10018 1501
rect -9902 1898 -9852 1910
rect -9902 1501 -9896 1898
rect -9858 1501 -9852 1898
rect -9902 1489 -9852 1501
rect -9736 1898 -9686 1910
rect -9736 1501 -9730 1898
rect -9692 1501 -9686 1898
rect -9736 1489 -9686 1501
rect -9570 1898 -9520 1910
rect -9570 1501 -9564 1898
rect -9526 1501 -9520 1898
rect -9570 1489 -9520 1501
rect -9404 1898 -9354 1910
rect -9404 1501 -9398 1898
rect -9360 1501 -9354 1898
rect -9404 1489 -9354 1501
rect -9238 1898 -9188 1910
rect -9238 1501 -9232 1898
rect -9194 1501 -9188 1898
rect -9238 1489 -9188 1501
rect -9072 1898 -9022 1910
rect -9072 1501 -9066 1898
rect -9028 1501 -9022 1898
rect -9072 1489 -9022 1501
rect -8906 1898 -8856 1910
rect -8906 1501 -8900 1898
rect -8862 1501 -8856 1898
rect -8906 1489 -8856 1501
rect -8740 1898 -8690 1910
rect -8740 1501 -8734 1898
rect -8696 1501 -8690 1898
rect -8740 1489 -8690 1501
rect -8574 1898 -8524 1910
rect -8574 1501 -8568 1898
rect -8530 1501 -8524 1898
rect -8574 1489 -8524 1501
rect -8408 1898 -8358 1910
rect -8408 1501 -8402 1898
rect -8364 1501 -8358 1898
rect -8408 1489 -8358 1501
rect -8242 1898 -8192 1910
rect -8242 1501 -8236 1898
rect -8198 1501 -8192 1898
rect -8242 1489 -8192 1501
rect -8076 1898 -8026 1910
rect -8076 1501 -8070 1898
rect -8032 1501 -8026 1898
rect -8076 1489 -8026 1501
rect -7910 1898 -7860 1910
rect -7910 1501 -7904 1898
rect -7866 1501 -7860 1898
rect -7910 1489 -7860 1501
rect -7744 1898 -7694 1910
rect -7744 1501 -7738 1898
rect -7700 1501 -7694 1898
rect -7744 1489 -7694 1501
rect -7578 1898 -7528 1910
rect -7578 1501 -7572 1898
rect -7534 1501 -7528 1898
rect -7578 1489 -7528 1501
rect -7412 1898 -7362 1910
rect -7412 1501 -7406 1898
rect -7368 1501 -7362 1898
rect -7412 1489 -7362 1501
rect -7246 1898 -7196 1910
rect -7246 1501 -7240 1898
rect -7202 1501 -7196 1898
rect -7246 1489 -7196 1501
rect -7080 1898 -7030 1910
rect -7080 1501 -7074 1898
rect -7036 1501 -7030 1898
rect -7080 1489 -7030 1501
rect -6914 1898 -6864 1910
rect -6914 1501 -6908 1898
rect -6870 1501 -6864 1898
rect -6914 1489 -6864 1501
rect -6748 1898 -6698 1910
rect -6748 1501 -6742 1898
rect -6704 1501 -6698 1898
rect -6748 1489 -6698 1501
rect -6582 1898 -6532 1910
rect -6582 1501 -6576 1898
rect -6538 1501 -6532 1898
rect -6582 1489 -6532 1501
rect -6416 1898 -6366 1910
rect -6416 1501 -6410 1898
rect -6372 1501 -6366 1898
rect -6416 1489 -6366 1501
rect -6250 1898 -6200 1910
rect -6250 1501 -6244 1898
rect -6206 1501 -6200 1898
rect -6250 1489 -6200 1501
rect -6084 1898 -6034 1910
rect -6084 1501 -6078 1898
rect -6040 1501 -6034 1898
rect -6084 1489 -6034 1501
rect -5918 1898 -5868 1910
rect -5918 1501 -5912 1898
rect -5874 1501 -5868 1898
rect -5918 1489 -5868 1501
rect -5752 1898 -5702 1910
rect -5752 1501 -5746 1898
rect -5708 1501 -5702 1898
rect -5752 1489 -5702 1501
rect -5586 1898 -5536 1910
rect -5586 1501 -5580 1898
rect -5542 1501 -5536 1898
rect -5586 1489 -5536 1501
rect -5420 1898 -5370 1910
rect -5420 1501 -5414 1898
rect -5376 1501 -5370 1898
rect -5420 1489 -5370 1501
rect -5254 1898 -5204 1910
rect -5254 1501 -5248 1898
rect -5210 1501 -5204 1898
rect -5254 1489 -5204 1501
rect -5088 1898 -5038 1910
rect -5088 1501 -5082 1898
rect -5044 1501 -5038 1898
rect -5088 1489 -5038 1501
rect -4922 1898 -4872 1910
rect -4922 1501 -4916 1898
rect -4878 1501 -4872 1898
rect -4922 1489 -4872 1501
rect -4756 1898 -4706 1910
rect -4756 1501 -4750 1898
rect -4712 1501 -4706 1898
rect -4756 1489 -4706 1501
rect -4590 1898 -4540 1910
rect -4590 1501 -4584 1898
rect -4546 1501 -4540 1898
rect -4590 1489 -4540 1501
rect -4424 1898 -4374 1910
rect -4424 1501 -4418 1898
rect -4380 1501 -4374 1898
rect -4424 1489 -4374 1501
rect -4258 1898 -4208 1910
rect -4258 1501 -4252 1898
rect -4214 1501 -4208 1898
rect -4258 1489 -4208 1501
rect -4092 1898 -4042 1910
rect -4092 1501 -4086 1898
rect -4048 1501 -4042 1898
rect -4092 1489 -4042 1501
rect -3926 1898 -3876 1910
rect -3926 1501 -3920 1898
rect -3882 1501 -3876 1898
rect -3926 1489 -3876 1501
rect -3760 1898 -3710 1910
rect -3760 1501 -3754 1898
rect -3716 1501 -3710 1898
rect -3760 1489 -3710 1501
rect -3594 1898 -3544 1910
rect -3594 1501 -3588 1898
rect -3550 1501 -3544 1898
rect -3594 1489 -3544 1501
rect -3428 1898 -3378 1910
rect -3428 1501 -3422 1898
rect -3384 1501 -3378 1898
rect -3428 1489 -3378 1501
rect -3262 1898 -3212 1910
rect -3262 1501 -3256 1898
rect -3218 1501 -3212 1898
rect -3262 1489 -3212 1501
rect -3096 1898 -3046 1910
rect -3096 1501 -3090 1898
rect -3052 1501 -3046 1898
rect -3096 1489 -3046 1501
rect -2930 1898 -2880 1910
rect -2930 1501 -2924 1898
rect -2886 1501 -2880 1898
rect -2930 1489 -2880 1501
rect -2764 1898 -2714 1910
rect -2764 1501 -2758 1898
rect -2720 1501 -2714 1898
rect -2764 1489 -2714 1501
rect -2598 1898 -2548 1910
rect -2598 1501 -2592 1898
rect -2554 1501 -2548 1898
rect -2598 1489 -2548 1501
rect -2432 1898 -2382 1910
rect -2432 1501 -2426 1898
rect -2388 1501 -2382 1898
rect -2432 1489 -2382 1501
rect -2266 1898 -2216 1910
rect -2266 1501 -2260 1898
rect -2222 1501 -2216 1898
rect -2266 1489 -2216 1501
rect -2100 1898 -2050 1910
rect -2100 1501 -2094 1898
rect -2056 1501 -2050 1898
rect -2100 1489 -2050 1501
rect -1934 1898 -1884 1910
rect -1934 1501 -1928 1898
rect -1890 1501 -1884 1898
rect -1934 1489 -1884 1501
rect -1768 1898 -1718 1910
rect -1768 1501 -1762 1898
rect -1724 1501 -1718 1898
rect -1768 1489 -1718 1501
rect -1602 1898 -1552 1910
rect -1602 1501 -1596 1898
rect -1558 1501 -1552 1898
rect -1602 1489 -1552 1501
rect -1436 1898 -1386 1910
rect -1436 1501 -1430 1898
rect -1392 1501 -1386 1898
rect -1436 1489 -1386 1501
rect -1270 1898 -1220 1910
rect -1270 1501 -1264 1898
rect -1226 1501 -1220 1898
rect -1270 1489 -1220 1501
rect -1104 1898 -1054 1910
rect -1104 1501 -1098 1898
rect -1060 1501 -1054 1898
rect -1104 1489 -1054 1501
rect -938 1898 -888 1910
rect -938 1501 -932 1898
rect -894 1501 -888 1898
rect -938 1489 -888 1501
rect -772 1898 -722 1910
rect -772 1501 -766 1898
rect -728 1501 -722 1898
rect -772 1489 -722 1501
rect -606 1898 -556 1910
rect -606 1501 -600 1898
rect -562 1501 -556 1898
rect -606 1489 -556 1501
rect -440 1898 -390 1910
rect -440 1501 -434 1898
rect -396 1501 -390 1898
rect -440 1489 -390 1501
rect -274 1898 -224 1910
rect -274 1501 -268 1898
rect -230 1501 -224 1898
rect -274 1489 -224 1501
rect -108 1898 -58 1910
rect -108 1501 -102 1898
rect -64 1501 -58 1898
rect -108 1489 -58 1501
rect 58 1898 108 1910
rect 58 1501 64 1898
rect 102 1501 108 1898
rect 58 1489 108 1501
rect 224 1898 274 1910
rect 224 1501 230 1898
rect 268 1501 274 1898
rect 224 1489 274 1501
rect 390 1898 440 1910
rect 390 1501 396 1898
rect 434 1501 440 1898
rect 390 1489 440 1501
rect 556 1898 606 1910
rect 556 1501 562 1898
rect 600 1501 606 1898
rect 556 1489 606 1501
rect 722 1898 772 1910
rect 722 1501 728 1898
rect 766 1501 772 1898
rect 722 1489 772 1501
rect 888 1898 938 1910
rect 888 1501 894 1898
rect 932 1501 938 1898
rect 888 1489 938 1501
rect 1054 1898 1104 1910
rect 1054 1501 1060 1898
rect 1098 1501 1104 1898
rect 1054 1489 1104 1501
rect 1220 1898 1270 1910
rect 1220 1501 1226 1898
rect 1264 1501 1270 1898
rect 1220 1489 1270 1501
rect 1386 1898 1436 1910
rect 1386 1501 1392 1898
rect 1430 1501 1436 1898
rect 1386 1489 1436 1501
rect 1552 1898 1602 1910
rect 1552 1501 1558 1898
rect 1596 1501 1602 1898
rect 1552 1489 1602 1501
rect 1718 1898 1768 1910
rect 1718 1501 1724 1898
rect 1762 1501 1768 1898
rect 1718 1489 1768 1501
rect 1884 1898 1934 1910
rect 1884 1501 1890 1898
rect 1928 1501 1934 1898
rect 1884 1489 1934 1501
rect 2050 1898 2100 1910
rect 2050 1501 2056 1898
rect 2094 1501 2100 1898
rect 2050 1489 2100 1501
rect 2216 1898 2266 1910
rect 2216 1501 2222 1898
rect 2260 1501 2266 1898
rect 2216 1489 2266 1501
rect 2382 1898 2432 1910
rect 2382 1501 2388 1898
rect 2426 1501 2432 1898
rect 2382 1489 2432 1501
rect 2548 1898 2598 1910
rect 2548 1501 2554 1898
rect 2592 1501 2598 1898
rect 2548 1489 2598 1501
rect 2714 1898 2764 1910
rect 2714 1501 2720 1898
rect 2758 1501 2764 1898
rect 2714 1489 2764 1501
rect 2880 1898 2930 1910
rect 2880 1501 2886 1898
rect 2924 1501 2930 1898
rect 2880 1489 2930 1501
rect 3046 1898 3096 1910
rect 3046 1501 3052 1898
rect 3090 1501 3096 1898
rect 3046 1489 3096 1501
rect 3212 1898 3262 1910
rect 3212 1501 3218 1898
rect 3256 1501 3262 1898
rect 3212 1489 3262 1501
rect 3378 1898 3428 1910
rect 3378 1501 3384 1898
rect 3422 1501 3428 1898
rect 3378 1489 3428 1501
rect 3544 1898 3594 1910
rect 3544 1501 3550 1898
rect 3588 1501 3594 1898
rect 3544 1489 3594 1501
rect 3710 1898 3760 1910
rect 3710 1501 3716 1898
rect 3754 1501 3760 1898
rect 3710 1489 3760 1501
rect 3876 1898 3926 1910
rect 3876 1501 3882 1898
rect 3920 1501 3926 1898
rect 3876 1489 3926 1501
rect 4042 1898 4092 1910
rect 4042 1501 4048 1898
rect 4086 1501 4092 1898
rect 4042 1489 4092 1501
rect 4208 1898 4258 1910
rect 4208 1501 4214 1898
rect 4252 1501 4258 1898
rect 4208 1489 4258 1501
rect 4374 1898 4424 1910
rect 4374 1501 4380 1898
rect 4418 1501 4424 1898
rect 4374 1489 4424 1501
rect 4540 1898 4590 1910
rect 4540 1501 4546 1898
rect 4584 1501 4590 1898
rect 4540 1489 4590 1501
rect 4706 1898 4756 1910
rect 4706 1501 4712 1898
rect 4750 1501 4756 1898
rect 4706 1489 4756 1501
rect 4872 1898 4922 1910
rect 4872 1501 4878 1898
rect 4916 1501 4922 1898
rect 4872 1489 4922 1501
rect 5038 1898 5088 1910
rect 5038 1501 5044 1898
rect 5082 1501 5088 1898
rect 5038 1489 5088 1501
rect 5204 1898 5254 1910
rect 5204 1501 5210 1898
rect 5248 1501 5254 1898
rect 5204 1489 5254 1501
rect 5370 1898 5420 1910
rect 5370 1501 5376 1898
rect 5414 1501 5420 1898
rect 5370 1489 5420 1501
rect 5536 1898 5586 1910
rect 5536 1501 5542 1898
rect 5580 1501 5586 1898
rect 5536 1489 5586 1501
rect 5702 1898 5752 1910
rect 5702 1501 5708 1898
rect 5746 1501 5752 1898
rect 5702 1489 5752 1501
rect 5868 1898 5918 1910
rect 5868 1501 5874 1898
rect 5912 1501 5918 1898
rect 5868 1489 5918 1501
rect 6034 1898 6084 1910
rect 6034 1501 6040 1898
rect 6078 1501 6084 1898
rect 6034 1489 6084 1501
rect 6200 1898 6250 1910
rect 6200 1501 6206 1898
rect 6244 1501 6250 1898
rect 6200 1489 6250 1501
rect 6366 1898 6416 1910
rect 6366 1501 6372 1898
rect 6410 1501 6416 1898
rect 6366 1489 6416 1501
rect 6532 1898 6582 1910
rect 6532 1501 6538 1898
rect 6576 1501 6582 1898
rect 6532 1489 6582 1501
rect 6698 1898 6748 1910
rect 6698 1501 6704 1898
rect 6742 1501 6748 1898
rect 6698 1489 6748 1501
rect 6864 1898 6914 1910
rect 6864 1501 6870 1898
rect 6908 1501 6914 1898
rect 6864 1489 6914 1501
rect 7030 1898 7080 1910
rect 7030 1501 7036 1898
rect 7074 1501 7080 1898
rect 7030 1489 7080 1501
rect 7196 1898 7246 1910
rect 7196 1501 7202 1898
rect 7240 1501 7246 1898
rect 7196 1489 7246 1501
rect 7362 1898 7412 1910
rect 7362 1501 7368 1898
rect 7406 1501 7412 1898
rect 7362 1489 7412 1501
rect 7528 1898 7578 1910
rect 7528 1501 7534 1898
rect 7572 1501 7578 1898
rect 7528 1489 7578 1501
rect 7694 1898 7744 1910
rect 7694 1501 7700 1898
rect 7738 1501 7744 1898
rect 7694 1489 7744 1501
rect 7860 1898 7910 1910
rect 7860 1501 7866 1898
rect 7904 1501 7910 1898
rect 7860 1489 7910 1501
rect 8026 1898 8076 1910
rect 8026 1501 8032 1898
rect 8070 1501 8076 1898
rect 8026 1489 8076 1501
rect 8192 1898 8242 1910
rect 8192 1501 8198 1898
rect 8236 1501 8242 1898
rect 8192 1489 8242 1501
rect 8358 1898 8408 1910
rect 8358 1501 8364 1898
rect 8402 1501 8408 1898
rect 8358 1489 8408 1501
rect 8524 1898 8574 1910
rect 8524 1501 8530 1898
rect 8568 1501 8574 1898
rect 8524 1489 8574 1501
rect 8690 1898 8740 1910
rect 8690 1501 8696 1898
rect 8734 1501 8740 1898
rect 8690 1489 8740 1501
rect 8856 1898 8906 1910
rect 8856 1501 8862 1898
rect 8900 1501 8906 1898
rect 8856 1489 8906 1501
rect 9022 1898 9072 1910
rect 9022 1501 9028 1898
rect 9066 1501 9072 1898
rect 9022 1489 9072 1501
rect 9188 1898 9238 1910
rect 9188 1501 9194 1898
rect 9232 1501 9238 1898
rect 9188 1489 9238 1501
rect 9354 1898 9404 1910
rect 9354 1501 9360 1898
rect 9398 1501 9404 1898
rect 9354 1489 9404 1501
rect 9520 1898 9570 1910
rect 9520 1501 9526 1898
rect 9564 1501 9570 1898
rect 9520 1489 9570 1501
rect 9686 1898 9736 1910
rect 9686 1501 9692 1898
rect 9730 1501 9736 1898
rect 9686 1489 9736 1501
rect 9852 1898 9902 1910
rect 9852 1501 9858 1898
rect 9896 1501 9902 1898
rect 9852 1489 9902 1501
rect 10018 1898 10068 1910
rect 10018 1501 10024 1898
rect 10062 1501 10068 1898
rect 10018 1489 10068 1501
rect 10184 1898 10234 1910
rect 10184 1501 10190 1898
rect 10228 1501 10234 1898
rect 10184 1489 10234 1501
rect 10350 1898 10400 1910
rect 10350 1501 10356 1898
rect 10394 1501 10400 1898
rect 10350 1489 10400 1501
rect 10516 1898 10566 1910
rect 10516 1501 10522 1898
rect 10560 1501 10566 1898
rect 10516 1489 10566 1501
rect 10682 1898 10732 1910
rect 10682 1501 10688 1898
rect 10726 1501 10732 1898
rect 10682 1489 10732 1501
rect 10848 1898 10898 1910
rect 10848 1501 10854 1898
rect 10892 1501 10898 1898
rect 10848 1489 10898 1501
rect 11014 1898 11064 1910
rect 11014 1501 11020 1898
rect 11058 1501 11064 1898
rect 11014 1489 11064 1501
rect 11180 1898 11230 1910
rect 11180 1501 11186 1898
rect 11224 1501 11230 1898
rect 11180 1489 11230 1501
rect 11346 1898 11396 1910
rect 11346 1501 11352 1898
rect 11390 1501 11396 1898
rect 11346 1489 11396 1501
rect 11512 1898 11562 1910
rect 11512 1501 11518 1898
rect 11556 1501 11562 1898
rect 11512 1489 11562 1501
rect 11678 1898 11728 1910
rect 11678 1501 11684 1898
rect 11722 1501 11728 1898
rect 11678 1489 11728 1501
rect 11844 1898 11894 1910
rect 11844 1501 11850 1898
rect 11888 1501 11894 1898
rect 11844 1489 11894 1501
rect 12010 1898 12060 1910
rect 12010 1501 12016 1898
rect 12054 1501 12060 1898
rect 12010 1489 12060 1501
rect 12176 1898 12226 1910
rect 12176 1501 12182 1898
rect 12220 1501 12226 1898
rect 12176 1489 12226 1501
rect 12342 1898 12392 1910
rect 12342 1501 12348 1898
rect 12386 1501 12392 1898
rect 12342 1489 12392 1501
rect 12508 1898 12558 1910
rect 12508 1501 12514 1898
rect 12552 1501 12558 1898
rect 12508 1489 12558 1501
rect 12674 1898 12724 1910
rect 12674 1501 12680 1898
rect 12718 1501 12724 1898
rect 12674 1489 12724 1501
rect 12840 1898 12890 1910
rect 12840 1501 12846 1898
rect 12884 1501 12890 1898
rect 12840 1489 12890 1501
rect 13006 1898 13056 1910
rect 13006 1501 13012 1898
rect 13050 1501 13056 1898
rect 13006 1489 13056 1501
rect 13172 1898 13222 1910
rect 13172 1501 13178 1898
rect 13216 1501 13222 1898
rect 13172 1489 13222 1501
rect 13338 1898 13388 1910
rect 13338 1501 13344 1898
rect 13382 1501 13388 1898
rect 13338 1489 13388 1501
rect 13504 1898 13554 1910
rect 13504 1501 13510 1898
rect 13548 1501 13554 1898
rect 13504 1489 13554 1501
rect 13670 1898 13720 1910
rect 13670 1501 13676 1898
rect 13714 1501 13720 1898
rect 13670 1489 13720 1501
rect 13836 1898 13886 1910
rect 13836 1501 13842 1898
rect 13880 1501 13886 1898
rect 13836 1489 13886 1501
rect -13886 -1501 -13836 -1489
rect -13886 -1898 -13880 -1501
rect -13842 -1898 -13836 -1501
rect -13886 -1910 -13836 -1898
rect -13720 -1501 -13670 -1489
rect -13720 -1898 -13714 -1501
rect -13676 -1898 -13670 -1501
rect -13720 -1910 -13670 -1898
rect -13554 -1501 -13504 -1489
rect -13554 -1898 -13548 -1501
rect -13510 -1898 -13504 -1501
rect -13554 -1910 -13504 -1898
rect -13388 -1501 -13338 -1489
rect -13388 -1898 -13382 -1501
rect -13344 -1898 -13338 -1501
rect -13388 -1910 -13338 -1898
rect -13222 -1501 -13172 -1489
rect -13222 -1898 -13216 -1501
rect -13178 -1898 -13172 -1501
rect -13222 -1910 -13172 -1898
rect -13056 -1501 -13006 -1489
rect -13056 -1898 -13050 -1501
rect -13012 -1898 -13006 -1501
rect -13056 -1910 -13006 -1898
rect -12890 -1501 -12840 -1489
rect -12890 -1898 -12884 -1501
rect -12846 -1898 -12840 -1501
rect -12890 -1910 -12840 -1898
rect -12724 -1501 -12674 -1489
rect -12724 -1898 -12718 -1501
rect -12680 -1898 -12674 -1501
rect -12724 -1910 -12674 -1898
rect -12558 -1501 -12508 -1489
rect -12558 -1898 -12552 -1501
rect -12514 -1898 -12508 -1501
rect -12558 -1910 -12508 -1898
rect -12392 -1501 -12342 -1489
rect -12392 -1898 -12386 -1501
rect -12348 -1898 -12342 -1501
rect -12392 -1910 -12342 -1898
rect -12226 -1501 -12176 -1489
rect -12226 -1898 -12220 -1501
rect -12182 -1898 -12176 -1501
rect -12226 -1910 -12176 -1898
rect -12060 -1501 -12010 -1489
rect -12060 -1898 -12054 -1501
rect -12016 -1898 -12010 -1501
rect -12060 -1910 -12010 -1898
rect -11894 -1501 -11844 -1489
rect -11894 -1898 -11888 -1501
rect -11850 -1898 -11844 -1501
rect -11894 -1910 -11844 -1898
rect -11728 -1501 -11678 -1489
rect -11728 -1898 -11722 -1501
rect -11684 -1898 -11678 -1501
rect -11728 -1910 -11678 -1898
rect -11562 -1501 -11512 -1489
rect -11562 -1898 -11556 -1501
rect -11518 -1898 -11512 -1501
rect -11562 -1910 -11512 -1898
rect -11396 -1501 -11346 -1489
rect -11396 -1898 -11390 -1501
rect -11352 -1898 -11346 -1501
rect -11396 -1910 -11346 -1898
rect -11230 -1501 -11180 -1489
rect -11230 -1898 -11224 -1501
rect -11186 -1898 -11180 -1501
rect -11230 -1910 -11180 -1898
rect -11064 -1501 -11014 -1489
rect -11064 -1898 -11058 -1501
rect -11020 -1898 -11014 -1501
rect -11064 -1910 -11014 -1898
rect -10898 -1501 -10848 -1489
rect -10898 -1898 -10892 -1501
rect -10854 -1898 -10848 -1501
rect -10898 -1910 -10848 -1898
rect -10732 -1501 -10682 -1489
rect -10732 -1898 -10726 -1501
rect -10688 -1898 -10682 -1501
rect -10732 -1910 -10682 -1898
rect -10566 -1501 -10516 -1489
rect -10566 -1898 -10560 -1501
rect -10522 -1898 -10516 -1501
rect -10566 -1910 -10516 -1898
rect -10400 -1501 -10350 -1489
rect -10400 -1898 -10394 -1501
rect -10356 -1898 -10350 -1501
rect -10400 -1910 -10350 -1898
rect -10234 -1501 -10184 -1489
rect -10234 -1898 -10228 -1501
rect -10190 -1898 -10184 -1501
rect -10234 -1910 -10184 -1898
rect -10068 -1501 -10018 -1489
rect -10068 -1898 -10062 -1501
rect -10024 -1898 -10018 -1501
rect -10068 -1910 -10018 -1898
rect -9902 -1501 -9852 -1489
rect -9902 -1898 -9896 -1501
rect -9858 -1898 -9852 -1501
rect -9902 -1910 -9852 -1898
rect -9736 -1501 -9686 -1489
rect -9736 -1898 -9730 -1501
rect -9692 -1898 -9686 -1501
rect -9736 -1910 -9686 -1898
rect -9570 -1501 -9520 -1489
rect -9570 -1898 -9564 -1501
rect -9526 -1898 -9520 -1501
rect -9570 -1910 -9520 -1898
rect -9404 -1501 -9354 -1489
rect -9404 -1898 -9398 -1501
rect -9360 -1898 -9354 -1501
rect -9404 -1910 -9354 -1898
rect -9238 -1501 -9188 -1489
rect -9238 -1898 -9232 -1501
rect -9194 -1898 -9188 -1501
rect -9238 -1910 -9188 -1898
rect -9072 -1501 -9022 -1489
rect -9072 -1898 -9066 -1501
rect -9028 -1898 -9022 -1501
rect -9072 -1910 -9022 -1898
rect -8906 -1501 -8856 -1489
rect -8906 -1898 -8900 -1501
rect -8862 -1898 -8856 -1501
rect -8906 -1910 -8856 -1898
rect -8740 -1501 -8690 -1489
rect -8740 -1898 -8734 -1501
rect -8696 -1898 -8690 -1501
rect -8740 -1910 -8690 -1898
rect -8574 -1501 -8524 -1489
rect -8574 -1898 -8568 -1501
rect -8530 -1898 -8524 -1501
rect -8574 -1910 -8524 -1898
rect -8408 -1501 -8358 -1489
rect -8408 -1898 -8402 -1501
rect -8364 -1898 -8358 -1501
rect -8408 -1910 -8358 -1898
rect -8242 -1501 -8192 -1489
rect -8242 -1898 -8236 -1501
rect -8198 -1898 -8192 -1501
rect -8242 -1910 -8192 -1898
rect -8076 -1501 -8026 -1489
rect -8076 -1898 -8070 -1501
rect -8032 -1898 -8026 -1501
rect -8076 -1910 -8026 -1898
rect -7910 -1501 -7860 -1489
rect -7910 -1898 -7904 -1501
rect -7866 -1898 -7860 -1501
rect -7910 -1910 -7860 -1898
rect -7744 -1501 -7694 -1489
rect -7744 -1898 -7738 -1501
rect -7700 -1898 -7694 -1501
rect -7744 -1910 -7694 -1898
rect -7578 -1501 -7528 -1489
rect -7578 -1898 -7572 -1501
rect -7534 -1898 -7528 -1501
rect -7578 -1910 -7528 -1898
rect -7412 -1501 -7362 -1489
rect -7412 -1898 -7406 -1501
rect -7368 -1898 -7362 -1501
rect -7412 -1910 -7362 -1898
rect -7246 -1501 -7196 -1489
rect -7246 -1898 -7240 -1501
rect -7202 -1898 -7196 -1501
rect -7246 -1910 -7196 -1898
rect -7080 -1501 -7030 -1489
rect -7080 -1898 -7074 -1501
rect -7036 -1898 -7030 -1501
rect -7080 -1910 -7030 -1898
rect -6914 -1501 -6864 -1489
rect -6914 -1898 -6908 -1501
rect -6870 -1898 -6864 -1501
rect -6914 -1910 -6864 -1898
rect -6748 -1501 -6698 -1489
rect -6748 -1898 -6742 -1501
rect -6704 -1898 -6698 -1501
rect -6748 -1910 -6698 -1898
rect -6582 -1501 -6532 -1489
rect -6582 -1898 -6576 -1501
rect -6538 -1898 -6532 -1501
rect -6582 -1910 -6532 -1898
rect -6416 -1501 -6366 -1489
rect -6416 -1898 -6410 -1501
rect -6372 -1898 -6366 -1501
rect -6416 -1910 -6366 -1898
rect -6250 -1501 -6200 -1489
rect -6250 -1898 -6244 -1501
rect -6206 -1898 -6200 -1501
rect -6250 -1910 -6200 -1898
rect -6084 -1501 -6034 -1489
rect -6084 -1898 -6078 -1501
rect -6040 -1898 -6034 -1501
rect -6084 -1910 -6034 -1898
rect -5918 -1501 -5868 -1489
rect -5918 -1898 -5912 -1501
rect -5874 -1898 -5868 -1501
rect -5918 -1910 -5868 -1898
rect -5752 -1501 -5702 -1489
rect -5752 -1898 -5746 -1501
rect -5708 -1898 -5702 -1501
rect -5752 -1910 -5702 -1898
rect -5586 -1501 -5536 -1489
rect -5586 -1898 -5580 -1501
rect -5542 -1898 -5536 -1501
rect -5586 -1910 -5536 -1898
rect -5420 -1501 -5370 -1489
rect -5420 -1898 -5414 -1501
rect -5376 -1898 -5370 -1501
rect -5420 -1910 -5370 -1898
rect -5254 -1501 -5204 -1489
rect -5254 -1898 -5248 -1501
rect -5210 -1898 -5204 -1501
rect -5254 -1910 -5204 -1898
rect -5088 -1501 -5038 -1489
rect -5088 -1898 -5082 -1501
rect -5044 -1898 -5038 -1501
rect -5088 -1910 -5038 -1898
rect -4922 -1501 -4872 -1489
rect -4922 -1898 -4916 -1501
rect -4878 -1898 -4872 -1501
rect -4922 -1910 -4872 -1898
rect -4756 -1501 -4706 -1489
rect -4756 -1898 -4750 -1501
rect -4712 -1898 -4706 -1501
rect -4756 -1910 -4706 -1898
rect -4590 -1501 -4540 -1489
rect -4590 -1898 -4584 -1501
rect -4546 -1898 -4540 -1501
rect -4590 -1910 -4540 -1898
rect -4424 -1501 -4374 -1489
rect -4424 -1898 -4418 -1501
rect -4380 -1898 -4374 -1501
rect -4424 -1910 -4374 -1898
rect -4258 -1501 -4208 -1489
rect -4258 -1898 -4252 -1501
rect -4214 -1898 -4208 -1501
rect -4258 -1910 -4208 -1898
rect -4092 -1501 -4042 -1489
rect -4092 -1898 -4086 -1501
rect -4048 -1898 -4042 -1501
rect -4092 -1910 -4042 -1898
rect -3926 -1501 -3876 -1489
rect -3926 -1898 -3920 -1501
rect -3882 -1898 -3876 -1501
rect -3926 -1910 -3876 -1898
rect -3760 -1501 -3710 -1489
rect -3760 -1898 -3754 -1501
rect -3716 -1898 -3710 -1501
rect -3760 -1910 -3710 -1898
rect -3594 -1501 -3544 -1489
rect -3594 -1898 -3588 -1501
rect -3550 -1898 -3544 -1501
rect -3594 -1910 -3544 -1898
rect -3428 -1501 -3378 -1489
rect -3428 -1898 -3422 -1501
rect -3384 -1898 -3378 -1501
rect -3428 -1910 -3378 -1898
rect -3262 -1501 -3212 -1489
rect -3262 -1898 -3256 -1501
rect -3218 -1898 -3212 -1501
rect -3262 -1910 -3212 -1898
rect -3096 -1501 -3046 -1489
rect -3096 -1898 -3090 -1501
rect -3052 -1898 -3046 -1501
rect -3096 -1910 -3046 -1898
rect -2930 -1501 -2880 -1489
rect -2930 -1898 -2924 -1501
rect -2886 -1898 -2880 -1501
rect -2930 -1910 -2880 -1898
rect -2764 -1501 -2714 -1489
rect -2764 -1898 -2758 -1501
rect -2720 -1898 -2714 -1501
rect -2764 -1910 -2714 -1898
rect -2598 -1501 -2548 -1489
rect -2598 -1898 -2592 -1501
rect -2554 -1898 -2548 -1501
rect -2598 -1910 -2548 -1898
rect -2432 -1501 -2382 -1489
rect -2432 -1898 -2426 -1501
rect -2388 -1898 -2382 -1501
rect -2432 -1910 -2382 -1898
rect -2266 -1501 -2216 -1489
rect -2266 -1898 -2260 -1501
rect -2222 -1898 -2216 -1501
rect -2266 -1910 -2216 -1898
rect -2100 -1501 -2050 -1489
rect -2100 -1898 -2094 -1501
rect -2056 -1898 -2050 -1501
rect -2100 -1910 -2050 -1898
rect -1934 -1501 -1884 -1489
rect -1934 -1898 -1928 -1501
rect -1890 -1898 -1884 -1501
rect -1934 -1910 -1884 -1898
rect -1768 -1501 -1718 -1489
rect -1768 -1898 -1762 -1501
rect -1724 -1898 -1718 -1501
rect -1768 -1910 -1718 -1898
rect -1602 -1501 -1552 -1489
rect -1602 -1898 -1596 -1501
rect -1558 -1898 -1552 -1501
rect -1602 -1910 -1552 -1898
rect -1436 -1501 -1386 -1489
rect -1436 -1898 -1430 -1501
rect -1392 -1898 -1386 -1501
rect -1436 -1910 -1386 -1898
rect -1270 -1501 -1220 -1489
rect -1270 -1898 -1264 -1501
rect -1226 -1898 -1220 -1501
rect -1270 -1910 -1220 -1898
rect -1104 -1501 -1054 -1489
rect -1104 -1898 -1098 -1501
rect -1060 -1898 -1054 -1501
rect -1104 -1910 -1054 -1898
rect -938 -1501 -888 -1489
rect -938 -1898 -932 -1501
rect -894 -1898 -888 -1501
rect -938 -1910 -888 -1898
rect -772 -1501 -722 -1489
rect -772 -1898 -766 -1501
rect -728 -1898 -722 -1501
rect -772 -1910 -722 -1898
rect -606 -1501 -556 -1489
rect -606 -1898 -600 -1501
rect -562 -1898 -556 -1501
rect -606 -1910 -556 -1898
rect -440 -1501 -390 -1489
rect -440 -1898 -434 -1501
rect -396 -1898 -390 -1501
rect -440 -1910 -390 -1898
rect -274 -1501 -224 -1489
rect -274 -1898 -268 -1501
rect -230 -1898 -224 -1501
rect -274 -1910 -224 -1898
rect -108 -1501 -58 -1489
rect -108 -1898 -102 -1501
rect -64 -1898 -58 -1501
rect -108 -1910 -58 -1898
rect 58 -1501 108 -1489
rect 58 -1898 64 -1501
rect 102 -1898 108 -1501
rect 58 -1910 108 -1898
rect 224 -1501 274 -1489
rect 224 -1898 230 -1501
rect 268 -1898 274 -1501
rect 224 -1910 274 -1898
rect 390 -1501 440 -1489
rect 390 -1898 396 -1501
rect 434 -1898 440 -1501
rect 390 -1910 440 -1898
rect 556 -1501 606 -1489
rect 556 -1898 562 -1501
rect 600 -1898 606 -1501
rect 556 -1910 606 -1898
rect 722 -1501 772 -1489
rect 722 -1898 728 -1501
rect 766 -1898 772 -1501
rect 722 -1910 772 -1898
rect 888 -1501 938 -1489
rect 888 -1898 894 -1501
rect 932 -1898 938 -1501
rect 888 -1910 938 -1898
rect 1054 -1501 1104 -1489
rect 1054 -1898 1060 -1501
rect 1098 -1898 1104 -1501
rect 1054 -1910 1104 -1898
rect 1220 -1501 1270 -1489
rect 1220 -1898 1226 -1501
rect 1264 -1898 1270 -1501
rect 1220 -1910 1270 -1898
rect 1386 -1501 1436 -1489
rect 1386 -1898 1392 -1501
rect 1430 -1898 1436 -1501
rect 1386 -1910 1436 -1898
rect 1552 -1501 1602 -1489
rect 1552 -1898 1558 -1501
rect 1596 -1898 1602 -1501
rect 1552 -1910 1602 -1898
rect 1718 -1501 1768 -1489
rect 1718 -1898 1724 -1501
rect 1762 -1898 1768 -1501
rect 1718 -1910 1768 -1898
rect 1884 -1501 1934 -1489
rect 1884 -1898 1890 -1501
rect 1928 -1898 1934 -1501
rect 1884 -1910 1934 -1898
rect 2050 -1501 2100 -1489
rect 2050 -1898 2056 -1501
rect 2094 -1898 2100 -1501
rect 2050 -1910 2100 -1898
rect 2216 -1501 2266 -1489
rect 2216 -1898 2222 -1501
rect 2260 -1898 2266 -1501
rect 2216 -1910 2266 -1898
rect 2382 -1501 2432 -1489
rect 2382 -1898 2388 -1501
rect 2426 -1898 2432 -1501
rect 2382 -1910 2432 -1898
rect 2548 -1501 2598 -1489
rect 2548 -1898 2554 -1501
rect 2592 -1898 2598 -1501
rect 2548 -1910 2598 -1898
rect 2714 -1501 2764 -1489
rect 2714 -1898 2720 -1501
rect 2758 -1898 2764 -1501
rect 2714 -1910 2764 -1898
rect 2880 -1501 2930 -1489
rect 2880 -1898 2886 -1501
rect 2924 -1898 2930 -1501
rect 2880 -1910 2930 -1898
rect 3046 -1501 3096 -1489
rect 3046 -1898 3052 -1501
rect 3090 -1898 3096 -1501
rect 3046 -1910 3096 -1898
rect 3212 -1501 3262 -1489
rect 3212 -1898 3218 -1501
rect 3256 -1898 3262 -1501
rect 3212 -1910 3262 -1898
rect 3378 -1501 3428 -1489
rect 3378 -1898 3384 -1501
rect 3422 -1898 3428 -1501
rect 3378 -1910 3428 -1898
rect 3544 -1501 3594 -1489
rect 3544 -1898 3550 -1501
rect 3588 -1898 3594 -1501
rect 3544 -1910 3594 -1898
rect 3710 -1501 3760 -1489
rect 3710 -1898 3716 -1501
rect 3754 -1898 3760 -1501
rect 3710 -1910 3760 -1898
rect 3876 -1501 3926 -1489
rect 3876 -1898 3882 -1501
rect 3920 -1898 3926 -1501
rect 3876 -1910 3926 -1898
rect 4042 -1501 4092 -1489
rect 4042 -1898 4048 -1501
rect 4086 -1898 4092 -1501
rect 4042 -1910 4092 -1898
rect 4208 -1501 4258 -1489
rect 4208 -1898 4214 -1501
rect 4252 -1898 4258 -1501
rect 4208 -1910 4258 -1898
rect 4374 -1501 4424 -1489
rect 4374 -1898 4380 -1501
rect 4418 -1898 4424 -1501
rect 4374 -1910 4424 -1898
rect 4540 -1501 4590 -1489
rect 4540 -1898 4546 -1501
rect 4584 -1898 4590 -1501
rect 4540 -1910 4590 -1898
rect 4706 -1501 4756 -1489
rect 4706 -1898 4712 -1501
rect 4750 -1898 4756 -1501
rect 4706 -1910 4756 -1898
rect 4872 -1501 4922 -1489
rect 4872 -1898 4878 -1501
rect 4916 -1898 4922 -1501
rect 4872 -1910 4922 -1898
rect 5038 -1501 5088 -1489
rect 5038 -1898 5044 -1501
rect 5082 -1898 5088 -1501
rect 5038 -1910 5088 -1898
rect 5204 -1501 5254 -1489
rect 5204 -1898 5210 -1501
rect 5248 -1898 5254 -1501
rect 5204 -1910 5254 -1898
rect 5370 -1501 5420 -1489
rect 5370 -1898 5376 -1501
rect 5414 -1898 5420 -1501
rect 5370 -1910 5420 -1898
rect 5536 -1501 5586 -1489
rect 5536 -1898 5542 -1501
rect 5580 -1898 5586 -1501
rect 5536 -1910 5586 -1898
rect 5702 -1501 5752 -1489
rect 5702 -1898 5708 -1501
rect 5746 -1898 5752 -1501
rect 5702 -1910 5752 -1898
rect 5868 -1501 5918 -1489
rect 5868 -1898 5874 -1501
rect 5912 -1898 5918 -1501
rect 5868 -1910 5918 -1898
rect 6034 -1501 6084 -1489
rect 6034 -1898 6040 -1501
rect 6078 -1898 6084 -1501
rect 6034 -1910 6084 -1898
rect 6200 -1501 6250 -1489
rect 6200 -1898 6206 -1501
rect 6244 -1898 6250 -1501
rect 6200 -1910 6250 -1898
rect 6366 -1501 6416 -1489
rect 6366 -1898 6372 -1501
rect 6410 -1898 6416 -1501
rect 6366 -1910 6416 -1898
rect 6532 -1501 6582 -1489
rect 6532 -1898 6538 -1501
rect 6576 -1898 6582 -1501
rect 6532 -1910 6582 -1898
rect 6698 -1501 6748 -1489
rect 6698 -1898 6704 -1501
rect 6742 -1898 6748 -1501
rect 6698 -1910 6748 -1898
rect 6864 -1501 6914 -1489
rect 6864 -1898 6870 -1501
rect 6908 -1898 6914 -1501
rect 6864 -1910 6914 -1898
rect 7030 -1501 7080 -1489
rect 7030 -1898 7036 -1501
rect 7074 -1898 7080 -1501
rect 7030 -1910 7080 -1898
rect 7196 -1501 7246 -1489
rect 7196 -1898 7202 -1501
rect 7240 -1898 7246 -1501
rect 7196 -1910 7246 -1898
rect 7362 -1501 7412 -1489
rect 7362 -1898 7368 -1501
rect 7406 -1898 7412 -1501
rect 7362 -1910 7412 -1898
rect 7528 -1501 7578 -1489
rect 7528 -1898 7534 -1501
rect 7572 -1898 7578 -1501
rect 7528 -1910 7578 -1898
rect 7694 -1501 7744 -1489
rect 7694 -1898 7700 -1501
rect 7738 -1898 7744 -1501
rect 7694 -1910 7744 -1898
rect 7860 -1501 7910 -1489
rect 7860 -1898 7866 -1501
rect 7904 -1898 7910 -1501
rect 7860 -1910 7910 -1898
rect 8026 -1501 8076 -1489
rect 8026 -1898 8032 -1501
rect 8070 -1898 8076 -1501
rect 8026 -1910 8076 -1898
rect 8192 -1501 8242 -1489
rect 8192 -1898 8198 -1501
rect 8236 -1898 8242 -1501
rect 8192 -1910 8242 -1898
rect 8358 -1501 8408 -1489
rect 8358 -1898 8364 -1501
rect 8402 -1898 8408 -1501
rect 8358 -1910 8408 -1898
rect 8524 -1501 8574 -1489
rect 8524 -1898 8530 -1501
rect 8568 -1898 8574 -1501
rect 8524 -1910 8574 -1898
rect 8690 -1501 8740 -1489
rect 8690 -1898 8696 -1501
rect 8734 -1898 8740 -1501
rect 8690 -1910 8740 -1898
rect 8856 -1501 8906 -1489
rect 8856 -1898 8862 -1501
rect 8900 -1898 8906 -1501
rect 8856 -1910 8906 -1898
rect 9022 -1501 9072 -1489
rect 9022 -1898 9028 -1501
rect 9066 -1898 9072 -1501
rect 9022 -1910 9072 -1898
rect 9188 -1501 9238 -1489
rect 9188 -1898 9194 -1501
rect 9232 -1898 9238 -1501
rect 9188 -1910 9238 -1898
rect 9354 -1501 9404 -1489
rect 9354 -1898 9360 -1501
rect 9398 -1898 9404 -1501
rect 9354 -1910 9404 -1898
rect 9520 -1501 9570 -1489
rect 9520 -1898 9526 -1501
rect 9564 -1898 9570 -1501
rect 9520 -1910 9570 -1898
rect 9686 -1501 9736 -1489
rect 9686 -1898 9692 -1501
rect 9730 -1898 9736 -1501
rect 9686 -1910 9736 -1898
rect 9852 -1501 9902 -1489
rect 9852 -1898 9858 -1501
rect 9896 -1898 9902 -1501
rect 9852 -1910 9902 -1898
rect 10018 -1501 10068 -1489
rect 10018 -1898 10024 -1501
rect 10062 -1898 10068 -1501
rect 10018 -1910 10068 -1898
rect 10184 -1501 10234 -1489
rect 10184 -1898 10190 -1501
rect 10228 -1898 10234 -1501
rect 10184 -1910 10234 -1898
rect 10350 -1501 10400 -1489
rect 10350 -1898 10356 -1501
rect 10394 -1898 10400 -1501
rect 10350 -1910 10400 -1898
rect 10516 -1501 10566 -1489
rect 10516 -1898 10522 -1501
rect 10560 -1898 10566 -1501
rect 10516 -1910 10566 -1898
rect 10682 -1501 10732 -1489
rect 10682 -1898 10688 -1501
rect 10726 -1898 10732 -1501
rect 10682 -1910 10732 -1898
rect 10848 -1501 10898 -1489
rect 10848 -1898 10854 -1501
rect 10892 -1898 10898 -1501
rect 10848 -1910 10898 -1898
rect 11014 -1501 11064 -1489
rect 11014 -1898 11020 -1501
rect 11058 -1898 11064 -1501
rect 11014 -1910 11064 -1898
rect 11180 -1501 11230 -1489
rect 11180 -1898 11186 -1501
rect 11224 -1898 11230 -1501
rect 11180 -1910 11230 -1898
rect 11346 -1501 11396 -1489
rect 11346 -1898 11352 -1501
rect 11390 -1898 11396 -1501
rect 11346 -1910 11396 -1898
rect 11512 -1501 11562 -1489
rect 11512 -1898 11518 -1501
rect 11556 -1898 11562 -1501
rect 11512 -1910 11562 -1898
rect 11678 -1501 11728 -1489
rect 11678 -1898 11684 -1501
rect 11722 -1898 11728 -1501
rect 11678 -1910 11728 -1898
rect 11844 -1501 11894 -1489
rect 11844 -1898 11850 -1501
rect 11888 -1898 11894 -1501
rect 11844 -1910 11894 -1898
rect 12010 -1501 12060 -1489
rect 12010 -1898 12016 -1501
rect 12054 -1898 12060 -1501
rect 12010 -1910 12060 -1898
rect 12176 -1501 12226 -1489
rect 12176 -1898 12182 -1501
rect 12220 -1898 12226 -1501
rect 12176 -1910 12226 -1898
rect 12342 -1501 12392 -1489
rect 12342 -1898 12348 -1501
rect 12386 -1898 12392 -1501
rect 12342 -1910 12392 -1898
rect 12508 -1501 12558 -1489
rect 12508 -1898 12514 -1501
rect 12552 -1898 12558 -1501
rect 12508 -1910 12558 -1898
rect 12674 -1501 12724 -1489
rect 12674 -1898 12680 -1501
rect 12718 -1898 12724 -1501
rect 12674 -1910 12724 -1898
rect 12840 -1501 12890 -1489
rect 12840 -1898 12846 -1501
rect 12884 -1898 12890 -1501
rect 12840 -1910 12890 -1898
rect 13006 -1501 13056 -1489
rect 13006 -1898 13012 -1501
rect 13050 -1898 13056 -1501
rect 13006 -1910 13056 -1898
rect 13172 -1501 13222 -1489
rect 13172 -1898 13178 -1501
rect 13216 -1898 13222 -1501
rect 13172 -1910 13222 -1898
rect 13338 -1501 13388 -1489
rect 13338 -1898 13344 -1501
rect 13382 -1898 13388 -1501
rect 13338 -1910 13388 -1898
rect 13504 -1501 13554 -1489
rect 13504 -1898 13510 -1501
rect 13548 -1898 13554 -1501
rect 13504 -1910 13554 -1898
rect 13670 -1501 13720 -1489
rect 13670 -1898 13676 -1501
rect 13714 -1898 13720 -1501
rect 13670 -1910 13720 -1898
rect 13836 -1501 13886 -1489
rect 13836 -1898 13842 -1501
rect 13880 -1898 13886 -1501
rect 13836 -1910 13886 -1898
<< properties >>
string FIXED_BBOX -14009 -2029 14009 2029
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 15.0 m 1 nx 168 wmin 0.350 lmin 0.50 class resistor rho 2000 val 86.789k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
