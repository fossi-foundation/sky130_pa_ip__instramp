magic
tech sky130A
magscale 1 2
timestamp 1729620069
<< pwell >>
rect -11818 -10582 11818 10582
<< psubdiff >>
rect -11782 10512 -11686 10546
rect 11686 10512 11782 10546
rect -11782 10450 -11748 10512
rect 11748 10450 11782 10512
rect -11782 -10512 -11748 -10450
rect 11748 -10512 11782 -10450
rect -11782 -10546 -11686 -10512
rect 11686 -10546 11782 -10512
<< psubdiffcont >>
rect -11686 10512 11686 10546
rect -11782 -10450 -11748 10450
rect 11748 -10450 11782 10450
rect -11686 -10546 11686 -10512
<< xpolycontact >>
rect -11652 9984 -11514 10416
rect -11652 -10416 -11514 -9984
rect -11418 9984 -11280 10416
rect -11418 -10416 -11280 -9984
rect -11184 9984 -11046 10416
rect -11184 -10416 -11046 -9984
rect -10950 9984 -10812 10416
rect -10950 -10416 -10812 -9984
rect -10716 9984 -10578 10416
rect -10716 -10416 -10578 -9984
rect -10482 9984 -10344 10416
rect -10482 -10416 -10344 -9984
rect -10248 9984 -10110 10416
rect -10248 -10416 -10110 -9984
rect -10014 9984 -9876 10416
rect -10014 -10416 -9876 -9984
rect -9780 9984 -9642 10416
rect -9780 -10416 -9642 -9984
rect -9546 9984 -9408 10416
rect -9546 -10416 -9408 -9984
rect -9312 9984 -9174 10416
rect -9312 -10416 -9174 -9984
rect -9078 9984 -8940 10416
rect -9078 -10416 -8940 -9984
rect -8844 9984 -8706 10416
rect -8844 -10416 -8706 -9984
rect -8610 9984 -8472 10416
rect -8610 -10416 -8472 -9984
rect -8376 9984 -8238 10416
rect -8376 -10416 -8238 -9984
rect -8142 9984 -8004 10416
rect -8142 -10416 -8004 -9984
rect -7908 9984 -7770 10416
rect -7908 -10416 -7770 -9984
rect -7674 9984 -7536 10416
rect -7674 -10416 -7536 -9984
rect -7440 9984 -7302 10416
rect -7440 -10416 -7302 -9984
rect -7206 9984 -7068 10416
rect -7206 -10416 -7068 -9984
rect -6972 9984 -6834 10416
rect -6972 -10416 -6834 -9984
rect -6738 9984 -6600 10416
rect -6738 -10416 -6600 -9984
rect -6504 9984 -6366 10416
rect -6504 -10416 -6366 -9984
rect -6270 9984 -6132 10416
rect -6270 -10416 -6132 -9984
rect -6036 9984 -5898 10416
rect -6036 -10416 -5898 -9984
rect -5802 9984 -5664 10416
rect -5802 -10416 -5664 -9984
rect -5568 9984 -5430 10416
rect -5568 -10416 -5430 -9984
rect -5334 9984 -5196 10416
rect -5334 -10416 -5196 -9984
rect -5100 9984 -4962 10416
rect -5100 -10416 -4962 -9984
rect -4866 9984 -4728 10416
rect -4866 -10416 -4728 -9984
rect -4632 9984 -4494 10416
rect -4632 -10416 -4494 -9984
rect -4398 9984 -4260 10416
rect -4398 -10416 -4260 -9984
rect -4164 9984 -4026 10416
rect -4164 -10416 -4026 -9984
rect -3930 9984 -3792 10416
rect -3930 -10416 -3792 -9984
rect -3696 9984 -3558 10416
rect -3696 -10416 -3558 -9984
rect -3462 9984 -3324 10416
rect -3462 -10416 -3324 -9984
rect -3228 9984 -3090 10416
rect -3228 -10416 -3090 -9984
rect -2994 9984 -2856 10416
rect -2994 -10416 -2856 -9984
rect -2760 9984 -2622 10416
rect -2760 -10416 -2622 -9984
rect -2526 9984 -2388 10416
rect -2526 -10416 -2388 -9984
rect -2292 9984 -2154 10416
rect -2292 -10416 -2154 -9984
rect -2058 9984 -1920 10416
rect -2058 -10416 -1920 -9984
rect -1824 9984 -1686 10416
rect -1824 -10416 -1686 -9984
rect -1590 9984 -1452 10416
rect -1590 -10416 -1452 -9984
rect -1356 9984 -1218 10416
rect -1356 -10416 -1218 -9984
rect -1122 9984 -984 10416
rect -1122 -10416 -984 -9984
rect -888 9984 -750 10416
rect -888 -10416 -750 -9984
rect -654 9984 -516 10416
rect -654 -10416 -516 -9984
rect -420 9984 -282 10416
rect -420 -10416 -282 -9984
rect -186 9984 -48 10416
rect -186 -10416 -48 -9984
rect 48 9984 186 10416
rect 48 -10416 186 -9984
rect 282 9984 420 10416
rect 282 -10416 420 -9984
rect 516 9984 654 10416
rect 516 -10416 654 -9984
rect 750 9984 888 10416
rect 750 -10416 888 -9984
rect 984 9984 1122 10416
rect 984 -10416 1122 -9984
rect 1218 9984 1356 10416
rect 1218 -10416 1356 -9984
rect 1452 9984 1590 10416
rect 1452 -10416 1590 -9984
rect 1686 9984 1824 10416
rect 1686 -10416 1824 -9984
rect 1920 9984 2058 10416
rect 1920 -10416 2058 -9984
rect 2154 9984 2292 10416
rect 2154 -10416 2292 -9984
rect 2388 9984 2526 10416
rect 2388 -10416 2526 -9984
rect 2622 9984 2760 10416
rect 2622 -10416 2760 -9984
rect 2856 9984 2994 10416
rect 2856 -10416 2994 -9984
rect 3090 9984 3228 10416
rect 3090 -10416 3228 -9984
rect 3324 9984 3462 10416
rect 3324 -10416 3462 -9984
rect 3558 9984 3696 10416
rect 3558 -10416 3696 -9984
rect 3792 9984 3930 10416
rect 3792 -10416 3930 -9984
rect 4026 9984 4164 10416
rect 4026 -10416 4164 -9984
rect 4260 9984 4398 10416
rect 4260 -10416 4398 -9984
rect 4494 9984 4632 10416
rect 4494 -10416 4632 -9984
rect 4728 9984 4866 10416
rect 4728 -10416 4866 -9984
rect 4962 9984 5100 10416
rect 4962 -10416 5100 -9984
rect 5196 9984 5334 10416
rect 5196 -10416 5334 -9984
rect 5430 9984 5568 10416
rect 5430 -10416 5568 -9984
rect 5664 9984 5802 10416
rect 5664 -10416 5802 -9984
rect 5898 9984 6036 10416
rect 5898 -10416 6036 -9984
rect 6132 9984 6270 10416
rect 6132 -10416 6270 -9984
rect 6366 9984 6504 10416
rect 6366 -10416 6504 -9984
rect 6600 9984 6738 10416
rect 6600 -10416 6738 -9984
rect 6834 9984 6972 10416
rect 6834 -10416 6972 -9984
rect 7068 9984 7206 10416
rect 7068 -10416 7206 -9984
rect 7302 9984 7440 10416
rect 7302 -10416 7440 -9984
rect 7536 9984 7674 10416
rect 7536 -10416 7674 -9984
rect 7770 9984 7908 10416
rect 7770 -10416 7908 -9984
rect 8004 9984 8142 10416
rect 8004 -10416 8142 -9984
rect 8238 9984 8376 10416
rect 8238 -10416 8376 -9984
rect 8472 9984 8610 10416
rect 8472 -10416 8610 -9984
rect 8706 9984 8844 10416
rect 8706 -10416 8844 -9984
rect 8940 9984 9078 10416
rect 8940 -10416 9078 -9984
rect 9174 9984 9312 10416
rect 9174 -10416 9312 -9984
rect 9408 9984 9546 10416
rect 9408 -10416 9546 -9984
rect 9642 9984 9780 10416
rect 9642 -10416 9780 -9984
rect 9876 9984 10014 10416
rect 9876 -10416 10014 -9984
rect 10110 9984 10248 10416
rect 10110 -10416 10248 -9984
rect 10344 9984 10482 10416
rect 10344 -10416 10482 -9984
rect 10578 9984 10716 10416
rect 10578 -10416 10716 -9984
rect 10812 9984 10950 10416
rect 10812 -10416 10950 -9984
rect 11046 9984 11184 10416
rect 11046 -10416 11184 -9984
rect 11280 9984 11418 10416
rect 11280 -10416 11418 -9984
rect 11514 9984 11652 10416
rect 11514 -10416 11652 -9984
<< ppolyres >>
rect -11652 -9984 -11514 9984
rect -11418 -9984 -11280 9984
rect -11184 -9984 -11046 9984
rect -10950 -9984 -10812 9984
rect -10716 -9984 -10578 9984
rect -10482 -9984 -10344 9984
rect -10248 -9984 -10110 9984
rect -10014 -9984 -9876 9984
rect -9780 -9984 -9642 9984
rect -9546 -9984 -9408 9984
rect -9312 -9984 -9174 9984
rect -9078 -9984 -8940 9984
rect -8844 -9984 -8706 9984
rect -8610 -9984 -8472 9984
rect -8376 -9984 -8238 9984
rect -8142 -9984 -8004 9984
rect -7908 -9984 -7770 9984
rect -7674 -9984 -7536 9984
rect -7440 -9984 -7302 9984
rect -7206 -9984 -7068 9984
rect -6972 -9984 -6834 9984
rect -6738 -9984 -6600 9984
rect -6504 -9984 -6366 9984
rect -6270 -9984 -6132 9984
rect -6036 -9984 -5898 9984
rect -5802 -9984 -5664 9984
rect -5568 -9984 -5430 9984
rect -5334 -9984 -5196 9984
rect -5100 -9984 -4962 9984
rect -4866 -9984 -4728 9984
rect -4632 -9984 -4494 9984
rect -4398 -9984 -4260 9984
rect -4164 -9984 -4026 9984
rect -3930 -9984 -3792 9984
rect -3696 -9984 -3558 9984
rect -3462 -9984 -3324 9984
rect -3228 -9984 -3090 9984
rect -2994 -9984 -2856 9984
rect -2760 -9984 -2622 9984
rect -2526 -9984 -2388 9984
rect -2292 -9984 -2154 9984
rect -2058 -9984 -1920 9984
rect -1824 -9984 -1686 9984
rect -1590 -9984 -1452 9984
rect -1356 -9984 -1218 9984
rect -1122 -9984 -984 9984
rect -888 -9984 -750 9984
rect -654 -9984 -516 9984
rect -420 -9984 -282 9984
rect -186 -9984 -48 9984
rect 48 -9984 186 9984
rect 282 -9984 420 9984
rect 516 -9984 654 9984
rect 750 -9984 888 9984
rect 984 -9984 1122 9984
rect 1218 -9984 1356 9984
rect 1452 -9984 1590 9984
rect 1686 -9984 1824 9984
rect 1920 -9984 2058 9984
rect 2154 -9984 2292 9984
rect 2388 -9984 2526 9984
rect 2622 -9984 2760 9984
rect 2856 -9984 2994 9984
rect 3090 -9984 3228 9984
rect 3324 -9984 3462 9984
rect 3558 -9984 3696 9984
rect 3792 -9984 3930 9984
rect 4026 -9984 4164 9984
rect 4260 -9984 4398 9984
rect 4494 -9984 4632 9984
rect 4728 -9984 4866 9984
rect 4962 -9984 5100 9984
rect 5196 -9984 5334 9984
rect 5430 -9984 5568 9984
rect 5664 -9984 5802 9984
rect 5898 -9984 6036 9984
rect 6132 -9984 6270 9984
rect 6366 -9984 6504 9984
rect 6600 -9984 6738 9984
rect 6834 -9984 6972 9984
rect 7068 -9984 7206 9984
rect 7302 -9984 7440 9984
rect 7536 -9984 7674 9984
rect 7770 -9984 7908 9984
rect 8004 -9984 8142 9984
rect 8238 -9984 8376 9984
rect 8472 -9984 8610 9984
rect 8706 -9984 8844 9984
rect 8940 -9984 9078 9984
rect 9174 -9984 9312 9984
rect 9408 -9984 9546 9984
rect 9642 -9984 9780 9984
rect 9876 -9984 10014 9984
rect 10110 -9984 10248 9984
rect 10344 -9984 10482 9984
rect 10578 -9984 10716 9984
rect 10812 -9984 10950 9984
rect 11046 -9984 11184 9984
rect 11280 -9984 11418 9984
rect 11514 -9984 11652 9984
<< locali >>
rect -11782 10512 -11686 10546
rect 11686 10512 11782 10546
rect -11782 10450 -11748 10512
rect 11748 10450 11782 10512
rect -11782 -10512 -11748 -10450
rect 11748 -10512 11782 -10450
rect -11782 -10546 -11686 -10512
rect 11686 -10546 11782 -10512
<< viali >>
rect -11636 10001 -11530 10398
rect -11402 10001 -11296 10398
rect -11168 10001 -11062 10398
rect -10934 10001 -10828 10398
rect -10700 10001 -10594 10398
rect -10466 10001 -10360 10398
rect -10232 10001 -10126 10398
rect -9998 10001 -9892 10398
rect -9764 10001 -9658 10398
rect -9530 10001 -9424 10398
rect -9296 10001 -9190 10398
rect -9062 10001 -8956 10398
rect -8828 10001 -8722 10398
rect -8594 10001 -8488 10398
rect -8360 10001 -8254 10398
rect -8126 10001 -8020 10398
rect -7892 10001 -7786 10398
rect -7658 10001 -7552 10398
rect -7424 10001 -7318 10398
rect -7190 10001 -7084 10398
rect -6956 10001 -6850 10398
rect -6722 10001 -6616 10398
rect -6488 10001 -6382 10398
rect -6254 10001 -6148 10398
rect -6020 10001 -5914 10398
rect -5786 10001 -5680 10398
rect -5552 10001 -5446 10398
rect -5318 10001 -5212 10398
rect -5084 10001 -4978 10398
rect -4850 10001 -4744 10398
rect -4616 10001 -4510 10398
rect -4382 10001 -4276 10398
rect -4148 10001 -4042 10398
rect -3914 10001 -3808 10398
rect -3680 10001 -3574 10398
rect -3446 10001 -3340 10398
rect -3212 10001 -3106 10398
rect -2978 10001 -2872 10398
rect -2744 10001 -2638 10398
rect -2510 10001 -2404 10398
rect -2276 10001 -2170 10398
rect -2042 10001 -1936 10398
rect -1808 10001 -1702 10398
rect -1574 10001 -1468 10398
rect -1340 10001 -1234 10398
rect -1106 10001 -1000 10398
rect -872 10001 -766 10398
rect -638 10001 -532 10398
rect -404 10001 -298 10398
rect -170 10001 -64 10398
rect 64 10001 170 10398
rect 298 10001 404 10398
rect 532 10001 638 10398
rect 766 10001 872 10398
rect 1000 10001 1106 10398
rect 1234 10001 1340 10398
rect 1468 10001 1574 10398
rect 1702 10001 1808 10398
rect 1936 10001 2042 10398
rect 2170 10001 2276 10398
rect 2404 10001 2510 10398
rect 2638 10001 2744 10398
rect 2872 10001 2978 10398
rect 3106 10001 3212 10398
rect 3340 10001 3446 10398
rect 3574 10001 3680 10398
rect 3808 10001 3914 10398
rect 4042 10001 4148 10398
rect 4276 10001 4382 10398
rect 4510 10001 4616 10398
rect 4744 10001 4850 10398
rect 4978 10001 5084 10398
rect 5212 10001 5318 10398
rect 5446 10001 5552 10398
rect 5680 10001 5786 10398
rect 5914 10001 6020 10398
rect 6148 10001 6254 10398
rect 6382 10001 6488 10398
rect 6616 10001 6722 10398
rect 6850 10001 6956 10398
rect 7084 10001 7190 10398
rect 7318 10001 7424 10398
rect 7552 10001 7658 10398
rect 7786 10001 7892 10398
rect 8020 10001 8126 10398
rect 8254 10001 8360 10398
rect 8488 10001 8594 10398
rect 8722 10001 8828 10398
rect 8956 10001 9062 10398
rect 9190 10001 9296 10398
rect 9424 10001 9530 10398
rect 9658 10001 9764 10398
rect 9892 10001 9998 10398
rect 10126 10001 10232 10398
rect 10360 10001 10466 10398
rect 10594 10001 10700 10398
rect 10828 10001 10934 10398
rect 11062 10001 11168 10398
rect 11296 10001 11402 10398
rect 11530 10001 11636 10398
rect -11636 -10398 -11530 -10001
rect -11402 -10398 -11296 -10001
rect -11168 -10398 -11062 -10001
rect -10934 -10398 -10828 -10001
rect -10700 -10398 -10594 -10001
rect -10466 -10398 -10360 -10001
rect -10232 -10398 -10126 -10001
rect -9998 -10398 -9892 -10001
rect -9764 -10398 -9658 -10001
rect -9530 -10398 -9424 -10001
rect -9296 -10398 -9190 -10001
rect -9062 -10398 -8956 -10001
rect -8828 -10398 -8722 -10001
rect -8594 -10398 -8488 -10001
rect -8360 -10398 -8254 -10001
rect -8126 -10398 -8020 -10001
rect -7892 -10398 -7786 -10001
rect -7658 -10398 -7552 -10001
rect -7424 -10398 -7318 -10001
rect -7190 -10398 -7084 -10001
rect -6956 -10398 -6850 -10001
rect -6722 -10398 -6616 -10001
rect -6488 -10398 -6382 -10001
rect -6254 -10398 -6148 -10001
rect -6020 -10398 -5914 -10001
rect -5786 -10398 -5680 -10001
rect -5552 -10398 -5446 -10001
rect -5318 -10398 -5212 -10001
rect -5084 -10398 -4978 -10001
rect -4850 -10398 -4744 -10001
rect -4616 -10398 -4510 -10001
rect -4382 -10398 -4276 -10001
rect -4148 -10398 -4042 -10001
rect -3914 -10398 -3808 -10001
rect -3680 -10398 -3574 -10001
rect -3446 -10398 -3340 -10001
rect -3212 -10398 -3106 -10001
rect -2978 -10398 -2872 -10001
rect -2744 -10398 -2638 -10001
rect -2510 -10398 -2404 -10001
rect -2276 -10398 -2170 -10001
rect -2042 -10398 -1936 -10001
rect -1808 -10398 -1702 -10001
rect -1574 -10398 -1468 -10001
rect -1340 -10398 -1234 -10001
rect -1106 -10398 -1000 -10001
rect -872 -10398 -766 -10001
rect -638 -10398 -532 -10001
rect -404 -10398 -298 -10001
rect -170 -10398 -64 -10001
rect 64 -10398 170 -10001
rect 298 -10398 404 -10001
rect 532 -10398 638 -10001
rect 766 -10398 872 -10001
rect 1000 -10398 1106 -10001
rect 1234 -10398 1340 -10001
rect 1468 -10398 1574 -10001
rect 1702 -10398 1808 -10001
rect 1936 -10398 2042 -10001
rect 2170 -10398 2276 -10001
rect 2404 -10398 2510 -10001
rect 2638 -10398 2744 -10001
rect 2872 -10398 2978 -10001
rect 3106 -10398 3212 -10001
rect 3340 -10398 3446 -10001
rect 3574 -10398 3680 -10001
rect 3808 -10398 3914 -10001
rect 4042 -10398 4148 -10001
rect 4276 -10398 4382 -10001
rect 4510 -10398 4616 -10001
rect 4744 -10398 4850 -10001
rect 4978 -10398 5084 -10001
rect 5212 -10398 5318 -10001
rect 5446 -10398 5552 -10001
rect 5680 -10398 5786 -10001
rect 5914 -10398 6020 -10001
rect 6148 -10398 6254 -10001
rect 6382 -10398 6488 -10001
rect 6616 -10398 6722 -10001
rect 6850 -10398 6956 -10001
rect 7084 -10398 7190 -10001
rect 7318 -10398 7424 -10001
rect 7552 -10398 7658 -10001
rect 7786 -10398 7892 -10001
rect 8020 -10398 8126 -10001
rect 8254 -10398 8360 -10001
rect 8488 -10398 8594 -10001
rect 8722 -10398 8828 -10001
rect 8956 -10398 9062 -10001
rect 9190 -10398 9296 -10001
rect 9424 -10398 9530 -10001
rect 9658 -10398 9764 -10001
rect 9892 -10398 9998 -10001
rect 10126 -10398 10232 -10001
rect 10360 -10398 10466 -10001
rect 10594 -10398 10700 -10001
rect 10828 -10398 10934 -10001
rect 11062 -10398 11168 -10001
rect 11296 -10398 11402 -10001
rect 11530 -10398 11636 -10001
<< metal1 >>
rect -11642 10398 -11524 10410
rect -11642 10001 -11636 10398
rect -11530 10001 -11524 10398
rect -11642 9989 -11524 10001
rect -11408 10398 -11290 10410
rect -11408 10001 -11402 10398
rect -11296 10001 -11290 10398
rect -11408 9989 -11290 10001
rect -11174 10398 -11056 10410
rect -11174 10001 -11168 10398
rect -11062 10001 -11056 10398
rect -11174 9989 -11056 10001
rect -10940 10398 -10822 10410
rect -10940 10001 -10934 10398
rect -10828 10001 -10822 10398
rect -10940 9989 -10822 10001
rect -10706 10398 -10588 10410
rect -10706 10001 -10700 10398
rect -10594 10001 -10588 10398
rect -10706 9989 -10588 10001
rect -10472 10398 -10354 10410
rect -10472 10001 -10466 10398
rect -10360 10001 -10354 10398
rect -10472 9989 -10354 10001
rect -10238 10398 -10120 10410
rect -10238 10001 -10232 10398
rect -10126 10001 -10120 10398
rect -10238 9989 -10120 10001
rect -10004 10398 -9886 10410
rect -10004 10001 -9998 10398
rect -9892 10001 -9886 10398
rect -10004 9989 -9886 10001
rect -9770 10398 -9652 10410
rect -9770 10001 -9764 10398
rect -9658 10001 -9652 10398
rect -9770 9989 -9652 10001
rect -9536 10398 -9418 10410
rect -9536 10001 -9530 10398
rect -9424 10001 -9418 10398
rect -9536 9989 -9418 10001
rect -9302 10398 -9184 10410
rect -9302 10001 -9296 10398
rect -9190 10001 -9184 10398
rect -9302 9989 -9184 10001
rect -9068 10398 -8950 10410
rect -9068 10001 -9062 10398
rect -8956 10001 -8950 10398
rect -9068 9989 -8950 10001
rect -8834 10398 -8716 10410
rect -8834 10001 -8828 10398
rect -8722 10001 -8716 10398
rect -8834 9989 -8716 10001
rect -8600 10398 -8482 10410
rect -8600 10001 -8594 10398
rect -8488 10001 -8482 10398
rect -8600 9989 -8482 10001
rect -8366 10398 -8248 10410
rect -8366 10001 -8360 10398
rect -8254 10001 -8248 10398
rect -8366 9989 -8248 10001
rect -8132 10398 -8014 10410
rect -8132 10001 -8126 10398
rect -8020 10001 -8014 10398
rect -8132 9989 -8014 10001
rect -7898 10398 -7780 10410
rect -7898 10001 -7892 10398
rect -7786 10001 -7780 10398
rect -7898 9989 -7780 10001
rect -7664 10398 -7546 10410
rect -7664 10001 -7658 10398
rect -7552 10001 -7546 10398
rect -7664 9989 -7546 10001
rect -7430 10398 -7312 10410
rect -7430 10001 -7424 10398
rect -7318 10001 -7312 10398
rect -7430 9989 -7312 10001
rect -7196 10398 -7078 10410
rect -7196 10001 -7190 10398
rect -7084 10001 -7078 10398
rect -7196 9989 -7078 10001
rect -6962 10398 -6844 10410
rect -6962 10001 -6956 10398
rect -6850 10001 -6844 10398
rect -6962 9989 -6844 10001
rect -6728 10398 -6610 10410
rect -6728 10001 -6722 10398
rect -6616 10001 -6610 10398
rect -6728 9989 -6610 10001
rect -6494 10398 -6376 10410
rect -6494 10001 -6488 10398
rect -6382 10001 -6376 10398
rect -6494 9989 -6376 10001
rect -6260 10398 -6142 10410
rect -6260 10001 -6254 10398
rect -6148 10001 -6142 10398
rect -6260 9989 -6142 10001
rect -6026 10398 -5908 10410
rect -6026 10001 -6020 10398
rect -5914 10001 -5908 10398
rect -6026 9989 -5908 10001
rect -5792 10398 -5674 10410
rect -5792 10001 -5786 10398
rect -5680 10001 -5674 10398
rect -5792 9989 -5674 10001
rect -5558 10398 -5440 10410
rect -5558 10001 -5552 10398
rect -5446 10001 -5440 10398
rect -5558 9989 -5440 10001
rect -5324 10398 -5206 10410
rect -5324 10001 -5318 10398
rect -5212 10001 -5206 10398
rect -5324 9989 -5206 10001
rect -5090 10398 -4972 10410
rect -5090 10001 -5084 10398
rect -4978 10001 -4972 10398
rect -5090 9989 -4972 10001
rect -4856 10398 -4738 10410
rect -4856 10001 -4850 10398
rect -4744 10001 -4738 10398
rect -4856 9989 -4738 10001
rect -4622 10398 -4504 10410
rect -4622 10001 -4616 10398
rect -4510 10001 -4504 10398
rect -4622 9989 -4504 10001
rect -4388 10398 -4270 10410
rect -4388 10001 -4382 10398
rect -4276 10001 -4270 10398
rect -4388 9989 -4270 10001
rect -4154 10398 -4036 10410
rect -4154 10001 -4148 10398
rect -4042 10001 -4036 10398
rect -4154 9989 -4036 10001
rect -3920 10398 -3802 10410
rect -3920 10001 -3914 10398
rect -3808 10001 -3802 10398
rect -3920 9989 -3802 10001
rect -3686 10398 -3568 10410
rect -3686 10001 -3680 10398
rect -3574 10001 -3568 10398
rect -3686 9989 -3568 10001
rect -3452 10398 -3334 10410
rect -3452 10001 -3446 10398
rect -3340 10001 -3334 10398
rect -3452 9989 -3334 10001
rect -3218 10398 -3100 10410
rect -3218 10001 -3212 10398
rect -3106 10001 -3100 10398
rect -3218 9989 -3100 10001
rect -2984 10398 -2866 10410
rect -2984 10001 -2978 10398
rect -2872 10001 -2866 10398
rect -2984 9989 -2866 10001
rect -2750 10398 -2632 10410
rect -2750 10001 -2744 10398
rect -2638 10001 -2632 10398
rect -2750 9989 -2632 10001
rect -2516 10398 -2398 10410
rect -2516 10001 -2510 10398
rect -2404 10001 -2398 10398
rect -2516 9989 -2398 10001
rect -2282 10398 -2164 10410
rect -2282 10001 -2276 10398
rect -2170 10001 -2164 10398
rect -2282 9989 -2164 10001
rect -2048 10398 -1930 10410
rect -2048 10001 -2042 10398
rect -1936 10001 -1930 10398
rect -2048 9989 -1930 10001
rect -1814 10398 -1696 10410
rect -1814 10001 -1808 10398
rect -1702 10001 -1696 10398
rect -1814 9989 -1696 10001
rect -1580 10398 -1462 10410
rect -1580 10001 -1574 10398
rect -1468 10001 -1462 10398
rect -1580 9989 -1462 10001
rect -1346 10398 -1228 10410
rect -1346 10001 -1340 10398
rect -1234 10001 -1228 10398
rect -1346 9989 -1228 10001
rect -1112 10398 -994 10410
rect -1112 10001 -1106 10398
rect -1000 10001 -994 10398
rect -1112 9989 -994 10001
rect -878 10398 -760 10410
rect -878 10001 -872 10398
rect -766 10001 -760 10398
rect -878 9989 -760 10001
rect -644 10398 -526 10410
rect -644 10001 -638 10398
rect -532 10001 -526 10398
rect -644 9989 -526 10001
rect -410 10398 -292 10410
rect -410 10001 -404 10398
rect -298 10001 -292 10398
rect -410 9989 -292 10001
rect -176 10398 -58 10410
rect -176 10001 -170 10398
rect -64 10001 -58 10398
rect -176 9989 -58 10001
rect 58 10398 176 10410
rect 58 10001 64 10398
rect 170 10001 176 10398
rect 58 9989 176 10001
rect 292 10398 410 10410
rect 292 10001 298 10398
rect 404 10001 410 10398
rect 292 9989 410 10001
rect 526 10398 644 10410
rect 526 10001 532 10398
rect 638 10001 644 10398
rect 526 9989 644 10001
rect 760 10398 878 10410
rect 760 10001 766 10398
rect 872 10001 878 10398
rect 760 9989 878 10001
rect 994 10398 1112 10410
rect 994 10001 1000 10398
rect 1106 10001 1112 10398
rect 994 9989 1112 10001
rect 1228 10398 1346 10410
rect 1228 10001 1234 10398
rect 1340 10001 1346 10398
rect 1228 9989 1346 10001
rect 1462 10398 1580 10410
rect 1462 10001 1468 10398
rect 1574 10001 1580 10398
rect 1462 9989 1580 10001
rect 1696 10398 1814 10410
rect 1696 10001 1702 10398
rect 1808 10001 1814 10398
rect 1696 9989 1814 10001
rect 1930 10398 2048 10410
rect 1930 10001 1936 10398
rect 2042 10001 2048 10398
rect 1930 9989 2048 10001
rect 2164 10398 2282 10410
rect 2164 10001 2170 10398
rect 2276 10001 2282 10398
rect 2164 9989 2282 10001
rect 2398 10398 2516 10410
rect 2398 10001 2404 10398
rect 2510 10001 2516 10398
rect 2398 9989 2516 10001
rect 2632 10398 2750 10410
rect 2632 10001 2638 10398
rect 2744 10001 2750 10398
rect 2632 9989 2750 10001
rect 2866 10398 2984 10410
rect 2866 10001 2872 10398
rect 2978 10001 2984 10398
rect 2866 9989 2984 10001
rect 3100 10398 3218 10410
rect 3100 10001 3106 10398
rect 3212 10001 3218 10398
rect 3100 9989 3218 10001
rect 3334 10398 3452 10410
rect 3334 10001 3340 10398
rect 3446 10001 3452 10398
rect 3334 9989 3452 10001
rect 3568 10398 3686 10410
rect 3568 10001 3574 10398
rect 3680 10001 3686 10398
rect 3568 9989 3686 10001
rect 3802 10398 3920 10410
rect 3802 10001 3808 10398
rect 3914 10001 3920 10398
rect 3802 9989 3920 10001
rect 4036 10398 4154 10410
rect 4036 10001 4042 10398
rect 4148 10001 4154 10398
rect 4036 9989 4154 10001
rect 4270 10398 4388 10410
rect 4270 10001 4276 10398
rect 4382 10001 4388 10398
rect 4270 9989 4388 10001
rect 4504 10398 4622 10410
rect 4504 10001 4510 10398
rect 4616 10001 4622 10398
rect 4504 9989 4622 10001
rect 4738 10398 4856 10410
rect 4738 10001 4744 10398
rect 4850 10001 4856 10398
rect 4738 9989 4856 10001
rect 4972 10398 5090 10410
rect 4972 10001 4978 10398
rect 5084 10001 5090 10398
rect 4972 9989 5090 10001
rect 5206 10398 5324 10410
rect 5206 10001 5212 10398
rect 5318 10001 5324 10398
rect 5206 9989 5324 10001
rect 5440 10398 5558 10410
rect 5440 10001 5446 10398
rect 5552 10001 5558 10398
rect 5440 9989 5558 10001
rect 5674 10398 5792 10410
rect 5674 10001 5680 10398
rect 5786 10001 5792 10398
rect 5674 9989 5792 10001
rect 5908 10398 6026 10410
rect 5908 10001 5914 10398
rect 6020 10001 6026 10398
rect 5908 9989 6026 10001
rect 6142 10398 6260 10410
rect 6142 10001 6148 10398
rect 6254 10001 6260 10398
rect 6142 9989 6260 10001
rect 6376 10398 6494 10410
rect 6376 10001 6382 10398
rect 6488 10001 6494 10398
rect 6376 9989 6494 10001
rect 6610 10398 6728 10410
rect 6610 10001 6616 10398
rect 6722 10001 6728 10398
rect 6610 9989 6728 10001
rect 6844 10398 6962 10410
rect 6844 10001 6850 10398
rect 6956 10001 6962 10398
rect 6844 9989 6962 10001
rect 7078 10398 7196 10410
rect 7078 10001 7084 10398
rect 7190 10001 7196 10398
rect 7078 9989 7196 10001
rect 7312 10398 7430 10410
rect 7312 10001 7318 10398
rect 7424 10001 7430 10398
rect 7312 9989 7430 10001
rect 7546 10398 7664 10410
rect 7546 10001 7552 10398
rect 7658 10001 7664 10398
rect 7546 9989 7664 10001
rect 7780 10398 7898 10410
rect 7780 10001 7786 10398
rect 7892 10001 7898 10398
rect 7780 9989 7898 10001
rect 8014 10398 8132 10410
rect 8014 10001 8020 10398
rect 8126 10001 8132 10398
rect 8014 9989 8132 10001
rect 8248 10398 8366 10410
rect 8248 10001 8254 10398
rect 8360 10001 8366 10398
rect 8248 9989 8366 10001
rect 8482 10398 8600 10410
rect 8482 10001 8488 10398
rect 8594 10001 8600 10398
rect 8482 9989 8600 10001
rect 8716 10398 8834 10410
rect 8716 10001 8722 10398
rect 8828 10001 8834 10398
rect 8716 9989 8834 10001
rect 8950 10398 9068 10410
rect 8950 10001 8956 10398
rect 9062 10001 9068 10398
rect 8950 9989 9068 10001
rect 9184 10398 9302 10410
rect 9184 10001 9190 10398
rect 9296 10001 9302 10398
rect 9184 9989 9302 10001
rect 9418 10398 9536 10410
rect 9418 10001 9424 10398
rect 9530 10001 9536 10398
rect 9418 9989 9536 10001
rect 9652 10398 9770 10410
rect 9652 10001 9658 10398
rect 9764 10001 9770 10398
rect 9652 9989 9770 10001
rect 9886 10398 10004 10410
rect 9886 10001 9892 10398
rect 9998 10001 10004 10398
rect 9886 9989 10004 10001
rect 10120 10398 10238 10410
rect 10120 10001 10126 10398
rect 10232 10001 10238 10398
rect 10120 9989 10238 10001
rect 10354 10398 10472 10410
rect 10354 10001 10360 10398
rect 10466 10001 10472 10398
rect 10354 9989 10472 10001
rect 10588 10398 10706 10410
rect 10588 10001 10594 10398
rect 10700 10001 10706 10398
rect 10588 9989 10706 10001
rect 10822 10398 10940 10410
rect 10822 10001 10828 10398
rect 10934 10001 10940 10398
rect 10822 9989 10940 10001
rect 11056 10398 11174 10410
rect 11056 10001 11062 10398
rect 11168 10001 11174 10398
rect 11056 9989 11174 10001
rect 11290 10398 11408 10410
rect 11290 10001 11296 10398
rect 11402 10001 11408 10398
rect 11290 9989 11408 10001
rect 11524 10398 11642 10410
rect 11524 10001 11530 10398
rect 11636 10001 11642 10398
rect 11524 9989 11642 10001
rect -11642 -10001 -11524 -9989
rect -11642 -10398 -11636 -10001
rect -11530 -10398 -11524 -10001
rect -11642 -10410 -11524 -10398
rect -11408 -10001 -11290 -9989
rect -11408 -10398 -11402 -10001
rect -11296 -10398 -11290 -10001
rect -11408 -10410 -11290 -10398
rect -11174 -10001 -11056 -9989
rect -11174 -10398 -11168 -10001
rect -11062 -10398 -11056 -10001
rect -11174 -10410 -11056 -10398
rect -10940 -10001 -10822 -9989
rect -10940 -10398 -10934 -10001
rect -10828 -10398 -10822 -10001
rect -10940 -10410 -10822 -10398
rect -10706 -10001 -10588 -9989
rect -10706 -10398 -10700 -10001
rect -10594 -10398 -10588 -10001
rect -10706 -10410 -10588 -10398
rect -10472 -10001 -10354 -9989
rect -10472 -10398 -10466 -10001
rect -10360 -10398 -10354 -10001
rect -10472 -10410 -10354 -10398
rect -10238 -10001 -10120 -9989
rect -10238 -10398 -10232 -10001
rect -10126 -10398 -10120 -10001
rect -10238 -10410 -10120 -10398
rect -10004 -10001 -9886 -9989
rect -10004 -10398 -9998 -10001
rect -9892 -10398 -9886 -10001
rect -10004 -10410 -9886 -10398
rect -9770 -10001 -9652 -9989
rect -9770 -10398 -9764 -10001
rect -9658 -10398 -9652 -10001
rect -9770 -10410 -9652 -10398
rect -9536 -10001 -9418 -9989
rect -9536 -10398 -9530 -10001
rect -9424 -10398 -9418 -10001
rect -9536 -10410 -9418 -10398
rect -9302 -10001 -9184 -9989
rect -9302 -10398 -9296 -10001
rect -9190 -10398 -9184 -10001
rect -9302 -10410 -9184 -10398
rect -9068 -10001 -8950 -9989
rect -9068 -10398 -9062 -10001
rect -8956 -10398 -8950 -10001
rect -9068 -10410 -8950 -10398
rect -8834 -10001 -8716 -9989
rect -8834 -10398 -8828 -10001
rect -8722 -10398 -8716 -10001
rect -8834 -10410 -8716 -10398
rect -8600 -10001 -8482 -9989
rect -8600 -10398 -8594 -10001
rect -8488 -10398 -8482 -10001
rect -8600 -10410 -8482 -10398
rect -8366 -10001 -8248 -9989
rect -8366 -10398 -8360 -10001
rect -8254 -10398 -8248 -10001
rect -8366 -10410 -8248 -10398
rect -8132 -10001 -8014 -9989
rect -8132 -10398 -8126 -10001
rect -8020 -10398 -8014 -10001
rect -8132 -10410 -8014 -10398
rect -7898 -10001 -7780 -9989
rect -7898 -10398 -7892 -10001
rect -7786 -10398 -7780 -10001
rect -7898 -10410 -7780 -10398
rect -7664 -10001 -7546 -9989
rect -7664 -10398 -7658 -10001
rect -7552 -10398 -7546 -10001
rect -7664 -10410 -7546 -10398
rect -7430 -10001 -7312 -9989
rect -7430 -10398 -7424 -10001
rect -7318 -10398 -7312 -10001
rect -7430 -10410 -7312 -10398
rect -7196 -10001 -7078 -9989
rect -7196 -10398 -7190 -10001
rect -7084 -10398 -7078 -10001
rect -7196 -10410 -7078 -10398
rect -6962 -10001 -6844 -9989
rect -6962 -10398 -6956 -10001
rect -6850 -10398 -6844 -10001
rect -6962 -10410 -6844 -10398
rect -6728 -10001 -6610 -9989
rect -6728 -10398 -6722 -10001
rect -6616 -10398 -6610 -10001
rect -6728 -10410 -6610 -10398
rect -6494 -10001 -6376 -9989
rect -6494 -10398 -6488 -10001
rect -6382 -10398 -6376 -10001
rect -6494 -10410 -6376 -10398
rect -6260 -10001 -6142 -9989
rect -6260 -10398 -6254 -10001
rect -6148 -10398 -6142 -10001
rect -6260 -10410 -6142 -10398
rect -6026 -10001 -5908 -9989
rect -6026 -10398 -6020 -10001
rect -5914 -10398 -5908 -10001
rect -6026 -10410 -5908 -10398
rect -5792 -10001 -5674 -9989
rect -5792 -10398 -5786 -10001
rect -5680 -10398 -5674 -10001
rect -5792 -10410 -5674 -10398
rect -5558 -10001 -5440 -9989
rect -5558 -10398 -5552 -10001
rect -5446 -10398 -5440 -10001
rect -5558 -10410 -5440 -10398
rect -5324 -10001 -5206 -9989
rect -5324 -10398 -5318 -10001
rect -5212 -10398 -5206 -10001
rect -5324 -10410 -5206 -10398
rect -5090 -10001 -4972 -9989
rect -5090 -10398 -5084 -10001
rect -4978 -10398 -4972 -10001
rect -5090 -10410 -4972 -10398
rect -4856 -10001 -4738 -9989
rect -4856 -10398 -4850 -10001
rect -4744 -10398 -4738 -10001
rect -4856 -10410 -4738 -10398
rect -4622 -10001 -4504 -9989
rect -4622 -10398 -4616 -10001
rect -4510 -10398 -4504 -10001
rect -4622 -10410 -4504 -10398
rect -4388 -10001 -4270 -9989
rect -4388 -10398 -4382 -10001
rect -4276 -10398 -4270 -10001
rect -4388 -10410 -4270 -10398
rect -4154 -10001 -4036 -9989
rect -4154 -10398 -4148 -10001
rect -4042 -10398 -4036 -10001
rect -4154 -10410 -4036 -10398
rect -3920 -10001 -3802 -9989
rect -3920 -10398 -3914 -10001
rect -3808 -10398 -3802 -10001
rect -3920 -10410 -3802 -10398
rect -3686 -10001 -3568 -9989
rect -3686 -10398 -3680 -10001
rect -3574 -10398 -3568 -10001
rect -3686 -10410 -3568 -10398
rect -3452 -10001 -3334 -9989
rect -3452 -10398 -3446 -10001
rect -3340 -10398 -3334 -10001
rect -3452 -10410 -3334 -10398
rect -3218 -10001 -3100 -9989
rect -3218 -10398 -3212 -10001
rect -3106 -10398 -3100 -10001
rect -3218 -10410 -3100 -10398
rect -2984 -10001 -2866 -9989
rect -2984 -10398 -2978 -10001
rect -2872 -10398 -2866 -10001
rect -2984 -10410 -2866 -10398
rect -2750 -10001 -2632 -9989
rect -2750 -10398 -2744 -10001
rect -2638 -10398 -2632 -10001
rect -2750 -10410 -2632 -10398
rect -2516 -10001 -2398 -9989
rect -2516 -10398 -2510 -10001
rect -2404 -10398 -2398 -10001
rect -2516 -10410 -2398 -10398
rect -2282 -10001 -2164 -9989
rect -2282 -10398 -2276 -10001
rect -2170 -10398 -2164 -10001
rect -2282 -10410 -2164 -10398
rect -2048 -10001 -1930 -9989
rect -2048 -10398 -2042 -10001
rect -1936 -10398 -1930 -10001
rect -2048 -10410 -1930 -10398
rect -1814 -10001 -1696 -9989
rect -1814 -10398 -1808 -10001
rect -1702 -10398 -1696 -10001
rect -1814 -10410 -1696 -10398
rect -1580 -10001 -1462 -9989
rect -1580 -10398 -1574 -10001
rect -1468 -10398 -1462 -10001
rect -1580 -10410 -1462 -10398
rect -1346 -10001 -1228 -9989
rect -1346 -10398 -1340 -10001
rect -1234 -10398 -1228 -10001
rect -1346 -10410 -1228 -10398
rect -1112 -10001 -994 -9989
rect -1112 -10398 -1106 -10001
rect -1000 -10398 -994 -10001
rect -1112 -10410 -994 -10398
rect -878 -10001 -760 -9989
rect -878 -10398 -872 -10001
rect -766 -10398 -760 -10001
rect -878 -10410 -760 -10398
rect -644 -10001 -526 -9989
rect -644 -10398 -638 -10001
rect -532 -10398 -526 -10001
rect -644 -10410 -526 -10398
rect -410 -10001 -292 -9989
rect -410 -10398 -404 -10001
rect -298 -10398 -292 -10001
rect -410 -10410 -292 -10398
rect -176 -10001 -58 -9989
rect -176 -10398 -170 -10001
rect -64 -10398 -58 -10001
rect -176 -10410 -58 -10398
rect 58 -10001 176 -9989
rect 58 -10398 64 -10001
rect 170 -10398 176 -10001
rect 58 -10410 176 -10398
rect 292 -10001 410 -9989
rect 292 -10398 298 -10001
rect 404 -10398 410 -10001
rect 292 -10410 410 -10398
rect 526 -10001 644 -9989
rect 526 -10398 532 -10001
rect 638 -10398 644 -10001
rect 526 -10410 644 -10398
rect 760 -10001 878 -9989
rect 760 -10398 766 -10001
rect 872 -10398 878 -10001
rect 760 -10410 878 -10398
rect 994 -10001 1112 -9989
rect 994 -10398 1000 -10001
rect 1106 -10398 1112 -10001
rect 994 -10410 1112 -10398
rect 1228 -10001 1346 -9989
rect 1228 -10398 1234 -10001
rect 1340 -10398 1346 -10001
rect 1228 -10410 1346 -10398
rect 1462 -10001 1580 -9989
rect 1462 -10398 1468 -10001
rect 1574 -10398 1580 -10001
rect 1462 -10410 1580 -10398
rect 1696 -10001 1814 -9989
rect 1696 -10398 1702 -10001
rect 1808 -10398 1814 -10001
rect 1696 -10410 1814 -10398
rect 1930 -10001 2048 -9989
rect 1930 -10398 1936 -10001
rect 2042 -10398 2048 -10001
rect 1930 -10410 2048 -10398
rect 2164 -10001 2282 -9989
rect 2164 -10398 2170 -10001
rect 2276 -10398 2282 -10001
rect 2164 -10410 2282 -10398
rect 2398 -10001 2516 -9989
rect 2398 -10398 2404 -10001
rect 2510 -10398 2516 -10001
rect 2398 -10410 2516 -10398
rect 2632 -10001 2750 -9989
rect 2632 -10398 2638 -10001
rect 2744 -10398 2750 -10001
rect 2632 -10410 2750 -10398
rect 2866 -10001 2984 -9989
rect 2866 -10398 2872 -10001
rect 2978 -10398 2984 -10001
rect 2866 -10410 2984 -10398
rect 3100 -10001 3218 -9989
rect 3100 -10398 3106 -10001
rect 3212 -10398 3218 -10001
rect 3100 -10410 3218 -10398
rect 3334 -10001 3452 -9989
rect 3334 -10398 3340 -10001
rect 3446 -10398 3452 -10001
rect 3334 -10410 3452 -10398
rect 3568 -10001 3686 -9989
rect 3568 -10398 3574 -10001
rect 3680 -10398 3686 -10001
rect 3568 -10410 3686 -10398
rect 3802 -10001 3920 -9989
rect 3802 -10398 3808 -10001
rect 3914 -10398 3920 -10001
rect 3802 -10410 3920 -10398
rect 4036 -10001 4154 -9989
rect 4036 -10398 4042 -10001
rect 4148 -10398 4154 -10001
rect 4036 -10410 4154 -10398
rect 4270 -10001 4388 -9989
rect 4270 -10398 4276 -10001
rect 4382 -10398 4388 -10001
rect 4270 -10410 4388 -10398
rect 4504 -10001 4622 -9989
rect 4504 -10398 4510 -10001
rect 4616 -10398 4622 -10001
rect 4504 -10410 4622 -10398
rect 4738 -10001 4856 -9989
rect 4738 -10398 4744 -10001
rect 4850 -10398 4856 -10001
rect 4738 -10410 4856 -10398
rect 4972 -10001 5090 -9989
rect 4972 -10398 4978 -10001
rect 5084 -10398 5090 -10001
rect 4972 -10410 5090 -10398
rect 5206 -10001 5324 -9989
rect 5206 -10398 5212 -10001
rect 5318 -10398 5324 -10001
rect 5206 -10410 5324 -10398
rect 5440 -10001 5558 -9989
rect 5440 -10398 5446 -10001
rect 5552 -10398 5558 -10001
rect 5440 -10410 5558 -10398
rect 5674 -10001 5792 -9989
rect 5674 -10398 5680 -10001
rect 5786 -10398 5792 -10001
rect 5674 -10410 5792 -10398
rect 5908 -10001 6026 -9989
rect 5908 -10398 5914 -10001
rect 6020 -10398 6026 -10001
rect 5908 -10410 6026 -10398
rect 6142 -10001 6260 -9989
rect 6142 -10398 6148 -10001
rect 6254 -10398 6260 -10001
rect 6142 -10410 6260 -10398
rect 6376 -10001 6494 -9989
rect 6376 -10398 6382 -10001
rect 6488 -10398 6494 -10001
rect 6376 -10410 6494 -10398
rect 6610 -10001 6728 -9989
rect 6610 -10398 6616 -10001
rect 6722 -10398 6728 -10001
rect 6610 -10410 6728 -10398
rect 6844 -10001 6962 -9989
rect 6844 -10398 6850 -10001
rect 6956 -10398 6962 -10001
rect 6844 -10410 6962 -10398
rect 7078 -10001 7196 -9989
rect 7078 -10398 7084 -10001
rect 7190 -10398 7196 -10001
rect 7078 -10410 7196 -10398
rect 7312 -10001 7430 -9989
rect 7312 -10398 7318 -10001
rect 7424 -10398 7430 -10001
rect 7312 -10410 7430 -10398
rect 7546 -10001 7664 -9989
rect 7546 -10398 7552 -10001
rect 7658 -10398 7664 -10001
rect 7546 -10410 7664 -10398
rect 7780 -10001 7898 -9989
rect 7780 -10398 7786 -10001
rect 7892 -10398 7898 -10001
rect 7780 -10410 7898 -10398
rect 8014 -10001 8132 -9989
rect 8014 -10398 8020 -10001
rect 8126 -10398 8132 -10001
rect 8014 -10410 8132 -10398
rect 8248 -10001 8366 -9989
rect 8248 -10398 8254 -10001
rect 8360 -10398 8366 -10001
rect 8248 -10410 8366 -10398
rect 8482 -10001 8600 -9989
rect 8482 -10398 8488 -10001
rect 8594 -10398 8600 -10001
rect 8482 -10410 8600 -10398
rect 8716 -10001 8834 -9989
rect 8716 -10398 8722 -10001
rect 8828 -10398 8834 -10001
rect 8716 -10410 8834 -10398
rect 8950 -10001 9068 -9989
rect 8950 -10398 8956 -10001
rect 9062 -10398 9068 -10001
rect 8950 -10410 9068 -10398
rect 9184 -10001 9302 -9989
rect 9184 -10398 9190 -10001
rect 9296 -10398 9302 -10001
rect 9184 -10410 9302 -10398
rect 9418 -10001 9536 -9989
rect 9418 -10398 9424 -10001
rect 9530 -10398 9536 -10001
rect 9418 -10410 9536 -10398
rect 9652 -10001 9770 -9989
rect 9652 -10398 9658 -10001
rect 9764 -10398 9770 -10001
rect 9652 -10410 9770 -10398
rect 9886 -10001 10004 -9989
rect 9886 -10398 9892 -10001
rect 9998 -10398 10004 -10001
rect 9886 -10410 10004 -10398
rect 10120 -10001 10238 -9989
rect 10120 -10398 10126 -10001
rect 10232 -10398 10238 -10001
rect 10120 -10410 10238 -10398
rect 10354 -10001 10472 -9989
rect 10354 -10398 10360 -10001
rect 10466 -10398 10472 -10001
rect 10354 -10410 10472 -10398
rect 10588 -10001 10706 -9989
rect 10588 -10398 10594 -10001
rect 10700 -10398 10706 -10001
rect 10588 -10410 10706 -10398
rect 10822 -10001 10940 -9989
rect 10822 -10398 10828 -10001
rect 10934 -10398 10940 -10001
rect 10822 -10410 10940 -10398
rect 11056 -10001 11174 -9989
rect 11056 -10398 11062 -10001
rect 11168 -10398 11174 -10001
rect 11056 -10410 11174 -10398
rect 11290 -10001 11408 -9989
rect 11290 -10398 11296 -10001
rect 11402 -10398 11408 -10001
rect 11290 -10410 11408 -10398
rect 11524 -10001 11642 -9989
rect 11524 -10398 11530 -10001
rect 11636 -10398 11642 -10001
rect 11524 -10410 11642 -10398
<< properties >>
string FIXED_BBOX -11765 -10529 11765 10529
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 100.0 m 1 nx 100 wmin 0.690 lmin 0.50 class resistor rho 319.8 val 46.912k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
