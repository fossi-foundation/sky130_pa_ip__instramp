magic
tech sky130A
timestamp 1729620069
<< pwell >>
rect -164 -4642 164 4642
<< mvnmos >>
rect -50 4013 50 4513
rect -50 3404 50 3904
rect -50 2795 50 3295
rect -50 2186 50 2686
rect -50 1577 50 2077
rect -50 968 50 1468
rect -50 359 50 859
rect -50 -250 50 250
rect -50 -859 50 -359
rect -50 -1468 50 -968
rect -50 -2077 50 -1577
rect -50 -2686 50 -2186
rect -50 -3295 50 -2795
rect -50 -3904 50 -3404
rect -50 -4513 50 -4013
<< mvndiff >>
rect -79 4507 -50 4513
rect -79 4019 -73 4507
rect -56 4019 -50 4507
rect -79 4013 -50 4019
rect 50 4507 79 4513
rect 50 4019 56 4507
rect 73 4019 79 4507
rect 50 4013 79 4019
rect -79 3898 -50 3904
rect -79 3410 -73 3898
rect -56 3410 -50 3898
rect -79 3404 -50 3410
rect 50 3898 79 3904
rect 50 3410 56 3898
rect 73 3410 79 3898
rect 50 3404 79 3410
rect -79 3289 -50 3295
rect -79 2801 -73 3289
rect -56 2801 -50 3289
rect -79 2795 -50 2801
rect 50 3289 79 3295
rect 50 2801 56 3289
rect 73 2801 79 3289
rect 50 2795 79 2801
rect -79 2680 -50 2686
rect -79 2192 -73 2680
rect -56 2192 -50 2680
rect -79 2186 -50 2192
rect 50 2680 79 2686
rect 50 2192 56 2680
rect 73 2192 79 2680
rect 50 2186 79 2192
rect -79 2071 -50 2077
rect -79 1583 -73 2071
rect -56 1583 -50 2071
rect -79 1577 -50 1583
rect 50 2071 79 2077
rect 50 1583 56 2071
rect 73 1583 79 2071
rect 50 1577 79 1583
rect -79 1462 -50 1468
rect -79 974 -73 1462
rect -56 974 -50 1462
rect -79 968 -50 974
rect 50 1462 79 1468
rect 50 974 56 1462
rect 73 974 79 1462
rect 50 968 79 974
rect -79 853 -50 859
rect -79 365 -73 853
rect -56 365 -50 853
rect -79 359 -50 365
rect 50 853 79 859
rect 50 365 56 853
rect 73 365 79 853
rect 50 359 79 365
rect -79 244 -50 250
rect -79 -244 -73 244
rect -56 -244 -50 244
rect -79 -250 -50 -244
rect 50 244 79 250
rect 50 -244 56 244
rect 73 -244 79 244
rect 50 -250 79 -244
rect -79 -365 -50 -359
rect -79 -853 -73 -365
rect -56 -853 -50 -365
rect -79 -859 -50 -853
rect 50 -365 79 -359
rect 50 -853 56 -365
rect 73 -853 79 -365
rect 50 -859 79 -853
rect -79 -974 -50 -968
rect -79 -1462 -73 -974
rect -56 -1462 -50 -974
rect -79 -1468 -50 -1462
rect 50 -974 79 -968
rect 50 -1462 56 -974
rect 73 -1462 79 -974
rect 50 -1468 79 -1462
rect -79 -1583 -50 -1577
rect -79 -2071 -73 -1583
rect -56 -2071 -50 -1583
rect -79 -2077 -50 -2071
rect 50 -1583 79 -1577
rect 50 -2071 56 -1583
rect 73 -2071 79 -1583
rect 50 -2077 79 -2071
rect -79 -2192 -50 -2186
rect -79 -2680 -73 -2192
rect -56 -2680 -50 -2192
rect -79 -2686 -50 -2680
rect 50 -2192 79 -2186
rect 50 -2680 56 -2192
rect 73 -2680 79 -2192
rect 50 -2686 79 -2680
rect -79 -2801 -50 -2795
rect -79 -3289 -73 -2801
rect -56 -3289 -50 -2801
rect -79 -3295 -50 -3289
rect 50 -2801 79 -2795
rect 50 -3289 56 -2801
rect 73 -3289 79 -2801
rect 50 -3295 79 -3289
rect -79 -3410 -50 -3404
rect -79 -3898 -73 -3410
rect -56 -3898 -50 -3410
rect -79 -3904 -50 -3898
rect 50 -3410 79 -3404
rect 50 -3898 56 -3410
rect 73 -3898 79 -3410
rect 50 -3904 79 -3898
rect -79 -4019 -50 -4013
rect -79 -4507 -73 -4019
rect -56 -4507 -50 -4019
rect -79 -4513 -50 -4507
rect 50 -4019 79 -4013
rect 50 -4507 56 -4019
rect 73 -4507 79 -4019
rect 50 -4513 79 -4507
<< mvndiffc >>
rect -73 4019 -56 4507
rect 56 4019 73 4507
rect -73 3410 -56 3898
rect 56 3410 73 3898
rect -73 2801 -56 3289
rect 56 2801 73 3289
rect -73 2192 -56 2680
rect 56 2192 73 2680
rect -73 1583 -56 2071
rect 56 1583 73 2071
rect -73 974 -56 1462
rect 56 974 73 1462
rect -73 365 -56 853
rect 56 365 73 853
rect -73 -244 -56 244
rect 56 -244 73 244
rect -73 -853 -56 -365
rect 56 -853 73 -365
rect -73 -1462 -56 -974
rect 56 -1462 73 -974
rect -73 -2071 -56 -1583
rect 56 -2071 73 -1583
rect -73 -2680 -56 -2192
rect 56 -2680 73 -2192
rect -73 -3289 -56 -2801
rect 56 -3289 73 -2801
rect -73 -3898 -56 -3410
rect 56 -3898 73 -3410
rect -73 -4507 -56 -4019
rect 56 -4507 73 -4019
<< mvpsubdiff >>
rect -146 4618 146 4624
rect -146 4601 -92 4618
rect 92 4601 146 4618
rect -146 4595 146 4601
rect -146 4570 -117 4595
rect -146 -4570 -140 4570
rect -123 -4570 -117 4570
rect 117 4570 146 4595
rect -146 -4595 -117 -4570
rect 117 -4570 123 4570
rect 140 -4570 146 4570
rect 117 -4595 146 -4570
rect -146 -4601 146 -4595
rect -146 -4618 -92 -4601
rect 92 -4618 146 -4601
rect -146 -4624 146 -4618
<< mvpsubdiffcont >>
rect -92 4601 92 4618
rect -140 -4570 -123 4570
rect 123 -4570 140 4570
rect -92 -4618 92 -4601
<< poly >>
rect -50 4549 50 4557
rect -50 4532 -42 4549
rect 42 4532 50 4549
rect -50 4513 50 4532
rect -50 3994 50 4013
rect -50 3977 -42 3994
rect 42 3977 50 3994
rect -50 3969 50 3977
rect -50 3940 50 3948
rect -50 3923 -42 3940
rect 42 3923 50 3940
rect -50 3904 50 3923
rect -50 3385 50 3404
rect -50 3368 -42 3385
rect 42 3368 50 3385
rect -50 3360 50 3368
rect -50 3331 50 3339
rect -50 3314 -42 3331
rect 42 3314 50 3331
rect -50 3295 50 3314
rect -50 2776 50 2795
rect -50 2759 -42 2776
rect 42 2759 50 2776
rect -50 2751 50 2759
rect -50 2722 50 2730
rect -50 2705 -42 2722
rect 42 2705 50 2722
rect -50 2686 50 2705
rect -50 2167 50 2186
rect -50 2150 -42 2167
rect 42 2150 50 2167
rect -50 2142 50 2150
rect -50 2113 50 2121
rect -50 2096 -42 2113
rect 42 2096 50 2113
rect -50 2077 50 2096
rect -50 1558 50 1577
rect -50 1541 -42 1558
rect 42 1541 50 1558
rect -50 1533 50 1541
rect -50 1504 50 1512
rect -50 1487 -42 1504
rect 42 1487 50 1504
rect -50 1468 50 1487
rect -50 949 50 968
rect -50 932 -42 949
rect 42 932 50 949
rect -50 924 50 932
rect -50 895 50 903
rect -50 878 -42 895
rect 42 878 50 895
rect -50 859 50 878
rect -50 340 50 359
rect -50 323 -42 340
rect 42 323 50 340
rect -50 315 50 323
rect -50 286 50 294
rect -50 269 -42 286
rect 42 269 50 286
rect -50 250 50 269
rect -50 -269 50 -250
rect -50 -286 -42 -269
rect 42 -286 50 -269
rect -50 -294 50 -286
rect -50 -323 50 -315
rect -50 -340 -42 -323
rect 42 -340 50 -323
rect -50 -359 50 -340
rect -50 -878 50 -859
rect -50 -895 -42 -878
rect 42 -895 50 -878
rect -50 -903 50 -895
rect -50 -932 50 -924
rect -50 -949 -42 -932
rect 42 -949 50 -932
rect -50 -968 50 -949
rect -50 -1487 50 -1468
rect -50 -1504 -42 -1487
rect 42 -1504 50 -1487
rect -50 -1512 50 -1504
rect -50 -1541 50 -1533
rect -50 -1558 -42 -1541
rect 42 -1558 50 -1541
rect -50 -1577 50 -1558
rect -50 -2096 50 -2077
rect -50 -2113 -42 -2096
rect 42 -2113 50 -2096
rect -50 -2121 50 -2113
rect -50 -2150 50 -2142
rect -50 -2167 -42 -2150
rect 42 -2167 50 -2150
rect -50 -2186 50 -2167
rect -50 -2705 50 -2686
rect -50 -2722 -42 -2705
rect 42 -2722 50 -2705
rect -50 -2730 50 -2722
rect -50 -2759 50 -2751
rect -50 -2776 -42 -2759
rect 42 -2776 50 -2759
rect -50 -2795 50 -2776
rect -50 -3314 50 -3295
rect -50 -3331 -42 -3314
rect 42 -3331 50 -3314
rect -50 -3339 50 -3331
rect -50 -3368 50 -3360
rect -50 -3385 -42 -3368
rect 42 -3385 50 -3368
rect -50 -3404 50 -3385
rect -50 -3923 50 -3904
rect -50 -3940 -42 -3923
rect 42 -3940 50 -3923
rect -50 -3948 50 -3940
rect -50 -3977 50 -3969
rect -50 -3994 -42 -3977
rect 42 -3994 50 -3977
rect -50 -4013 50 -3994
rect -50 -4532 50 -4513
rect -50 -4549 -42 -4532
rect 42 -4549 50 -4532
rect -50 -4557 50 -4549
<< polycont >>
rect -42 4532 42 4549
rect -42 3977 42 3994
rect -42 3923 42 3940
rect -42 3368 42 3385
rect -42 3314 42 3331
rect -42 2759 42 2776
rect -42 2705 42 2722
rect -42 2150 42 2167
rect -42 2096 42 2113
rect -42 1541 42 1558
rect -42 1487 42 1504
rect -42 932 42 949
rect -42 878 42 895
rect -42 323 42 340
rect -42 269 42 286
rect -42 -286 42 -269
rect -42 -340 42 -323
rect -42 -895 42 -878
rect -42 -949 42 -932
rect -42 -1504 42 -1487
rect -42 -1558 42 -1541
rect -42 -2113 42 -2096
rect -42 -2167 42 -2150
rect -42 -2722 42 -2705
rect -42 -2776 42 -2759
rect -42 -3331 42 -3314
rect -42 -3385 42 -3368
rect -42 -3940 42 -3923
rect -42 -3994 42 -3977
rect -42 -4549 42 -4532
<< locali >>
rect -140 4601 -92 4618
rect 92 4601 140 4618
rect -140 4570 -123 4601
rect 123 4570 140 4601
rect -50 4532 -42 4549
rect 42 4532 50 4549
rect -73 4507 -56 4515
rect -73 4011 -56 4019
rect 56 4507 73 4515
rect 56 4011 73 4019
rect -50 3977 -42 3994
rect 42 3977 50 3994
rect -50 3923 -42 3940
rect 42 3923 50 3940
rect -73 3898 -56 3906
rect -73 3402 -56 3410
rect 56 3898 73 3906
rect 56 3402 73 3410
rect -50 3368 -42 3385
rect 42 3368 50 3385
rect -50 3314 -42 3331
rect 42 3314 50 3331
rect -73 3289 -56 3297
rect -73 2793 -56 2801
rect 56 3289 73 3297
rect 56 2793 73 2801
rect -50 2759 -42 2776
rect 42 2759 50 2776
rect -50 2705 -42 2722
rect 42 2705 50 2722
rect -73 2680 -56 2688
rect -73 2184 -56 2192
rect 56 2680 73 2688
rect 56 2184 73 2192
rect -50 2150 -42 2167
rect 42 2150 50 2167
rect -50 2096 -42 2113
rect 42 2096 50 2113
rect -73 2071 -56 2079
rect -73 1575 -56 1583
rect 56 2071 73 2079
rect 56 1575 73 1583
rect -50 1541 -42 1558
rect 42 1541 50 1558
rect -50 1487 -42 1504
rect 42 1487 50 1504
rect -73 1462 -56 1470
rect -73 966 -56 974
rect 56 1462 73 1470
rect 56 966 73 974
rect -50 932 -42 949
rect 42 932 50 949
rect -50 878 -42 895
rect 42 878 50 895
rect -73 853 -56 861
rect -73 357 -56 365
rect 56 853 73 861
rect 56 357 73 365
rect -50 323 -42 340
rect 42 323 50 340
rect -50 269 -42 286
rect 42 269 50 286
rect -73 244 -56 252
rect -73 -252 -56 -244
rect 56 244 73 252
rect 56 -252 73 -244
rect -50 -286 -42 -269
rect 42 -286 50 -269
rect -50 -340 -42 -323
rect 42 -340 50 -323
rect -73 -365 -56 -357
rect -73 -861 -56 -853
rect 56 -365 73 -357
rect 56 -861 73 -853
rect -50 -895 -42 -878
rect 42 -895 50 -878
rect -50 -949 -42 -932
rect 42 -949 50 -932
rect -73 -974 -56 -966
rect -73 -1470 -56 -1462
rect 56 -974 73 -966
rect 56 -1470 73 -1462
rect -50 -1504 -42 -1487
rect 42 -1504 50 -1487
rect -50 -1558 -42 -1541
rect 42 -1558 50 -1541
rect -73 -1583 -56 -1575
rect -73 -2079 -56 -2071
rect 56 -1583 73 -1575
rect 56 -2079 73 -2071
rect -50 -2113 -42 -2096
rect 42 -2113 50 -2096
rect -50 -2167 -42 -2150
rect 42 -2167 50 -2150
rect -73 -2192 -56 -2184
rect -73 -2688 -56 -2680
rect 56 -2192 73 -2184
rect 56 -2688 73 -2680
rect -50 -2722 -42 -2705
rect 42 -2722 50 -2705
rect -50 -2776 -42 -2759
rect 42 -2776 50 -2759
rect -73 -2801 -56 -2793
rect -73 -3297 -56 -3289
rect 56 -2801 73 -2793
rect 56 -3297 73 -3289
rect -50 -3331 -42 -3314
rect 42 -3331 50 -3314
rect -50 -3385 -42 -3368
rect 42 -3385 50 -3368
rect -73 -3410 -56 -3402
rect -73 -3906 -56 -3898
rect 56 -3410 73 -3402
rect 56 -3906 73 -3898
rect -50 -3940 -42 -3923
rect 42 -3940 50 -3923
rect -50 -3994 -42 -3977
rect 42 -3994 50 -3977
rect -73 -4019 -56 -4011
rect -73 -4515 -56 -4507
rect 56 -4019 73 -4011
rect 56 -4515 73 -4507
rect -50 -4549 -42 -4532
rect 42 -4549 50 -4532
rect -140 -4601 -123 -4570
rect 123 -4601 140 -4570
rect -140 -4618 -92 -4601
rect 92 -4618 140 -4601
<< viali >>
rect -42 4532 42 4549
rect -73 4019 -56 4507
rect 56 4019 73 4507
rect -42 3977 42 3994
rect -42 3923 42 3940
rect -73 3410 -56 3898
rect 56 3410 73 3898
rect -42 3368 42 3385
rect -42 3314 42 3331
rect -73 2801 -56 3289
rect 56 2801 73 3289
rect -42 2759 42 2776
rect -42 2705 42 2722
rect -73 2192 -56 2680
rect 56 2192 73 2680
rect -42 2150 42 2167
rect -42 2096 42 2113
rect -73 1583 -56 2071
rect 56 1583 73 2071
rect -42 1541 42 1558
rect -42 1487 42 1504
rect -73 974 -56 1462
rect 56 974 73 1462
rect -42 932 42 949
rect -42 878 42 895
rect -73 365 -56 853
rect 56 365 73 853
rect -42 323 42 340
rect -42 269 42 286
rect -73 -244 -56 244
rect 56 -244 73 244
rect -42 -286 42 -269
rect -42 -340 42 -323
rect -73 -853 -56 -365
rect 56 -853 73 -365
rect -42 -895 42 -878
rect -42 -949 42 -932
rect -73 -1462 -56 -974
rect 56 -1462 73 -974
rect -42 -1504 42 -1487
rect -42 -1558 42 -1541
rect -73 -2071 -56 -1583
rect 56 -2071 73 -1583
rect -42 -2113 42 -2096
rect -42 -2167 42 -2150
rect -73 -2680 -56 -2192
rect 56 -2680 73 -2192
rect -42 -2722 42 -2705
rect -42 -2776 42 -2759
rect -73 -3289 -56 -2801
rect 56 -3289 73 -2801
rect -42 -3331 42 -3314
rect -42 -3385 42 -3368
rect -73 -3898 -56 -3410
rect 56 -3898 73 -3410
rect -42 -3940 42 -3923
rect -42 -3994 42 -3977
rect -73 -4507 -56 -4019
rect 56 -4507 73 -4019
rect -42 -4549 42 -4532
<< metal1 >>
rect -48 4549 48 4552
rect -48 4532 -42 4549
rect 42 4532 48 4549
rect -48 4529 48 4532
rect -76 4507 -53 4513
rect -76 4019 -73 4507
rect -56 4019 -53 4507
rect -76 4013 -53 4019
rect 53 4507 76 4513
rect 53 4019 56 4507
rect 73 4019 76 4507
rect 53 4013 76 4019
rect -48 3994 48 3997
rect -48 3977 -42 3994
rect 42 3977 48 3994
rect -48 3974 48 3977
rect -48 3940 48 3943
rect -48 3923 -42 3940
rect 42 3923 48 3940
rect -48 3920 48 3923
rect -76 3898 -53 3904
rect -76 3410 -73 3898
rect -56 3410 -53 3898
rect -76 3404 -53 3410
rect 53 3898 76 3904
rect 53 3410 56 3898
rect 73 3410 76 3898
rect 53 3404 76 3410
rect -48 3385 48 3388
rect -48 3368 -42 3385
rect 42 3368 48 3385
rect -48 3365 48 3368
rect -48 3331 48 3334
rect -48 3314 -42 3331
rect 42 3314 48 3331
rect -48 3311 48 3314
rect -76 3289 -53 3295
rect -76 2801 -73 3289
rect -56 2801 -53 3289
rect -76 2795 -53 2801
rect 53 3289 76 3295
rect 53 2801 56 3289
rect 73 2801 76 3289
rect 53 2795 76 2801
rect -48 2776 48 2779
rect -48 2759 -42 2776
rect 42 2759 48 2776
rect -48 2756 48 2759
rect -48 2722 48 2725
rect -48 2705 -42 2722
rect 42 2705 48 2722
rect -48 2702 48 2705
rect -76 2680 -53 2686
rect -76 2192 -73 2680
rect -56 2192 -53 2680
rect -76 2186 -53 2192
rect 53 2680 76 2686
rect 53 2192 56 2680
rect 73 2192 76 2680
rect 53 2186 76 2192
rect -48 2167 48 2170
rect -48 2150 -42 2167
rect 42 2150 48 2167
rect -48 2147 48 2150
rect -48 2113 48 2116
rect -48 2096 -42 2113
rect 42 2096 48 2113
rect -48 2093 48 2096
rect -76 2071 -53 2077
rect -76 1583 -73 2071
rect -56 1583 -53 2071
rect -76 1577 -53 1583
rect 53 2071 76 2077
rect 53 1583 56 2071
rect 73 1583 76 2071
rect 53 1577 76 1583
rect -48 1558 48 1561
rect -48 1541 -42 1558
rect 42 1541 48 1558
rect -48 1538 48 1541
rect -48 1504 48 1507
rect -48 1487 -42 1504
rect 42 1487 48 1504
rect -48 1484 48 1487
rect -76 1462 -53 1468
rect -76 974 -73 1462
rect -56 974 -53 1462
rect -76 968 -53 974
rect 53 1462 76 1468
rect 53 974 56 1462
rect 73 974 76 1462
rect 53 968 76 974
rect -48 949 48 952
rect -48 932 -42 949
rect 42 932 48 949
rect -48 929 48 932
rect -48 895 48 898
rect -48 878 -42 895
rect 42 878 48 895
rect -48 875 48 878
rect -76 853 -53 859
rect -76 365 -73 853
rect -56 365 -53 853
rect -76 359 -53 365
rect 53 853 76 859
rect 53 365 56 853
rect 73 365 76 853
rect 53 359 76 365
rect -48 340 48 343
rect -48 323 -42 340
rect 42 323 48 340
rect -48 320 48 323
rect -48 286 48 289
rect -48 269 -42 286
rect 42 269 48 286
rect -48 266 48 269
rect -76 244 -53 250
rect -76 -244 -73 244
rect -56 -244 -53 244
rect -76 -250 -53 -244
rect 53 244 76 250
rect 53 -244 56 244
rect 73 -244 76 244
rect 53 -250 76 -244
rect -48 -269 48 -266
rect -48 -286 -42 -269
rect 42 -286 48 -269
rect -48 -289 48 -286
rect -48 -323 48 -320
rect -48 -340 -42 -323
rect 42 -340 48 -323
rect -48 -343 48 -340
rect -76 -365 -53 -359
rect -76 -853 -73 -365
rect -56 -853 -53 -365
rect -76 -859 -53 -853
rect 53 -365 76 -359
rect 53 -853 56 -365
rect 73 -853 76 -365
rect 53 -859 76 -853
rect -48 -878 48 -875
rect -48 -895 -42 -878
rect 42 -895 48 -878
rect -48 -898 48 -895
rect -48 -932 48 -929
rect -48 -949 -42 -932
rect 42 -949 48 -932
rect -48 -952 48 -949
rect -76 -974 -53 -968
rect -76 -1462 -73 -974
rect -56 -1462 -53 -974
rect -76 -1468 -53 -1462
rect 53 -974 76 -968
rect 53 -1462 56 -974
rect 73 -1462 76 -974
rect 53 -1468 76 -1462
rect -48 -1487 48 -1484
rect -48 -1504 -42 -1487
rect 42 -1504 48 -1487
rect -48 -1507 48 -1504
rect -48 -1541 48 -1538
rect -48 -1558 -42 -1541
rect 42 -1558 48 -1541
rect -48 -1561 48 -1558
rect -76 -1583 -53 -1577
rect -76 -2071 -73 -1583
rect -56 -2071 -53 -1583
rect -76 -2077 -53 -2071
rect 53 -1583 76 -1577
rect 53 -2071 56 -1583
rect 73 -2071 76 -1583
rect 53 -2077 76 -2071
rect -48 -2096 48 -2093
rect -48 -2113 -42 -2096
rect 42 -2113 48 -2096
rect -48 -2116 48 -2113
rect -48 -2150 48 -2147
rect -48 -2167 -42 -2150
rect 42 -2167 48 -2150
rect -48 -2170 48 -2167
rect -76 -2192 -53 -2186
rect -76 -2680 -73 -2192
rect -56 -2680 -53 -2192
rect -76 -2686 -53 -2680
rect 53 -2192 76 -2186
rect 53 -2680 56 -2192
rect 73 -2680 76 -2192
rect 53 -2686 76 -2680
rect -48 -2705 48 -2702
rect -48 -2722 -42 -2705
rect 42 -2722 48 -2705
rect -48 -2725 48 -2722
rect -48 -2759 48 -2756
rect -48 -2776 -42 -2759
rect 42 -2776 48 -2759
rect -48 -2779 48 -2776
rect -76 -2801 -53 -2795
rect -76 -3289 -73 -2801
rect -56 -3289 -53 -2801
rect -76 -3295 -53 -3289
rect 53 -2801 76 -2795
rect 53 -3289 56 -2801
rect 73 -3289 76 -2801
rect 53 -3295 76 -3289
rect -48 -3314 48 -3311
rect -48 -3331 -42 -3314
rect 42 -3331 48 -3314
rect -48 -3334 48 -3331
rect -48 -3368 48 -3365
rect -48 -3385 -42 -3368
rect 42 -3385 48 -3368
rect -48 -3388 48 -3385
rect -76 -3410 -53 -3404
rect -76 -3898 -73 -3410
rect -56 -3898 -53 -3410
rect -76 -3904 -53 -3898
rect 53 -3410 76 -3404
rect 53 -3898 56 -3410
rect 73 -3898 76 -3410
rect 53 -3904 76 -3898
rect -48 -3923 48 -3920
rect -48 -3940 -42 -3923
rect 42 -3940 48 -3923
rect -48 -3943 48 -3940
rect -48 -3977 48 -3974
rect -48 -3994 -42 -3977
rect 42 -3994 48 -3977
rect -48 -3997 48 -3994
rect -76 -4019 -53 -4013
rect -76 -4507 -73 -4019
rect -56 -4507 -53 -4019
rect -76 -4513 -53 -4507
rect 53 -4019 76 -4013
rect 53 -4507 56 -4019
rect 73 -4507 76 -4019
rect 53 -4513 76 -4507
rect -48 -4532 48 -4529
rect -48 -4549 -42 -4532
rect 42 -4549 48 -4532
rect -48 -4552 48 -4549
<< properties >>
string FIXED_BBOX -131 -4609 131 4609
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 1.0 m 15 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 ad {int((nf+1)/2) * W/nf * 0.29} as {int((nf+2)/2) * W/nf * 0.29} pd {2*int((nf+1)/2) * (W/nf + 0.29)} ps {2*int((nf+2)/2) * (W/nf + 0.29)} nrd {0.29 / W} nrs {0.29 / W} sa 0 sb 0 sd 0 mult 15
<< end >>
