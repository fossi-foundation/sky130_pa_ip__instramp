magic
tech sky130A
magscale 1 2
timestamp 1730948043
<< pwell >>
rect -616 -1582 616 1582
<< psubdiff >>
rect -580 1512 -484 1546
rect 484 1512 580 1546
rect -580 1450 -546 1512
rect 546 1450 580 1512
rect -580 -1512 -546 -1450
rect 546 -1512 580 -1450
rect -580 -1546 -484 -1512
rect 484 -1546 580 -1512
<< psubdiffcont >>
rect -484 1512 484 1546
rect -580 -1450 -546 1450
rect 546 -1450 580 1450
rect -484 -1546 484 -1512
<< xpolycontact >>
rect -450 984 -380 1416
rect -450 -1416 -380 -984
rect -284 984 -214 1416
rect -284 -1416 -214 -984
rect -118 984 -48 1416
rect -118 -1416 -48 -984
rect 48 984 118 1416
rect 48 -1416 118 -984
rect 214 984 284 1416
rect 214 -1416 284 -984
rect 380 984 450 1416
rect 380 -1416 450 -984
<< xpolyres >>
rect -450 -984 -380 984
rect -284 -984 -214 984
rect -118 -984 -48 984
rect 48 -984 118 984
rect 214 -984 284 984
rect 380 -984 450 984
<< locali >>
rect -580 1512 -484 1546
rect 484 1512 580 1546
rect -580 1450 -546 1512
rect 546 1450 580 1512
rect -580 -1512 -546 -1450
rect 546 -1512 580 -1450
rect -580 -1546 -484 -1512
rect 484 -1546 580 -1512
<< viali >>
rect -434 1001 -396 1398
rect -268 1001 -230 1398
rect -102 1001 -64 1398
rect 64 1001 102 1398
rect 230 1001 268 1398
rect 396 1001 434 1398
rect -434 -1398 -396 -1001
rect -268 -1398 -230 -1001
rect -102 -1398 -64 -1001
rect 64 -1398 102 -1001
rect 230 -1398 268 -1001
rect 396 -1398 434 -1001
<< metal1 >>
rect -440 1398 -390 1410
rect -440 1001 -434 1398
rect -396 1001 -390 1398
rect -440 989 -390 1001
rect -274 1398 -224 1410
rect -274 1001 -268 1398
rect -230 1001 -224 1398
rect -274 989 -224 1001
rect -108 1398 -58 1410
rect -108 1001 -102 1398
rect -64 1001 -58 1398
rect -108 989 -58 1001
rect 58 1398 108 1410
rect 58 1001 64 1398
rect 102 1001 108 1398
rect 58 989 108 1001
rect 224 1398 274 1410
rect 224 1001 230 1398
rect 268 1001 274 1398
rect 224 989 274 1001
rect 390 1398 440 1410
rect 390 1001 396 1398
rect 434 1001 440 1398
rect 390 989 440 1001
rect -440 -1001 -390 -989
rect -440 -1398 -434 -1001
rect -396 -1398 -390 -1001
rect -440 -1410 -390 -1398
rect -274 -1001 -224 -989
rect -274 -1398 -268 -1001
rect -230 -1398 -224 -1001
rect -274 -1410 -224 -1398
rect -108 -1001 -58 -989
rect -108 -1398 -102 -1001
rect -64 -1398 -58 -1001
rect -108 -1410 -58 -1398
rect 58 -1001 108 -989
rect 58 -1398 64 -1001
rect 102 -1398 108 -1001
rect 58 -1410 108 -1398
rect 224 -1001 274 -989
rect 224 -1398 230 -1001
rect 268 -1398 274 -1001
rect 224 -1410 274 -1398
rect 390 -1001 440 -989
rect 390 -1398 396 -1001
rect 434 -1398 440 -1001
rect 390 -1410 440 -1398
<< properties >>
string FIXED_BBOX -563 -1529 563 1529
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 10 m 1 nx 6 wmin 0.350 lmin 0.50 class resistor rho 2000 val 58.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
