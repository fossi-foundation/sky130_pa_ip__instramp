magic
tech sky130A
magscale 1 2
timestamp 1729620069
<< pwell >>
rect -1084 -2585 1084 2585
<< mvnmos >>
rect -856 1327 -656 2327
rect -478 1327 -278 2327
rect -100 1327 100 2327
rect 278 1327 478 2327
rect 656 1327 856 2327
rect -856 109 -656 1109
rect -478 109 -278 1109
rect -100 109 100 1109
rect 278 109 478 1109
rect 656 109 856 1109
rect -856 -1109 -656 -109
rect -478 -1109 -278 -109
rect -100 -1109 100 -109
rect 278 -1109 478 -109
rect 656 -1109 856 -109
rect -856 -2327 -656 -1327
rect -478 -2327 -278 -1327
rect -100 -2327 100 -1327
rect 278 -2327 478 -1327
rect 656 -2327 856 -1327
<< mvndiff >>
rect -914 2315 -856 2327
rect -914 1339 -902 2315
rect -868 1339 -856 2315
rect -914 1327 -856 1339
rect -656 2315 -598 2327
rect -656 1339 -644 2315
rect -610 1339 -598 2315
rect -656 1327 -598 1339
rect -536 2315 -478 2327
rect -536 1339 -524 2315
rect -490 1339 -478 2315
rect -536 1327 -478 1339
rect -278 2315 -220 2327
rect -278 1339 -266 2315
rect -232 1339 -220 2315
rect -278 1327 -220 1339
rect -158 2315 -100 2327
rect -158 1339 -146 2315
rect -112 1339 -100 2315
rect -158 1327 -100 1339
rect 100 2315 158 2327
rect 100 1339 112 2315
rect 146 1339 158 2315
rect 100 1327 158 1339
rect 220 2315 278 2327
rect 220 1339 232 2315
rect 266 1339 278 2315
rect 220 1327 278 1339
rect 478 2315 536 2327
rect 478 1339 490 2315
rect 524 1339 536 2315
rect 478 1327 536 1339
rect 598 2315 656 2327
rect 598 1339 610 2315
rect 644 1339 656 2315
rect 598 1327 656 1339
rect 856 2315 914 2327
rect 856 1339 868 2315
rect 902 1339 914 2315
rect 856 1327 914 1339
rect -914 1097 -856 1109
rect -914 121 -902 1097
rect -868 121 -856 1097
rect -914 109 -856 121
rect -656 1097 -598 1109
rect -656 121 -644 1097
rect -610 121 -598 1097
rect -656 109 -598 121
rect -536 1097 -478 1109
rect -536 121 -524 1097
rect -490 121 -478 1097
rect -536 109 -478 121
rect -278 1097 -220 1109
rect -278 121 -266 1097
rect -232 121 -220 1097
rect -278 109 -220 121
rect -158 1097 -100 1109
rect -158 121 -146 1097
rect -112 121 -100 1097
rect -158 109 -100 121
rect 100 1097 158 1109
rect 100 121 112 1097
rect 146 121 158 1097
rect 100 109 158 121
rect 220 1097 278 1109
rect 220 121 232 1097
rect 266 121 278 1097
rect 220 109 278 121
rect 478 1097 536 1109
rect 478 121 490 1097
rect 524 121 536 1097
rect 478 109 536 121
rect 598 1097 656 1109
rect 598 121 610 1097
rect 644 121 656 1097
rect 598 109 656 121
rect 856 1097 914 1109
rect 856 121 868 1097
rect 902 121 914 1097
rect 856 109 914 121
rect -914 -121 -856 -109
rect -914 -1097 -902 -121
rect -868 -1097 -856 -121
rect -914 -1109 -856 -1097
rect -656 -121 -598 -109
rect -656 -1097 -644 -121
rect -610 -1097 -598 -121
rect -656 -1109 -598 -1097
rect -536 -121 -478 -109
rect -536 -1097 -524 -121
rect -490 -1097 -478 -121
rect -536 -1109 -478 -1097
rect -278 -121 -220 -109
rect -278 -1097 -266 -121
rect -232 -1097 -220 -121
rect -278 -1109 -220 -1097
rect -158 -121 -100 -109
rect -158 -1097 -146 -121
rect -112 -1097 -100 -121
rect -158 -1109 -100 -1097
rect 100 -121 158 -109
rect 100 -1097 112 -121
rect 146 -1097 158 -121
rect 100 -1109 158 -1097
rect 220 -121 278 -109
rect 220 -1097 232 -121
rect 266 -1097 278 -121
rect 220 -1109 278 -1097
rect 478 -121 536 -109
rect 478 -1097 490 -121
rect 524 -1097 536 -121
rect 478 -1109 536 -1097
rect 598 -121 656 -109
rect 598 -1097 610 -121
rect 644 -1097 656 -121
rect 598 -1109 656 -1097
rect 856 -121 914 -109
rect 856 -1097 868 -121
rect 902 -1097 914 -121
rect 856 -1109 914 -1097
rect -914 -1339 -856 -1327
rect -914 -2315 -902 -1339
rect -868 -2315 -856 -1339
rect -914 -2327 -856 -2315
rect -656 -1339 -598 -1327
rect -656 -2315 -644 -1339
rect -610 -2315 -598 -1339
rect -656 -2327 -598 -2315
rect -536 -1339 -478 -1327
rect -536 -2315 -524 -1339
rect -490 -2315 -478 -1339
rect -536 -2327 -478 -2315
rect -278 -1339 -220 -1327
rect -278 -2315 -266 -1339
rect -232 -2315 -220 -1339
rect -278 -2327 -220 -2315
rect -158 -1339 -100 -1327
rect -158 -2315 -146 -1339
rect -112 -2315 -100 -1339
rect -158 -2327 -100 -2315
rect 100 -1339 158 -1327
rect 100 -2315 112 -1339
rect 146 -2315 158 -1339
rect 100 -2327 158 -2315
rect 220 -1339 278 -1327
rect 220 -2315 232 -1339
rect 266 -2315 278 -1339
rect 220 -2327 278 -2315
rect 478 -1339 536 -1327
rect 478 -2315 490 -1339
rect 524 -2315 536 -1339
rect 478 -2327 536 -2315
rect 598 -1339 656 -1327
rect 598 -2315 610 -1339
rect 644 -2315 656 -1339
rect 598 -2327 656 -2315
rect 856 -1339 914 -1327
rect 856 -2315 868 -1339
rect 902 -2315 914 -1339
rect 856 -2327 914 -2315
<< mvndiffc >>
rect -902 1339 -868 2315
rect -644 1339 -610 2315
rect -524 1339 -490 2315
rect -266 1339 -232 2315
rect -146 1339 -112 2315
rect 112 1339 146 2315
rect 232 1339 266 2315
rect 490 1339 524 2315
rect 610 1339 644 2315
rect 868 1339 902 2315
rect -902 121 -868 1097
rect -644 121 -610 1097
rect -524 121 -490 1097
rect -266 121 -232 1097
rect -146 121 -112 1097
rect 112 121 146 1097
rect 232 121 266 1097
rect 490 121 524 1097
rect 610 121 644 1097
rect 868 121 902 1097
rect -902 -1097 -868 -121
rect -644 -1097 -610 -121
rect -524 -1097 -490 -121
rect -266 -1097 -232 -121
rect -146 -1097 -112 -121
rect 112 -1097 146 -121
rect 232 -1097 266 -121
rect 490 -1097 524 -121
rect 610 -1097 644 -121
rect 868 -1097 902 -121
rect -902 -2315 -868 -1339
rect -644 -2315 -610 -1339
rect -524 -2315 -490 -1339
rect -266 -2315 -232 -1339
rect -146 -2315 -112 -1339
rect 112 -2315 146 -1339
rect 232 -2315 266 -1339
rect 490 -2315 524 -1339
rect 610 -2315 644 -1339
rect 868 -2315 902 -1339
<< mvpsubdiff >>
rect -1048 2537 1048 2549
rect -1048 2503 -940 2537
rect 940 2503 1048 2537
rect -1048 2491 1048 2503
rect -1048 2441 -990 2491
rect -1048 -2441 -1036 2441
rect -1002 -2441 -990 2441
rect 990 2441 1048 2491
rect -1048 -2491 -990 -2441
rect 990 -2441 1002 2441
rect 1036 -2441 1048 2441
rect 990 -2491 1048 -2441
rect -1048 -2503 1048 -2491
rect -1048 -2537 -940 -2503
rect 940 -2537 1048 -2503
rect -1048 -2549 1048 -2537
<< mvpsubdiffcont >>
rect -940 2503 940 2537
rect -1036 -2441 -1002 2441
rect 1002 -2441 1036 2441
rect -940 -2537 940 -2503
<< poly >>
rect -856 2399 -656 2415
rect -856 2365 -840 2399
rect -672 2365 -656 2399
rect -856 2327 -656 2365
rect -478 2399 -278 2415
rect -478 2365 -462 2399
rect -294 2365 -278 2399
rect -478 2327 -278 2365
rect -100 2399 100 2415
rect -100 2365 -84 2399
rect 84 2365 100 2399
rect -100 2327 100 2365
rect 278 2399 478 2415
rect 278 2365 294 2399
rect 462 2365 478 2399
rect 278 2327 478 2365
rect 656 2399 856 2415
rect 656 2365 672 2399
rect 840 2365 856 2399
rect 656 2327 856 2365
rect -856 1289 -656 1327
rect -856 1255 -840 1289
rect -672 1255 -656 1289
rect -856 1239 -656 1255
rect -478 1289 -278 1327
rect -478 1255 -462 1289
rect -294 1255 -278 1289
rect -478 1239 -278 1255
rect -100 1289 100 1327
rect -100 1255 -84 1289
rect 84 1255 100 1289
rect -100 1239 100 1255
rect 278 1289 478 1327
rect 278 1255 294 1289
rect 462 1255 478 1289
rect 278 1239 478 1255
rect 656 1289 856 1327
rect 656 1255 672 1289
rect 840 1255 856 1289
rect 656 1239 856 1255
rect -856 1181 -656 1197
rect -856 1147 -840 1181
rect -672 1147 -656 1181
rect -856 1109 -656 1147
rect -478 1181 -278 1197
rect -478 1147 -462 1181
rect -294 1147 -278 1181
rect -478 1109 -278 1147
rect -100 1181 100 1197
rect -100 1147 -84 1181
rect 84 1147 100 1181
rect -100 1109 100 1147
rect 278 1181 478 1197
rect 278 1147 294 1181
rect 462 1147 478 1181
rect 278 1109 478 1147
rect 656 1181 856 1197
rect 656 1147 672 1181
rect 840 1147 856 1181
rect 656 1109 856 1147
rect -856 71 -656 109
rect -856 37 -840 71
rect -672 37 -656 71
rect -856 21 -656 37
rect -478 71 -278 109
rect -478 37 -462 71
rect -294 37 -278 71
rect -478 21 -278 37
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect 278 71 478 109
rect 278 37 294 71
rect 462 37 478 71
rect 278 21 478 37
rect 656 71 856 109
rect 656 37 672 71
rect 840 37 856 71
rect 656 21 856 37
rect -856 -37 -656 -21
rect -856 -71 -840 -37
rect -672 -71 -656 -37
rect -856 -109 -656 -71
rect -478 -37 -278 -21
rect -478 -71 -462 -37
rect -294 -71 -278 -37
rect -478 -109 -278 -71
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect 278 -37 478 -21
rect 278 -71 294 -37
rect 462 -71 478 -37
rect 278 -109 478 -71
rect 656 -37 856 -21
rect 656 -71 672 -37
rect 840 -71 856 -37
rect 656 -109 856 -71
rect -856 -1147 -656 -1109
rect -856 -1181 -840 -1147
rect -672 -1181 -656 -1147
rect -856 -1197 -656 -1181
rect -478 -1147 -278 -1109
rect -478 -1181 -462 -1147
rect -294 -1181 -278 -1147
rect -478 -1197 -278 -1181
rect -100 -1147 100 -1109
rect -100 -1181 -84 -1147
rect 84 -1181 100 -1147
rect -100 -1197 100 -1181
rect 278 -1147 478 -1109
rect 278 -1181 294 -1147
rect 462 -1181 478 -1147
rect 278 -1197 478 -1181
rect 656 -1147 856 -1109
rect 656 -1181 672 -1147
rect 840 -1181 856 -1147
rect 656 -1197 856 -1181
rect -856 -1255 -656 -1239
rect -856 -1289 -840 -1255
rect -672 -1289 -656 -1255
rect -856 -1327 -656 -1289
rect -478 -1255 -278 -1239
rect -478 -1289 -462 -1255
rect -294 -1289 -278 -1255
rect -478 -1327 -278 -1289
rect -100 -1255 100 -1239
rect -100 -1289 -84 -1255
rect 84 -1289 100 -1255
rect -100 -1327 100 -1289
rect 278 -1255 478 -1239
rect 278 -1289 294 -1255
rect 462 -1289 478 -1255
rect 278 -1327 478 -1289
rect 656 -1255 856 -1239
rect 656 -1289 672 -1255
rect 840 -1289 856 -1255
rect 656 -1327 856 -1289
rect -856 -2365 -656 -2327
rect -856 -2399 -840 -2365
rect -672 -2399 -656 -2365
rect -856 -2415 -656 -2399
rect -478 -2365 -278 -2327
rect -478 -2399 -462 -2365
rect -294 -2399 -278 -2365
rect -478 -2415 -278 -2399
rect -100 -2365 100 -2327
rect -100 -2399 -84 -2365
rect 84 -2399 100 -2365
rect -100 -2415 100 -2399
rect 278 -2365 478 -2327
rect 278 -2399 294 -2365
rect 462 -2399 478 -2365
rect 278 -2415 478 -2399
rect 656 -2365 856 -2327
rect 656 -2399 672 -2365
rect 840 -2399 856 -2365
rect 656 -2415 856 -2399
<< polycont >>
rect -840 2365 -672 2399
rect -462 2365 -294 2399
rect -84 2365 84 2399
rect 294 2365 462 2399
rect 672 2365 840 2399
rect -840 1255 -672 1289
rect -462 1255 -294 1289
rect -84 1255 84 1289
rect 294 1255 462 1289
rect 672 1255 840 1289
rect -840 1147 -672 1181
rect -462 1147 -294 1181
rect -84 1147 84 1181
rect 294 1147 462 1181
rect 672 1147 840 1181
rect -840 37 -672 71
rect -462 37 -294 71
rect -84 37 84 71
rect 294 37 462 71
rect 672 37 840 71
rect -840 -71 -672 -37
rect -462 -71 -294 -37
rect -84 -71 84 -37
rect 294 -71 462 -37
rect 672 -71 840 -37
rect -840 -1181 -672 -1147
rect -462 -1181 -294 -1147
rect -84 -1181 84 -1147
rect 294 -1181 462 -1147
rect 672 -1181 840 -1147
rect -840 -1289 -672 -1255
rect -462 -1289 -294 -1255
rect -84 -1289 84 -1255
rect 294 -1289 462 -1255
rect 672 -1289 840 -1255
rect -840 -2399 -672 -2365
rect -462 -2399 -294 -2365
rect -84 -2399 84 -2365
rect 294 -2399 462 -2365
rect 672 -2399 840 -2365
<< locali >>
rect -1036 2503 -940 2537
rect 940 2503 1036 2537
rect -1036 2441 -1002 2503
rect 1002 2441 1036 2503
rect -856 2365 -840 2399
rect -672 2365 -656 2399
rect -478 2365 -462 2399
rect -294 2365 -278 2399
rect -100 2365 -84 2399
rect 84 2365 100 2399
rect 278 2365 294 2399
rect 462 2365 478 2399
rect 656 2365 672 2399
rect 840 2365 856 2399
rect -902 2315 -868 2331
rect -902 1323 -868 1339
rect -644 2315 -610 2331
rect -644 1323 -610 1339
rect -524 2315 -490 2331
rect -524 1323 -490 1339
rect -266 2315 -232 2331
rect -266 1323 -232 1339
rect -146 2315 -112 2331
rect -146 1323 -112 1339
rect 112 2315 146 2331
rect 112 1323 146 1339
rect 232 2315 266 2331
rect 232 1323 266 1339
rect 490 2315 524 2331
rect 490 1323 524 1339
rect 610 2315 644 2331
rect 610 1323 644 1339
rect 868 2315 902 2331
rect 868 1323 902 1339
rect -856 1255 -840 1289
rect -672 1255 -656 1289
rect -478 1255 -462 1289
rect -294 1255 -278 1289
rect -100 1255 -84 1289
rect 84 1255 100 1289
rect 278 1255 294 1289
rect 462 1255 478 1289
rect 656 1255 672 1289
rect 840 1255 856 1289
rect -856 1147 -840 1181
rect -672 1147 -656 1181
rect -478 1147 -462 1181
rect -294 1147 -278 1181
rect -100 1147 -84 1181
rect 84 1147 100 1181
rect 278 1147 294 1181
rect 462 1147 478 1181
rect 656 1147 672 1181
rect 840 1147 856 1181
rect -902 1097 -868 1113
rect -902 105 -868 121
rect -644 1097 -610 1113
rect -644 105 -610 121
rect -524 1097 -490 1113
rect -524 105 -490 121
rect -266 1097 -232 1113
rect -266 105 -232 121
rect -146 1097 -112 1113
rect -146 105 -112 121
rect 112 1097 146 1113
rect 112 105 146 121
rect 232 1097 266 1113
rect 232 105 266 121
rect 490 1097 524 1113
rect 490 105 524 121
rect 610 1097 644 1113
rect 610 105 644 121
rect 868 1097 902 1113
rect 868 105 902 121
rect -856 37 -840 71
rect -672 37 -656 71
rect -478 37 -462 71
rect -294 37 -278 71
rect -100 37 -84 71
rect 84 37 100 71
rect 278 37 294 71
rect 462 37 478 71
rect 656 37 672 71
rect 840 37 856 71
rect -856 -71 -840 -37
rect -672 -71 -656 -37
rect -478 -71 -462 -37
rect -294 -71 -278 -37
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect 278 -71 294 -37
rect 462 -71 478 -37
rect 656 -71 672 -37
rect 840 -71 856 -37
rect -902 -121 -868 -105
rect -902 -1113 -868 -1097
rect -644 -121 -610 -105
rect -644 -1113 -610 -1097
rect -524 -121 -490 -105
rect -524 -1113 -490 -1097
rect -266 -121 -232 -105
rect -266 -1113 -232 -1097
rect -146 -121 -112 -105
rect -146 -1113 -112 -1097
rect 112 -121 146 -105
rect 112 -1113 146 -1097
rect 232 -121 266 -105
rect 232 -1113 266 -1097
rect 490 -121 524 -105
rect 490 -1113 524 -1097
rect 610 -121 644 -105
rect 610 -1113 644 -1097
rect 868 -121 902 -105
rect 868 -1113 902 -1097
rect -856 -1181 -840 -1147
rect -672 -1181 -656 -1147
rect -478 -1181 -462 -1147
rect -294 -1181 -278 -1147
rect -100 -1181 -84 -1147
rect 84 -1181 100 -1147
rect 278 -1181 294 -1147
rect 462 -1181 478 -1147
rect 656 -1181 672 -1147
rect 840 -1181 856 -1147
rect -856 -1289 -840 -1255
rect -672 -1289 -656 -1255
rect -478 -1289 -462 -1255
rect -294 -1289 -278 -1255
rect -100 -1289 -84 -1255
rect 84 -1289 100 -1255
rect 278 -1289 294 -1255
rect 462 -1289 478 -1255
rect 656 -1289 672 -1255
rect 840 -1289 856 -1255
rect -902 -1339 -868 -1323
rect -902 -2331 -868 -2315
rect -644 -1339 -610 -1323
rect -644 -2331 -610 -2315
rect -524 -1339 -490 -1323
rect -524 -2331 -490 -2315
rect -266 -1339 -232 -1323
rect -266 -2331 -232 -2315
rect -146 -1339 -112 -1323
rect -146 -2331 -112 -2315
rect 112 -1339 146 -1323
rect 112 -2331 146 -2315
rect 232 -1339 266 -1323
rect 232 -2331 266 -2315
rect 490 -1339 524 -1323
rect 490 -2331 524 -2315
rect 610 -1339 644 -1323
rect 610 -2331 644 -2315
rect 868 -1339 902 -1323
rect 868 -2331 902 -2315
rect -856 -2399 -840 -2365
rect -672 -2399 -656 -2365
rect -478 -2399 -462 -2365
rect -294 -2399 -278 -2365
rect -100 -2399 -84 -2365
rect 84 -2399 100 -2365
rect 278 -2399 294 -2365
rect 462 -2399 478 -2365
rect 656 -2399 672 -2365
rect 840 -2399 856 -2365
rect -1036 -2503 -1002 -2441
rect 1002 -2503 1036 -2441
rect -1036 -2537 -940 -2503
rect 940 -2537 1036 -2503
<< viali >>
rect -840 2365 -672 2399
rect -462 2365 -294 2399
rect -84 2365 84 2399
rect 294 2365 462 2399
rect 672 2365 840 2399
rect -902 1339 -868 2315
rect -644 1339 -610 2315
rect -524 1339 -490 2315
rect -266 1339 -232 2315
rect -146 1339 -112 2315
rect 112 1339 146 2315
rect 232 1339 266 2315
rect 490 1339 524 2315
rect 610 1339 644 2315
rect 868 1339 902 2315
rect -840 1255 -672 1289
rect -462 1255 -294 1289
rect -84 1255 84 1289
rect 294 1255 462 1289
rect 672 1255 840 1289
rect -840 1147 -672 1181
rect -462 1147 -294 1181
rect -84 1147 84 1181
rect 294 1147 462 1181
rect 672 1147 840 1181
rect -902 121 -868 1097
rect -644 121 -610 1097
rect -524 121 -490 1097
rect -266 121 -232 1097
rect -146 121 -112 1097
rect 112 121 146 1097
rect 232 121 266 1097
rect 490 121 524 1097
rect 610 121 644 1097
rect 868 121 902 1097
rect -840 37 -672 71
rect -462 37 -294 71
rect -84 37 84 71
rect 294 37 462 71
rect 672 37 840 71
rect -840 -71 -672 -37
rect -462 -71 -294 -37
rect -84 -71 84 -37
rect 294 -71 462 -37
rect 672 -71 840 -37
rect -902 -1097 -868 -121
rect -644 -1097 -610 -121
rect -524 -1097 -490 -121
rect -266 -1097 -232 -121
rect -146 -1097 -112 -121
rect 112 -1097 146 -121
rect 232 -1097 266 -121
rect 490 -1097 524 -121
rect 610 -1097 644 -121
rect 868 -1097 902 -121
rect -840 -1181 -672 -1147
rect -462 -1181 -294 -1147
rect -84 -1181 84 -1147
rect 294 -1181 462 -1147
rect 672 -1181 840 -1147
rect -840 -1289 -672 -1255
rect -462 -1289 -294 -1255
rect -84 -1289 84 -1255
rect 294 -1289 462 -1255
rect 672 -1289 840 -1255
rect -902 -2315 -868 -1339
rect -644 -2315 -610 -1339
rect -524 -2315 -490 -1339
rect -266 -2315 -232 -1339
rect -146 -2315 -112 -1339
rect 112 -2315 146 -1339
rect 232 -2315 266 -1339
rect 490 -2315 524 -1339
rect 610 -2315 644 -1339
rect 868 -2315 902 -1339
rect -840 -2399 -672 -2365
rect -462 -2399 -294 -2365
rect -84 -2399 84 -2365
rect 294 -2399 462 -2365
rect 672 -2399 840 -2365
<< metal1 >>
rect -852 2399 -660 2405
rect -852 2365 -840 2399
rect -672 2365 -660 2399
rect -852 2359 -660 2365
rect -474 2399 -282 2405
rect -474 2365 -462 2399
rect -294 2365 -282 2399
rect -474 2359 -282 2365
rect -96 2399 96 2405
rect -96 2365 -84 2399
rect 84 2365 96 2399
rect -96 2359 96 2365
rect 282 2399 474 2405
rect 282 2365 294 2399
rect 462 2365 474 2399
rect 282 2359 474 2365
rect 660 2399 852 2405
rect 660 2365 672 2399
rect 840 2365 852 2399
rect 660 2359 852 2365
rect -908 2315 -862 2327
rect -908 1339 -902 2315
rect -868 1339 -862 2315
rect -908 1327 -862 1339
rect -650 2315 -604 2327
rect -650 1339 -644 2315
rect -610 1339 -604 2315
rect -650 1327 -604 1339
rect -530 2315 -484 2327
rect -530 1339 -524 2315
rect -490 1339 -484 2315
rect -530 1327 -484 1339
rect -272 2315 -226 2327
rect -272 1339 -266 2315
rect -232 1339 -226 2315
rect -272 1327 -226 1339
rect -152 2315 -106 2327
rect -152 1339 -146 2315
rect -112 1339 -106 2315
rect -152 1327 -106 1339
rect 106 2315 152 2327
rect 106 1339 112 2315
rect 146 1339 152 2315
rect 106 1327 152 1339
rect 226 2315 272 2327
rect 226 1339 232 2315
rect 266 1339 272 2315
rect 226 1327 272 1339
rect 484 2315 530 2327
rect 484 1339 490 2315
rect 524 1339 530 2315
rect 484 1327 530 1339
rect 604 2315 650 2327
rect 604 1339 610 2315
rect 644 1339 650 2315
rect 604 1327 650 1339
rect 862 2315 908 2327
rect 862 1339 868 2315
rect 902 1339 908 2315
rect 862 1327 908 1339
rect -852 1289 -660 1295
rect -852 1255 -840 1289
rect -672 1255 -660 1289
rect -852 1249 -660 1255
rect -474 1289 -282 1295
rect -474 1255 -462 1289
rect -294 1255 -282 1289
rect -474 1249 -282 1255
rect -96 1289 96 1295
rect -96 1255 -84 1289
rect 84 1255 96 1289
rect -96 1249 96 1255
rect 282 1289 474 1295
rect 282 1255 294 1289
rect 462 1255 474 1289
rect 282 1249 474 1255
rect 660 1289 852 1295
rect 660 1255 672 1289
rect 840 1255 852 1289
rect 660 1249 852 1255
rect -852 1181 -660 1187
rect -852 1147 -840 1181
rect -672 1147 -660 1181
rect -852 1141 -660 1147
rect -474 1181 -282 1187
rect -474 1147 -462 1181
rect -294 1147 -282 1181
rect -474 1141 -282 1147
rect -96 1181 96 1187
rect -96 1147 -84 1181
rect 84 1147 96 1181
rect -96 1141 96 1147
rect 282 1181 474 1187
rect 282 1147 294 1181
rect 462 1147 474 1181
rect 282 1141 474 1147
rect 660 1181 852 1187
rect 660 1147 672 1181
rect 840 1147 852 1181
rect 660 1141 852 1147
rect -908 1097 -862 1109
rect -908 121 -902 1097
rect -868 121 -862 1097
rect -908 109 -862 121
rect -650 1097 -604 1109
rect -650 121 -644 1097
rect -610 121 -604 1097
rect -650 109 -604 121
rect -530 1097 -484 1109
rect -530 121 -524 1097
rect -490 121 -484 1097
rect -530 109 -484 121
rect -272 1097 -226 1109
rect -272 121 -266 1097
rect -232 121 -226 1097
rect -272 109 -226 121
rect -152 1097 -106 1109
rect -152 121 -146 1097
rect -112 121 -106 1097
rect -152 109 -106 121
rect 106 1097 152 1109
rect 106 121 112 1097
rect 146 121 152 1097
rect 106 109 152 121
rect 226 1097 272 1109
rect 226 121 232 1097
rect 266 121 272 1097
rect 226 109 272 121
rect 484 1097 530 1109
rect 484 121 490 1097
rect 524 121 530 1097
rect 484 109 530 121
rect 604 1097 650 1109
rect 604 121 610 1097
rect 644 121 650 1097
rect 604 109 650 121
rect 862 1097 908 1109
rect 862 121 868 1097
rect 902 121 908 1097
rect 862 109 908 121
rect -852 71 -660 77
rect -852 37 -840 71
rect -672 37 -660 71
rect -852 31 -660 37
rect -474 71 -282 77
rect -474 37 -462 71
rect -294 37 -282 71
rect -474 31 -282 37
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect 282 71 474 77
rect 282 37 294 71
rect 462 37 474 71
rect 282 31 474 37
rect 660 71 852 77
rect 660 37 672 71
rect 840 37 852 71
rect 660 31 852 37
rect -852 -37 -660 -31
rect -852 -71 -840 -37
rect -672 -71 -660 -37
rect -852 -77 -660 -71
rect -474 -37 -282 -31
rect -474 -71 -462 -37
rect -294 -71 -282 -37
rect -474 -77 -282 -71
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect 282 -37 474 -31
rect 282 -71 294 -37
rect 462 -71 474 -37
rect 282 -77 474 -71
rect 660 -37 852 -31
rect 660 -71 672 -37
rect 840 -71 852 -37
rect 660 -77 852 -71
rect -908 -121 -862 -109
rect -908 -1097 -902 -121
rect -868 -1097 -862 -121
rect -908 -1109 -862 -1097
rect -650 -121 -604 -109
rect -650 -1097 -644 -121
rect -610 -1097 -604 -121
rect -650 -1109 -604 -1097
rect -530 -121 -484 -109
rect -530 -1097 -524 -121
rect -490 -1097 -484 -121
rect -530 -1109 -484 -1097
rect -272 -121 -226 -109
rect -272 -1097 -266 -121
rect -232 -1097 -226 -121
rect -272 -1109 -226 -1097
rect -152 -121 -106 -109
rect -152 -1097 -146 -121
rect -112 -1097 -106 -121
rect -152 -1109 -106 -1097
rect 106 -121 152 -109
rect 106 -1097 112 -121
rect 146 -1097 152 -121
rect 106 -1109 152 -1097
rect 226 -121 272 -109
rect 226 -1097 232 -121
rect 266 -1097 272 -121
rect 226 -1109 272 -1097
rect 484 -121 530 -109
rect 484 -1097 490 -121
rect 524 -1097 530 -121
rect 484 -1109 530 -1097
rect 604 -121 650 -109
rect 604 -1097 610 -121
rect 644 -1097 650 -121
rect 604 -1109 650 -1097
rect 862 -121 908 -109
rect 862 -1097 868 -121
rect 902 -1097 908 -121
rect 862 -1109 908 -1097
rect -852 -1147 -660 -1141
rect -852 -1181 -840 -1147
rect -672 -1181 -660 -1147
rect -852 -1187 -660 -1181
rect -474 -1147 -282 -1141
rect -474 -1181 -462 -1147
rect -294 -1181 -282 -1147
rect -474 -1187 -282 -1181
rect -96 -1147 96 -1141
rect -96 -1181 -84 -1147
rect 84 -1181 96 -1147
rect -96 -1187 96 -1181
rect 282 -1147 474 -1141
rect 282 -1181 294 -1147
rect 462 -1181 474 -1147
rect 282 -1187 474 -1181
rect 660 -1147 852 -1141
rect 660 -1181 672 -1147
rect 840 -1181 852 -1147
rect 660 -1187 852 -1181
rect -852 -1255 -660 -1249
rect -852 -1289 -840 -1255
rect -672 -1289 -660 -1255
rect -852 -1295 -660 -1289
rect -474 -1255 -282 -1249
rect -474 -1289 -462 -1255
rect -294 -1289 -282 -1255
rect -474 -1295 -282 -1289
rect -96 -1255 96 -1249
rect -96 -1289 -84 -1255
rect 84 -1289 96 -1255
rect -96 -1295 96 -1289
rect 282 -1255 474 -1249
rect 282 -1289 294 -1255
rect 462 -1289 474 -1255
rect 282 -1295 474 -1289
rect 660 -1255 852 -1249
rect 660 -1289 672 -1255
rect 840 -1289 852 -1255
rect 660 -1295 852 -1289
rect -908 -1339 -862 -1327
rect -908 -2315 -902 -1339
rect -868 -2315 -862 -1339
rect -908 -2327 -862 -2315
rect -650 -1339 -604 -1327
rect -650 -2315 -644 -1339
rect -610 -2315 -604 -1339
rect -650 -2327 -604 -2315
rect -530 -1339 -484 -1327
rect -530 -2315 -524 -1339
rect -490 -2315 -484 -1339
rect -530 -2327 -484 -2315
rect -272 -1339 -226 -1327
rect -272 -2315 -266 -1339
rect -232 -2315 -226 -1339
rect -272 -2327 -226 -2315
rect -152 -1339 -106 -1327
rect -152 -2315 -146 -1339
rect -112 -2315 -106 -1339
rect -152 -2327 -106 -2315
rect 106 -1339 152 -1327
rect 106 -2315 112 -1339
rect 146 -2315 152 -1339
rect 106 -2327 152 -2315
rect 226 -1339 272 -1327
rect 226 -2315 232 -1339
rect 266 -2315 272 -1339
rect 226 -2327 272 -2315
rect 484 -1339 530 -1327
rect 484 -2315 490 -1339
rect 524 -2315 530 -1339
rect 484 -2327 530 -2315
rect 604 -1339 650 -1327
rect 604 -2315 610 -1339
rect 644 -2315 650 -1339
rect 604 -2327 650 -2315
rect 862 -1339 908 -1327
rect 862 -2315 868 -1339
rect 902 -2315 908 -1339
rect 862 -2327 908 -2315
rect -852 -2365 -660 -2359
rect -852 -2399 -840 -2365
rect -672 -2399 -660 -2365
rect -852 -2405 -660 -2399
rect -474 -2365 -282 -2359
rect -474 -2399 -462 -2365
rect -294 -2399 -282 -2365
rect -474 -2405 -282 -2399
rect -96 -2365 96 -2359
rect -96 -2399 -84 -2365
rect 84 -2399 96 -2365
rect -96 -2405 96 -2399
rect 282 -2365 474 -2359
rect 282 -2399 294 -2365
rect 462 -2399 474 -2365
rect 282 -2405 474 -2399
rect 660 -2365 852 -2359
rect 660 -2399 672 -2365
rect 840 -2399 852 -2365
rect 660 -2405 852 -2399
<< properties >>
string FIXED_BBOX -1019 -2520 1019 2520
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 1.0 m 4 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
