magic
tech sky130A
magscale 1 2
timestamp 1729620069
<< pwell >>
rect -328 -121949 328 121949
<< mvnmos >>
rect -100 120691 100 121691
rect -100 119473 100 120473
rect -100 118255 100 119255
rect -100 117037 100 118037
rect -100 115819 100 116819
rect -100 114601 100 115601
rect -100 113383 100 114383
rect -100 112165 100 113165
rect -100 110947 100 111947
rect -100 109729 100 110729
rect -100 108511 100 109511
rect -100 107293 100 108293
rect -100 106075 100 107075
rect -100 104857 100 105857
rect -100 103639 100 104639
rect -100 102421 100 103421
rect -100 101203 100 102203
rect -100 99985 100 100985
rect -100 98767 100 99767
rect -100 97549 100 98549
rect -100 96331 100 97331
rect -100 95113 100 96113
rect -100 93895 100 94895
rect -100 92677 100 93677
rect -100 91459 100 92459
rect -100 90241 100 91241
rect -100 89023 100 90023
rect -100 87805 100 88805
rect -100 86587 100 87587
rect -100 85369 100 86369
rect -100 84151 100 85151
rect -100 82933 100 83933
rect -100 81715 100 82715
rect -100 80497 100 81497
rect -100 79279 100 80279
rect -100 78061 100 79061
rect -100 76843 100 77843
rect -100 75625 100 76625
rect -100 74407 100 75407
rect -100 73189 100 74189
rect -100 71971 100 72971
rect -100 70753 100 71753
rect -100 69535 100 70535
rect -100 68317 100 69317
rect -100 67099 100 68099
rect -100 65881 100 66881
rect -100 64663 100 65663
rect -100 63445 100 64445
rect -100 62227 100 63227
rect -100 61009 100 62009
rect -100 59791 100 60791
rect -100 58573 100 59573
rect -100 57355 100 58355
rect -100 56137 100 57137
rect -100 54919 100 55919
rect -100 53701 100 54701
rect -100 52483 100 53483
rect -100 51265 100 52265
rect -100 50047 100 51047
rect -100 48829 100 49829
rect -100 47611 100 48611
rect -100 46393 100 47393
rect -100 45175 100 46175
rect -100 43957 100 44957
rect -100 42739 100 43739
rect -100 41521 100 42521
rect -100 40303 100 41303
rect -100 39085 100 40085
rect -100 37867 100 38867
rect -100 36649 100 37649
rect -100 35431 100 36431
rect -100 34213 100 35213
rect -100 32995 100 33995
rect -100 31777 100 32777
rect -100 30559 100 31559
rect -100 29341 100 30341
rect -100 28123 100 29123
rect -100 26905 100 27905
rect -100 25687 100 26687
rect -100 24469 100 25469
rect -100 23251 100 24251
rect -100 22033 100 23033
rect -100 20815 100 21815
rect -100 19597 100 20597
rect -100 18379 100 19379
rect -100 17161 100 18161
rect -100 15943 100 16943
rect -100 14725 100 15725
rect -100 13507 100 14507
rect -100 12289 100 13289
rect -100 11071 100 12071
rect -100 9853 100 10853
rect -100 8635 100 9635
rect -100 7417 100 8417
rect -100 6199 100 7199
rect -100 4981 100 5981
rect -100 3763 100 4763
rect -100 2545 100 3545
rect -100 1327 100 2327
rect -100 109 100 1109
rect -100 -1109 100 -109
rect -100 -2327 100 -1327
rect -100 -3545 100 -2545
rect -100 -4763 100 -3763
rect -100 -5981 100 -4981
rect -100 -7199 100 -6199
rect -100 -8417 100 -7417
rect -100 -9635 100 -8635
rect -100 -10853 100 -9853
rect -100 -12071 100 -11071
rect -100 -13289 100 -12289
rect -100 -14507 100 -13507
rect -100 -15725 100 -14725
rect -100 -16943 100 -15943
rect -100 -18161 100 -17161
rect -100 -19379 100 -18379
rect -100 -20597 100 -19597
rect -100 -21815 100 -20815
rect -100 -23033 100 -22033
rect -100 -24251 100 -23251
rect -100 -25469 100 -24469
rect -100 -26687 100 -25687
rect -100 -27905 100 -26905
rect -100 -29123 100 -28123
rect -100 -30341 100 -29341
rect -100 -31559 100 -30559
rect -100 -32777 100 -31777
rect -100 -33995 100 -32995
rect -100 -35213 100 -34213
rect -100 -36431 100 -35431
rect -100 -37649 100 -36649
rect -100 -38867 100 -37867
rect -100 -40085 100 -39085
rect -100 -41303 100 -40303
rect -100 -42521 100 -41521
rect -100 -43739 100 -42739
rect -100 -44957 100 -43957
rect -100 -46175 100 -45175
rect -100 -47393 100 -46393
rect -100 -48611 100 -47611
rect -100 -49829 100 -48829
rect -100 -51047 100 -50047
rect -100 -52265 100 -51265
rect -100 -53483 100 -52483
rect -100 -54701 100 -53701
rect -100 -55919 100 -54919
rect -100 -57137 100 -56137
rect -100 -58355 100 -57355
rect -100 -59573 100 -58573
rect -100 -60791 100 -59791
rect -100 -62009 100 -61009
rect -100 -63227 100 -62227
rect -100 -64445 100 -63445
rect -100 -65663 100 -64663
rect -100 -66881 100 -65881
rect -100 -68099 100 -67099
rect -100 -69317 100 -68317
rect -100 -70535 100 -69535
rect -100 -71753 100 -70753
rect -100 -72971 100 -71971
rect -100 -74189 100 -73189
rect -100 -75407 100 -74407
rect -100 -76625 100 -75625
rect -100 -77843 100 -76843
rect -100 -79061 100 -78061
rect -100 -80279 100 -79279
rect -100 -81497 100 -80497
rect -100 -82715 100 -81715
rect -100 -83933 100 -82933
rect -100 -85151 100 -84151
rect -100 -86369 100 -85369
rect -100 -87587 100 -86587
rect -100 -88805 100 -87805
rect -100 -90023 100 -89023
rect -100 -91241 100 -90241
rect -100 -92459 100 -91459
rect -100 -93677 100 -92677
rect -100 -94895 100 -93895
rect -100 -96113 100 -95113
rect -100 -97331 100 -96331
rect -100 -98549 100 -97549
rect -100 -99767 100 -98767
rect -100 -100985 100 -99985
rect -100 -102203 100 -101203
rect -100 -103421 100 -102421
rect -100 -104639 100 -103639
rect -100 -105857 100 -104857
rect -100 -107075 100 -106075
rect -100 -108293 100 -107293
rect -100 -109511 100 -108511
rect -100 -110729 100 -109729
rect -100 -111947 100 -110947
rect -100 -113165 100 -112165
rect -100 -114383 100 -113383
rect -100 -115601 100 -114601
rect -100 -116819 100 -115819
rect -100 -118037 100 -117037
rect -100 -119255 100 -118255
rect -100 -120473 100 -119473
rect -100 -121691 100 -120691
<< mvndiff >>
rect -158 121679 -100 121691
rect -158 120703 -146 121679
rect -112 120703 -100 121679
rect -158 120691 -100 120703
rect 100 121679 158 121691
rect 100 120703 112 121679
rect 146 120703 158 121679
rect 100 120691 158 120703
rect -158 120461 -100 120473
rect -158 119485 -146 120461
rect -112 119485 -100 120461
rect -158 119473 -100 119485
rect 100 120461 158 120473
rect 100 119485 112 120461
rect 146 119485 158 120461
rect 100 119473 158 119485
rect -158 119243 -100 119255
rect -158 118267 -146 119243
rect -112 118267 -100 119243
rect -158 118255 -100 118267
rect 100 119243 158 119255
rect 100 118267 112 119243
rect 146 118267 158 119243
rect 100 118255 158 118267
rect -158 118025 -100 118037
rect -158 117049 -146 118025
rect -112 117049 -100 118025
rect -158 117037 -100 117049
rect 100 118025 158 118037
rect 100 117049 112 118025
rect 146 117049 158 118025
rect 100 117037 158 117049
rect -158 116807 -100 116819
rect -158 115831 -146 116807
rect -112 115831 -100 116807
rect -158 115819 -100 115831
rect 100 116807 158 116819
rect 100 115831 112 116807
rect 146 115831 158 116807
rect 100 115819 158 115831
rect -158 115589 -100 115601
rect -158 114613 -146 115589
rect -112 114613 -100 115589
rect -158 114601 -100 114613
rect 100 115589 158 115601
rect 100 114613 112 115589
rect 146 114613 158 115589
rect 100 114601 158 114613
rect -158 114371 -100 114383
rect -158 113395 -146 114371
rect -112 113395 -100 114371
rect -158 113383 -100 113395
rect 100 114371 158 114383
rect 100 113395 112 114371
rect 146 113395 158 114371
rect 100 113383 158 113395
rect -158 113153 -100 113165
rect -158 112177 -146 113153
rect -112 112177 -100 113153
rect -158 112165 -100 112177
rect 100 113153 158 113165
rect 100 112177 112 113153
rect 146 112177 158 113153
rect 100 112165 158 112177
rect -158 111935 -100 111947
rect -158 110959 -146 111935
rect -112 110959 -100 111935
rect -158 110947 -100 110959
rect 100 111935 158 111947
rect 100 110959 112 111935
rect 146 110959 158 111935
rect 100 110947 158 110959
rect -158 110717 -100 110729
rect -158 109741 -146 110717
rect -112 109741 -100 110717
rect -158 109729 -100 109741
rect 100 110717 158 110729
rect 100 109741 112 110717
rect 146 109741 158 110717
rect 100 109729 158 109741
rect -158 109499 -100 109511
rect -158 108523 -146 109499
rect -112 108523 -100 109499
rect -158 108511 -100 108523
rect 100 109499 158 109511
rect 100 108523 112 109499
rect 146 108523 158 109499
rect 100 108511 158 108523
rect -158 108281 -100 108293
rect -158 107305 -146 108281
rect -112 107305 -100 108281
rect -158 107293 -100 107305
rect 100 108281 158 108293
rect 100 107305 112 108281
rect 146 107305 158 108281
rect 100 107293 158 107305
rect -158 107063 -100 107075
rect -158 106087 -146 107063
rect -112 106087 -100 107063
rect -158 106075 -100 106087
rect 100 107063 158 107075
rect 100 106087 112 107063
rect 146 106087 158 107063
rect 100 106075 158 106087
rect -158 105845 -100 105857
rect -158 104869 -146 105845
rect -112 104869 -100 105845
rect -158 104857 -100 104869
rect 100 105845 158 105857
rect 100 104869 112 105845
rect 146 104869 158 105845
rect 100 104857 158 104869
rect -158 104627 -100 104639
rect -158 103651 -146 104627
rect -112 103651 -100 104627
rect -158 103639 -100 103651
rect 100 104627 158 104639
rect 100 103651 112 104627
rect 146 103651 158 104627
rect 100 103639 158 103651
rect -158 103409 -100 103421
rect -158 102433 -146 103409
rect -112 102433 -100 103409
rect -158 102421 -100 102433
rect 100 103409 158 103421
rect 100 102433 112 103409
rect 146 102433 158 103409
rect 100 102421 158 102433
rect -158 102191 -100 102203
rect -158 101215 -146 102191
rect -112 101215 -100 102191
rect -158 101203 -100 101215
rect 100 102191 158 102203
rect 100 101215 112 102191
rect 146 101215 158 102191
rect 100 101203 158 101215
rect -158 100973 -100 100985
rect -158 99997 -146 100973
rect -112 99997 -100 100973
rect -158 99985 -100 99997
rect 100 100973 158 100985
rect 100 99997 112 100973
rect 146 99997 158 100973
rect 100 99985 158 99997
rect -158 99755 -100 99767
rect -158 98779 -146 99755
rect -112 98779 -100 99755
rect -158 98767 -100 98779
rect 100 99755 158 99767
rect 100 98779 112 99755
rect 146 98779 158 99755
rect 100 98767 158 98779
rect -158 98537 -100 98549
rect -158 97561 -146 98537
rect -112 97561 -100 98537
rect -158 97549 -100 97561
rect 100 98537 158 98549
rect 100 97561 112 98537
rect 146 97561 158 98537
rect 100 97549 158 97561
rect -158 97319 -100 97331
rect -158 96343 -146 97319
rect -112 96343 -100 97319
rect -158 96331 -100 96343
rect 100 97319 158 97331
rect 100 96343 112 97319
rect 146 96343 158 97319
rect 100 96331 158 96343
rect -158 96101 -100 96113
rect -158 95125 -146 96101
rect -112 95125 -100 96101
rect -158 95113 -100 95125
rect 100 96101 158 96113
rect 100 95125 112 96101
rect 146 95125 158 96101
rect 100 95113 158 95125
rect -158 94883 -100 94895
rect -158 93907 -146 94883
rect -112 93907 -100 94883
rect -158 93895 -100 93907
rect 100 94883 158 94895
rect 100 93907 112 94883
rect 146 93907 158 94883
rect 100 93895 158 93907
rect -158 93665 -100 93677
rect -158 92689 -146 93665
rect -112 92689 -100 93665
rect -158 92677 -100 92689
rect 100 93665 158 93677
rect 100 92689 112 93665
rect 146 92689 158 93665
rect 100 92677 158 92689
rect -158 92447 -100 92459
rect -158 91471 -146 92447
rect -112 91471 -100 92447
rect -158 91459 -100 91471
rect 100 92447 158 92459
rect 100 91471 112 92447
rect 146 91471 158 92447
rect 100 91459 158 91471
rect -158 91229 -100 91241
rect -158 90253 -146 91229
rect -112 90253 -100 91229
rect -158 90241 -100 90253
rect 100 91229 158 91241
rect 100 90253 112 91229
rect 146 90253 158 91229
rect 100 90241 158 90253
rect -158 90011 -100 90023
rect -158 89035 -146 90011
rect -112 89035 -100 90011
rect -158 89023 -100 89035
rect 100 90011 158 90023
rect 100 89035 112 90011
rect 146 89035 158 90011
rect 100 89023 158 89035
rect -158 88793 -100 88805
rect -158 87817 -146 88793
rect -112 87817 -100 88793
rect -158 87805 -100 87817
rect 100 88793 158 88805
rect 100 87817 112 88793
rect 146 87817 158 88793
rect 100 87805 158 87817
rect -158 87575 -100 87587
rect -158 86599 -146 87575
rect -112 86599 -100 87575
rect -158 86587 -100 86599
rect 100 87575 158 87587
rect 100 86599 112 87575
rect 146 86599 158 87575
rect 100 86587 158 86599
rect -158 86357 -100 86369
rect -158 85381 -146 86357
rect -112 85381 -100 86357
rect -158 85369 -100 85381
rect 100 86357 158 86369
rect 100 85381 112 86357
rect 146 85381 158 86357
rect 100 85369 158 85381
rect -158 85139 -100 85151
rect -158 84163 -146 85139
rect -112 84163 -100 85139
rect -158 84151 -100 84163
rect 100 85139 158 85151
rect 100 84163 112 85139
rect 146 84163 158 85139
rect 100 84151 158 84163
rect -158 83921 -100 83933
rect -158 82945 -146 83921
rect -112 82945 -100 83921
rect -158 82933 -100 82945
rect 100 83921 158 83933
rect 100 82945 112 83921
rect 146 82945 158 83921
rect 100 82933 158 82945
rect -158 82703 -100 82715
rect -158 81727 -146 82703
rect -112 81727 -100 82703
rect -158 81715 -100 81727
rect 100 82703 158 82715
rect 100 81727 112 82703
rect 146 81727 158 82703
rect 100 81715 158 81727
rect -158 81485 -100 81497
rect -158 80509 -146 81485
rect -112 80509 -100 81485
rect -158 80497 -100 80509
rect 100 81485 158 81497
rect 100 80509 112 81485
rect 146 80509 158 81485
rect 100 80497 158 80509
rect -158 80267 -100 80279
rect -158 79291 -146 80267
rect -112 79291 -100 80267
rect -158 79279 -100 79291
rect 100 80267 158 80279
rect 100 79291 112 80267
rect 146 79291 158 80267
rect 100 79279 158 79291
rect -158 79049 -100 79061
rect -158 78073 -146 79049
rect -112 78073 -100 79049
rect -158 78061 -100 78073
rect 100 79049 158 79061
rect 100 78073 112 79049
rect 146 78073 158 79049
rect 100 78061 158 78073
rect -158 77831 -100 77843
rect -158 76855 -146 77831
rect -112 76855 -100 77831
rect -158 76843 -100 76855
rect 100 77831 158 77843
rect 100 76855 112 77831
rect 146 76855 158 77831
rect 100 76843 158 76855
rect -158 76613 -100 76625
rect -158 75637 -146 76613
rect -112 75637 -100 76613
rect -158 75625 -100 75637
rect 100 76613 158 76625
rect 100 75637 112 76613
rect 146 75637 158 76613
rect 100 75625 158 75637
rect -158 75395 -100 75407
rect -158 74419 -146 75395
rect -112 74419 -100 75395
rect -158 74407 -100 74419
rect 100 75395 158 75407
rect 100 74419 112 75395
rect 146 74419 158 75395
rect 100 74407 158 74419
rect -158 74177 -100 74189
rect -158 73201 -146 74177
rect -112 73201 -100 74177
rect -158 73189 -100 73201
rect 100 74177 158 74189
rect 100 73201 112 74177
rect 146 73201 158 74177
rect 100 73189 158 73201
rect -158 72959 -100 72971
rect -158 71983 -146 72959
rect -112 71983 -100 72959
rect -158 71971 -100 71983
rect 100 72959 158 72971
rect 100 71983 112 72959
rect 146 71983 158 72959
rect 100 71971 158 71983
rect -158 71741 -100 71753
rect -158 70765 -146 71741
rect -112 70765 -100 71741
rect -158 70753 -100 70765
rect 100 71741 158 71753
rect 100 70765 112 71741
rect 146 70765 158 71741
rect 100 70753 158 70765
rect -158 70523 -100 70535
rect -158 69547 -146 70523
rect -112 69547 -100 70523
rect -158 69535 -100 69547
rect 100 70523 158 70535
rect 100 69547 112 70523
rect 146 69547 158 70523
rect 100 69535 158 69547
rect -158 69305 -100 69317
rect -158 68329 -146 69305
rect -112 68329 -100 69305
rect -158 68317 -100 68329
rect 100 69305 158 69317
rect 100 68329 112 69305
rect 146 68329 158 69305
rect 100 68317 158 68329
rect -158 68087 -100 68099
rect -158 67111 -146 68087
rect -112 67111 -100 68087
rect -158 67099 -100 67111
rect 100 68087 158 68099
rect 100 67111 112 68087
rect 146 67111 158 68087
rect 100 67099 158 67111
rect -158 66869 -100 66881
rect -158 65893 -146 66869
rect -112 65893 -100 66869
rect -158 65881 -100 65893
rect 100 66869 158 66881
rect 100 65893 112 66869
rect 146 65893 158 66869
rect 100 65881 158 65893
rect -158 65651 -100 65663
rect -158 64675 -146 65651
rect -112 64675 -100 65651
rect -158 64663 -100 64675
rect 100 65651 158 65663
rect 100 64675 112 65651
rect 146 64675 158 65651
rect 100 64663 158 64675
rect -158 64433 -100 64445
rect -158 63457 -146 64433
rect -112 63457 -100 64433
rect -158 63445 -100 63457
rect 100 64433 158 64445
rect 100 63457 112 64433
rect 146 63457 158 64433
rect 100 63445 158 63457
rect -158 63215 -100 63227
rect -158 62239 -146 63215
rect -112 62239 -100 63215
rect -158 62227 -100 62239
rect 100 63215 158 63227
rect 100 62239 112 63215
rect 146 62239 158 63215
rect 100 62227 158 62239
rect -158 61997 -100 62009
rect -158 61021 -146 61997
rect -112 61021 -100 61997
rect -158 61009 -100 61021
rect 100 61997 158 62009
rect 100 61021 112 61997
rect 146 61021 158 61997
rect 100 61009 158 61021
rect -158 60779 -100 60791
rect -158 59803 -146 60779
rect -112 59803 -100 60779
rect -158 59791 -100 59803
rect 100 60779 158 60791
rect 100 59803 112 60779
rect 146 59803 158 60779
rect 100 59791 158 59803
rect -158 59561 -100 59573
rect -158 58585 -146 59561
rect -112 58585 -100 59561
rect -158 58573 -100 58585
rect 100 59561 158 59573
rect 100 58585 112 59561
rect 146 58585 158 59561
rect 100 58573 158 58585
rect -158 58343 -100 58355
rect -158 57367 -146 58343
rect -112 57367 -100 58343
rect -158 57355 -100 57367
rect 100 58343 158 58355
rect 100 57367 112 58343
rect 146 57367 158 58343
rect 100 57355 158 57367
rect -158 57125 -100 57137
rect -158 56149 -146 57125
rect -112 56149 -100 57125
rect -158 56137 -100 56149
rect 100 57125 158 57137
rect 100 56149 112 57125
rect 146 56149 158 57125
rect 100 56137 158 56149
rect -158 55907 -100 55919
rect -158 54931 -146 55907
rect -112 54931 -100 55907
rect -158 54919 -100 54931
rect 100 55907 158 55919
rect 100 54931 112 55907
rect 146 54931 158 55907
rect 100 54919 158 54931
rect -158 54689 -100 54701
rect -158 53713 -146 54689
rect -112 53713 -100 54689
rect -158 53701 -100 53713
rect 100 54689 158 54701
rect 100 53713 112 54689
rect 146 53713 158 54689
rect 100 53701 158 53713
rect -158 53471 -100 53483
rect -158 52495 -146 53471
rect -112 52495 -100 53471
rect -158 52483 -100 52495
rect 100 53471 158 53483
rect 100 52495 112 53471
rect 146 52495 158 53471
rect 100 52483 158 52495
rect -158 52253 -100 52265
rect -158 51277 -146 52253
rect -112 51277 -100 52253
rect -158 51265 -100 51277
rect 100 52253 158 52265
rect 100 51277 112 52253
rect 146 51277 158 52253
rect 100 51265 158 51277
rect -158 51035 -100 51047
rect -158 50059 -146 51035
rect -112 50059 -100 51035
rect -158 50047 -100 50059
rect 100 51035 158 51047
rect 100 50059 112 51035
rect 146 50059 158 51035
rect 100 50047 158 50059
rect -158 49817 -100 49829
rect -158 48841 -146 49817
rect -112 48841 -100 49817
rect -158 48829 -100 48841
rect 100 49817 158 49829
rect 100 48841 112 49817
rect 146 48841 158 49817
rect 100 48829 158 48841
rect -158 48599 -100 48611
rect -158 47623 -146 48599
rect -112 47623 -100 48599
rect -158 47611 -100 47623
rect 100 48599 158 48611
rect 100 47623 112 48599
rect 146 47623 158 48599
rect 100 47611 158 47623
rect -158 47381 -100 47393
rect -158 46405 -146 47381
rect -112 46405 -100 47381
rect -158 46393 -100 46405
rect 100 47381 158 47393
rect 100 46405 112 47381
rect 146 46405 158 47381
rect 100 46393 158 46405
rect -158 46163 -100 46175
rect -158 45187 -146 46163
rect -112 45187 -100 46163
rect -158 45175 -100 45187
rect 100 46163 158 46175
rect 100 45187 112 46163
rect 146 45187 158 46163
rect 100 45175 158 45187
rect -158 44945 -100 44957
rect -158 43969 -146 44945
rect -112 43969 -100 44945
rect -158 43957 -100 43969
rect 100 44945 158 44957
rect 100 43969 112 44945
rect 146 43969 158 44945
rect 100 43957 158 43969
rect -158 43727 -100 43739
rect -158 42751 -146 43727
rect -112 42751 -100 43727
rect -158 42739 -100 42751
rect 100 43727 158 43739
rect 100 42751 112 43727
rect 146 42751 158 43727
rect 100 42739 158 42751
rect -158 42509 -100 42521
rect -158 41533 -146 42509
rect -112 41533 -100 42509
rect -158 41521 -100 41533
rect 100 42509 158 42521
rect 100 41533 112 42509
rect 146 41533 158 42509
rect 100 41521 158 41533
rect -158 41291 -100 41303
rect -158 40315 -146 41291
rect -112 40315 -100 41291
rect -158 40303 -100 40315
rect 100 41291 158 41303
rect 100 40315 112 41291
rect 146 40315 158 41291
rect 100 40303 158 40315
rect -158 40073 -100 40085
rect -158 39097 -146 40073
rect -112 39097 -100 40073
rect -158 39085 -100 39097
rect 100 40073 158 40085
rect 100 39097 112 40073
rect 146 39097 158 40073
rect 100 39085 158 39097
rect -158 38855 -100 38867
rect -158 37879 -146 38855
rect -112 37879 -100 38855
rect -158 37867 -100 37879
rect 100 38855 158 38867
rect 100 37879 112 38855
rect 146 37879 158 38855
rect 100 37867 158 37879
rect -158 37637 -100 37649
rect -158 36661 -146 37637
rect -112 36661 -100 37637
rect -158 36649 -100 36661
rect 100 37637 158 37649
rect 100 36661 112 37637
rect 146 36661 158 37637
rect 100 36649 158 36661
rect -158 36419 -100 36431
rect -158 35443 -146 36419
rect -112 35443 -100 36419
rect -158 35431 -100 35443
rect 100 36419 158 36431
rect 100 35443 112 36419
rect 146 35443 158 36419
rect 100 35431 158 35443
rect -158 35201 -100 35213
rect -158 34225 -146 35201
rect -112 34225 -100 35201
rect -158 34213 -100 34225
rect 100 35201 158 35213
rect 100 34225 112 35201
rect 146 34225 158 35201
rect 100 34213 158 34225
rect -158 33983 -100 33995
rect -158 33007 -146 33983
rect -112 33007 -100 33983
rect -158 32995 -100 33007
rect 100 33983 158 33995
rect 100 33007 112 33983
rect 146 33007 158 33983
rect 100 32995 158 33007
rect -158 32765 -100 32777
rect -158 31789 -146 32765
rect -112 31789 -100 32765
rect -158 31777 -100 31789
rect 100 32765 158 32777
rect 100 31789 112 32765
rect 146 31789 158 32765
rect 100 31777 158 31789
rect -158 31547 -100 31559
rect -158 30571 -146 31547
rect -112 30571 -100 31547
rect -158 30559 -100 30571
rect 100 31547 158 31559
rect 100 30571 112 31547
rect 146 30571 158 31547
rect 100 30559 158 30571
rect -158 30329 -100 30341
rect -158 29353 -146 30329
rect -112 29353 -100 30329
rect -158 29341 -100 29353
rect 100 30329 158 30341
rect 100 29353 112 30329
rect 146 29353 158 30329
rect 100 29341 158 29353
rect -158 29111 -100 29123
rect -158 28135 -146 29111
rect -112 28135 -100 29111
rect -158 28123 -100 28135
rect 100 29111 158 29123
rect 100 28135 112 29111
rect 146 28135 158 29111
rect 100 28123 158 28135
rect -158 27893 -100 27905
rect -158 26917 -146 27893
rect -112 26917 -100 27893
rect -158 26905 -100 26917
rect 100 27893 158 27905
rect 100 26917 112 27893
rect 146 26917 158 27893
rect 100 26905 158 26917
rect -158 26675 -100 26687
rect -158 25699 -146 26675
rect -112 25699 -100 26675
rect -158 25687 -100 25699
rect 100 26675 158 26687
rect 100 25699 112 26675
rect 146 25699 158 26675
rect 100 25687 158 25699
rect -158 25457 -100 25469
rect -158 24481 -146 25457
rect -112 24481 -100 25457
rect -158 24469 -100 24481
rect 100 25457 158 25469
rect 100 24481 112 25457
rect 146 24481 158 25457
rect 100 24469 158 24481
rect -158 24239 -100 24251
rect -158 23263 -146 24239
rect -112 23263 -100 24239
rect -158 23251 -100 23263
rect 100 24239 158 24251
rect 100 23263 112 24239
rect 146 23263 158 24239
rect 100 23251 158 23263
rect -158 23021 -100 23033
rect -158 22045 -146 23021
rect -112 22045 -100 23021
rect -158 22033 -100 22045
rect 100 23021 158 23033
rect 100 22045 112 23021
rect 146 22045 158 23021
rect 100 22033 158 22045
rect -158 21803 -100 21815
rect -158 20827 -146 21803
rect -112 20827 -100 21803
rect -158 20815 -100 20827
rect 100 21803 158 21815
rect 100 20827 112 21803
rect 146 20827 158 21803
rect 100 20815 158 20827
rect -158 20585 -100 20597
rect -158 19609 -146 20585
rect -112 19609 -100 20585
rect -158 19597 -100 19609
rect 100 20585 158 20597
rect 100 19609 112 20585
rect 146 19609 158 20585
rect 100 19597 158 19609
rect -158 19367 -100 19379
rect -158 18391 -146 19367
rect -112 18391 -100 19367
rect -158 18379 -100 18391
rect 100 19367 158 19379
rect 100 18391 112 19367
rect 146 18391 158 19367
rect 100 18379 158 18391
rect -158 18149 -100 18161
rect -158 17173 -146 18149
rect -112 17173 -100 18149
rect -158 17161 -100 17173
rect 100 18149 158 18161
rect 100 17173 112 18149
rect 146 17173 158 18149
rect 100 17161 158 17173
rect -158 16931 -100 16943
rect -158 15955 -146 16931
rect -112 15955 -100 16931
rect -158 15943 -100 15955
rect 100 16931 158 16943
rect 100 15955 112 16931
rect 146 15955 158 16931
rect 100 15943 158 15955
rect -158 15713 -100 15725
rect -158 14737 -146 15713
rect -112 14737 -100 15713
rect -158 14725 -100 14737
rect 100 15713 158 15725
rect 100 14737 112 15713
rect 146 14737 158 15713
rect 100 14725 158 14737
rect -158 14495 -100 14507
rect -158 13519 -146 14495
rect -112 13519 -100 14495
rect -158 13507 -100 13519
rect 100 14495 158 14507
rect 100 13519 112 14495
rect 146 13519 158 14495
rect 100 13507 158 13519
rect -158 13277 -100 13289
rect -158 12301 -146 13277
rect -112 12301 -100 13277
rect -158 12289 -100 12301
rect 100 13277 158 13289
rect 100 12301 112 13277
rect 146 12301 158 13277
rect 100 12289 158 12301
rect -158 12059 -100 12071
rect -158 11083 -146 12059
rect -112 11083 -100 12059
rect -158 11071 -100 11083
rect 100 12059 158 12071
rect 100 11083 112 12059
rect 146 11083 158 12059
rect 100 11071 158 11083
rect -158 10841 -100 10853
rect -158 9865 -146 10841
rect -112 9865 -100 10841
rect -158 9853 -100 9865
rect 100 10841 158 10853
rect 100 9865 112 10841
rect 146 9865 158 10841
rect 100 9853 158 9865
rect -158 9623 -100 9635
rect -158 8647 -146 9623
rect -112 8647 -100 9623
rect -158 8635 -100 8647
rect 100 9623 158 9635
rect 100 8647 112 9623
rect 146 8647 158 9623
rect 100 8635 158 8647
rect -158 8405 -100 8417
rect -158 7429 -146 8405
rect -112 7429 -100 8405
rect -158 7417 -100 7429
rect 100 8405 158 8417
rect 100 7429 112 8405
rect 146 7429 158 8405
rect 100 7417 158 7429
rect -158 7187 -100 7199
rect -158 6211 -146 7187
rect -112 6211 -100 7187
rect -158 6199 -100 6211
rect 100 7187 158 7199
rect 100 6211 112 7187
rect 146 6211 158 7187
rect 100 6199 158 6211
rect -158 5969 -100 5981
rect -158 4993 -146 5969
rect -112 4993 -100 5969
rect -158 4981 -100 4993
rect 100 5969 158 5981
rect 100 4993 112 5969
rect 146 4993 158 5969
rect 100 4981 158 4993
rect -158 4751 -100 4763
rect -158 3775 -146 4751
rect -112 3775 -100 4751
rect -158 3763 -100 3775
rect 100 4751 158 4763
rect 100 3775 112 4751
rect 146 3775 158 4751
rect 100 3763 158 3775
rect -158 3533 -100 3545
rect -158 2557 -146 3533
rect -112 2557 -100 3533
rect -158 2545 -100 2557
rect 100 3533 158 3545
rect 100 2557 112 3533
rect 146 2557 158 3533
rect 100 2545 158 2557
rect -158 2315 -100 2327
rect -158 1339 -146 2315
rect -112 1339 -100 2315
rect -158 1327 -100 1339
rect 100 2315 158 2327
rect 100 1339 112 2315
rect 146 1339 158 2315
rect 100 1327 158 1339
rect -158 1097 -100 1109
rect -158 121 -146 1097
rect -112 121 -100 1097
rect -158 109 -100 121
rect 100 1097 158 1109
rect 100 121 112 1097
rect 146 121 158 1097
rect 100 109 158 121
rect -158 -121 -100 -109
rect -158 -1097 -146 -121
rect -112 -1097 -100 -121
rect -158 -1109 -100 -1097
rect 100 -121 158 -109
rect 100 -1097 112 -121
rect 146 -1097 158 -121
rect 100 -1109 158 -1097
rect -158 -1339 -100 -1327
rect -158 -2315 -146 -1339
rect -112 -2315 -100 -1339
rect -158 -2327 -100 -2315
rect 100 -1339 158 -1327
rect 100 -2315 112 -1339
rect 146 -2315 158 -1339
rect 100 -2327 158 -2315
rect -158 -2557 -100 -2545
rect -158 -3533 -146 -2557
rect -112 -3533 -100 -2557
rect -158 -3545 -100 -3533
rect 100 -2557 158 -2545
rect 100 -3533 112 -2557
rect 146 -3533 158 -2557
rect 100 -3545 158 -3533
rect -158 -3775 -100 -3763
rect -158 -4751 -146 -3775
rect -112 -4751 -100 -3775
rect -158 -4763 -100 -4751
rect 100 -3775 158 -3763
rect 100 -4751 112 -3775
rect 146 -4751 158 -3775
rect 100 -4763 158 -4751
rect -158 -4993 -100 -4981
rect -158 -5969 -146 -4993
rect -112 -5969 -100 -4993
rect -158 -5981 -100 -5969
rect 100 -4993 158 -4981
rect 100 -5969 112 -4993
rect 146 -5969 158 -4993
rect 100 -5981 158 -5969
rect -158 -6211 -100 -6199
rect -158 -7187 -146 -6211
rect -112 -7187 -100 -6211
rect -158 -7199 -100 -7187
rect 100 -6211 158 -6199
rect 100 -7187 112 -6211
rect 146 -7187 158 -6211
rect 100 -7199 158 -7187
rect -158 -7429 -100 -7417
rect -158 -8405 -146 -7429
rect -112 -8405 -100 -7429
rect -158 -8417 -100 -8405
rect 100 -7429 158 -7417
rect 100 -8405 112 -7429
rect 146 -8405 158 -7429
rect 100 -8417 158 -8405
rect -158 -8647 -100 -8635
rect -158 -9623 -146 -8647
rect -112 -9623 -100 -8647
rect -158 -9635 -100 -9623
rect 100 -8647 158 -8635
rect 100 -9623 112 -8647
rect 146 -9623 158 -8647
rect 100 -9635 158 -9623
rect -158 -9865 -100 -9853
rect -158 -10841 -146 -9865
rect -112 -10841 -100 -9865
rect -158 -10853 -100 -10841
rect 100 -9865 158 -9853
rect 100 -10841 112 -9865
rect 146 -10841 158 -9865
rect 100 -10853 158 -10841
rect -158 -11083 -100 -11071
rect -158 -12059 -146 -11083
rect -112 -12059 -100 -11083
rect -158 -12071 -100 -12059
rect 100 -11083 158 -11071
rect 100 -12059 112 -11083
rect 146 -12059 158 -11083
rect 100 -12071 158 -12059
rect -158 -12301 -100 -12289
rect -158 -13277 -146 -12301
rect -112 -13277 -100 -12301
rect -158 -13289 -100 -13277
rect 100 -12301 158 -12289
rect 100 -13277 112 -12301
rect 146 -13277 158 -12301
rect 100 -13289 158 -13277
rect -158 -13519 -100 -13507
rect -158 -14495 -146 -13519
rect -112 -14495 -100 -13519
rect -158 -14507 -100 -14495
rect 100 -13519 158 -13507
rect 100 -14495 112 -13519
rect 146 -14495 158 -13519
rect 100 -14507 158 -14495
rect -158 -14737 -100 -14725
rect -158 -15713 -146 -14737
rect -112 -15713 -100 -14737
rect -158 -15725 -100 -15713
rect 100 -14737 158 -14725
rect 100 -15713 112 -14737
rect 146 -15713 158 -14737
rect 100 -15725 158 -15713
rect -158 -15955 -100 -15943
rect -158 -16931 -146 -15955
rect -112 -16931 -100 -15955
rect -158 -16943 -100 -16931
rect 100 -15955 158 -15943
rect 100 -16931 112 -15955
rect 146 -16931 158 -15955
rect 100 -16943 158 -16931
rect -158 -17173 -100 -17161
rect -158 -18149 -146 -17173
rect -112 -18149 -100 -17173
rect -158 -18161 -100 -18149
rect 100 -17173 158 -17161
rect 100 -18149 112 -17173
rect 146 -18149 158 -17173
rect 100 -18161 158 -18149
rect -158 -18391 -100 -18379
rect -158 -19367 -146 -18391
rect -112 -19367 -100 -18391
rect -158 -19379 -100 -19367
rect 100 -18391 158 -18379
rect 100 -19367 112 -18391
rect 146 -19367 158 -18391
rect 100 -19379 158 -19367
rect -158 -19609 -100 -19597
rect -158 -20585 -146 -19609
rect -112 -20585 -100 -19609
rect -158 -20597 -100 -20585
rect 100 -19609 158 -19597
rect 100 -20585 112 -19609
rect 146 -20585 158 -19609
rect 100 -20597 158 -20585
rect -158 -20827 -100 -20815
rect -158 -21803 -146 -20827
rect -112 -21803 -100 -20827
rect -158 -21815 -100 -21803
rect 100 -20827 158 -20815
rect 100 -21803 112 -20827
rect 146 -21803 158 -20827
rect 100 -21815 158 -21803
rect -158 -22045 -100 -22033
rect -158 -23021 -146 -22045
rect -112 -23021 -100 -22045
rect -158 -23033 -100 -23021
rect 100 -22045 158 -22033
rect 100 -23021 112 -22045
rect 146 -23021 158 -22045
rect 100 -23033 158 -23021
rect -158 -23263 -100 -23251
rect -158 -24239 -146 -23263
rect -112 -24239 -100 -23263
rect -158 -24251 -100 -24239
rect 100 -23263 158 -23251
rect 100 -24239 112 -23263
rect 146 -24239 158 -23263
rect 100 -24251 158 -24239
rect -158 -24481 -100 -24469
rect -158 -25457 -146 -24481
rect -112 -25457 -100 -24481
rect -158 -25469 -100 -25457
rect 100 -24481 158 -24469
rect 100 -25457 112 -24481
rect 146 -25457 158 -24481
rect 100 -25469 158 -25457
rect -158 -25699 -100 -25687
rect -158 -26675 -146 -25699
rect -112 -26675 -100 -25699
rect -158 -26687 -100 -26675
rect 100 -25699 158 -25687
rect 100 -26675 112 -25699
rect 146 -26675 158 -25699
rect 100 -26687 158 -26675
rect -158 -26917 -100 -26905
rect -158 -27893 -146 -26917
rect -112 -27893 -100 -26917
rect -158 -27905 -100 -27893
rect 100 -26917 158 -26905
rect 100 -27893 112 -26917
rect 146 -27893 158 -26917
rect 100 -27905 158 -27893
rect -158 -28135 -100 -28123
rect -158 -29111 -146 -28135
rect -112 -29111 -100 -28135
rect -158 -29123 -100 -29111
rect 100 -28135 158 -28123
rect 100 -29111 112 -28135
rect 146 -29111 158 -28135
rect 100 -29123 158 -29111
rect -158 -29353 -100 -29341
rect -158 -30329 -146 -29353
rect -112 -30329 -100 -29353
rect -158 -30341 -100 -30329
rect 100 -29353 158 -29341
rect 100 -30329 112 -29353
rect 146 -30329 158 -29353
rect 100 -30341 158 -30329
rect -158 -30571 -100 -30559
rect -158 -31547 -146 -30571
rect -112 -31547 -100 -30571
rect -158 -31559 -100 -31547
rect 100 -30571 158 -30559
rect 100 -31547 112 -30571
rect 146 -31547 158 -30571
rect 100 -31559 158 -31547
rect -158 -31789 -100 -31777
rect -158 -32765 -146 -31789
rect -112 -32765 -100 -31789
rect -158 -32777 -100 -32765
rect 100 -31789 158 -31777
rect 100 -32765 112 -31789
rect 146 -32765 158 -31789
rect 100 -32777 158 -32765
rect -158 -33007 -100 -32995
rect -158 -33983 -146 -33007
rect -112 -33983 -100 -33007
rect -158 -33995 -100 -33983
rect 100 -33007 158 -32995
rect 100 -33983 112 -33007
rect 146 -33983 158 -33007
rect 100 -33995 158 -33983
rect -158 -34225 -100 -34213
rect -158 -35201 -146 -34225
rect -112 -35201 -100 -34225
rect -158 -35213 -100 -35201
rect 100 -34225 158 -34213
rect 100 -35201 112 -34225
rect 146 -35201 158 -34225
rect 100 -35213 158 -35201
rect -158 -35443 -100 -35431
rect -158 -36419 -146 -35443
rect -112 -36419 -100 -35443
rect -158 -36431 -100 -36419
rect 100 -35443 158 -35431
rect 100 -36419 112 -35443
rect 146 -36419 158 -35443
rect 100 -36431 158 -36419
rect -158 -36661 -100 -36649
rect -158 -37637 -146 -36661
rect -112 -37637 -100 -36661
rect -158 -37649 -100 -37637
rect 100 -36661 158 -36649
rect 100 -37637 112 -36661
rect 146 -37637 158 -36661
rect 100 -37649 158 -37637
rect -158 -37879 -100 -37867
rect -158 -38855 -146 -37879
rect -112 -38855 -100 -37879
rect -158 -38867 -100 -38855
rect 100 -37879 158 -37867
rect 100 -38855 112 -37879
rect 146 -38855 158 -37879
rect 100 -38867 158 -38855
rect -158 -39097 -100 -39085
rect -158 -40073 -146 -39097
rect -112 -40073 -100 -39097
rect -158 -40085 -100 -40073
rect 100 -39097 158 -39085
rect 100 -40073 112 -39097
rect 146 -40073 158 -39097
rect 100 -40085 158 -40073
rect -158 -40315 -100 -40303
rect -158 -41291 -146 -40315
rect -112 -41291 -100 -40315
rect -158 -41303 -100 -41291
rect 100 -40315 158 -40303
rect 100 -41291 112 -40315
rect 146 -41291 158 -40315
rect 100 -41303 158 -41291
rect -158 -41533 -100 -41521
rect -158 -42509 -146 -41533
rect -112 -42509 -100 -41533
rect -158 -42521 -100 -42509
rect 100 -41533 158 -41521
rect 100 -42509 112 -41533
rect 146 -42509 158 -41533
rect 100 -42521 158 -42509
rect -158 -42751 -100 -42739
rect -158 -43727 -146 -42751
rect -112 -43727 -100 -42751
rect -158 -43739 -100 -43727
rect 100 -42751 158 -42739
rect 100 -43727 112 -42751
rect 146 -43727 158 -42751
rect 100 -43739 158 -43727
rect -158 -43969 -100 -43957
rect -158 -44945 -146 -43969
rect -112 -44945 -100 -43969
rect -158 -44957 -100 -44945
rect 100 -43969 158 -43957
rect 100 -44945 112 -43969
rect 146 -44945 158 -43969
rect 100 -44957 158 -44945
rect -158 -45187 -100 -45175
rect -158 -46163 -146 -45187
rect -112 -46163 -100 -45187
rect -158 -46175 -100 -46163
rect 100 -45187 158 -45175
rect 100 -46163 112 -45187
rect 146 -46163 158 -45187
rect 100 -46175 158 -46163
rect -158 -46405 -100 -46393
rect -158 -47381 -146 -46405
rect -112 -47381 -100 -46405
rect -158 -47393 -100 -47381
rect 100 -46405 158 -46393
rect 100 -47381 112 -46405
rect 146 -47381 158 -46405
rect 100 -47393 158 -47381
rect -158 -47623 -100 -47611
rect -158 -48599 -146 -47623
rect -112 -48599 -100 -47623
rect -158 -48611 -100 -48599
rect 100 -47623 158 -47611
rect 100 -48599 112 -47623
rect 146 -48599 158 -47623
rect 100 -48611 158 -48599
rect -158 -48841 -100 -48829
rect -158 -49817 -146 -48841
rect -112 -49817 -100 -48841
rect -158 -49829 -100 -49817
rect 100 -48841 158 -48829
rect 100 -49817 112 -48841
rect 146 -49817 158 -48841
rect 100 -49829 158 -49817
rect -158 -50059 -100 -50047
rect -158 -51035 -146 -50059
rect -112 -51035 -100 -50059
rect -158 -51047 -100 -51035
rect 100 -50059 158 -50047
rect 100 -51035 112 -50059
rect 146 -51035 158 -50059
rect 100 -51047 158 -51035
rect -158 -51277 -100 -51265
rect -158 -52253 -146 -51277
rect -112 -52253 -100 -51277
rect -158 -52265 -100 -52253
rect 100 -51277 158 -51265
rect 100 -52253 112 -51277
rect 146 -52253 158 -51277
rect 100 -52265 158 -52253
rect -158 -52495 -100 -52483
rect -158 -53471 -146 -52495
rect -112 -53471 -100 -52495
rect -158 -53483 -100 -53471
rect 100 -52495 158 -52483
rect 100 -53471 112 -52495
rect 146 -53471 158 -52495
rect 100 -53483 158 -53471
rect -158 -53713 -100 -53701
rect -158 -54689 -146 -53713
rect -112 -54689 -100 -53713
rect -158 -54701 -100 -54689
rect 100 -53713 158 -53701
rect 100 -54689 112 -53713
rect 146 -54689 158 -53713
rect 100 -54701 158 -54689
rect -158 -54931 -100 -54919
rect -158 -55907 -146 -54931
rect -112 -55907 -100 -54931
rect -158 -55919 -100 -55907
rect 100 -54931 158 -54919
rect 100 -55907 112 -54931
rect 146 -55907 158 -54931
rect 100 -55919 158 -55907
rect -158 -56149 -100 -56137
rect -158 -57125 -146 -56149
rect -112 -57125 -100 -56149
rect -158 -57137 -100 -57125
rect 100 -56149 158 -56137
rect 100 -57125 112 -56149
rect 146 -57125 158 -56149
rect 100 -57137 158 -57125
rect -158 -57367 -100 -57355
rect -158 -58343 -146 -57367
rect -112 -58343 -100 -57367
rect -158 -58355 -100 -58343
rect 100 -57367 158 -57355
rect 100 -58343 112 -57367
rect 146 -58343 158 -57367
rect 100 -58355 158 -58343
rect -158 -58585 -100 -58573
rect -158 -59561 -146 -58585
rect -112 -59561 -100 -58585
rect -158 -59573 -100 -59561
rect 100 -58585 158 -58573
rect 100 -59561 112 -58585
rect 146 -59561 158 -58585
rect 100 -59573 158 -59561
rect -158 -59803 -100 -59791
rect -158 -60779 -146 -59803
rect -112 -60779 -100 -59803
rect -158 -60791 -100 -60779
rect 100 -59803 158 -59791
rect 100 -60779 112 -59803
rect 146 -60779 158 -59803
rect 100 -60791 158 -60779
rect -158 -61021 -100 -61009
rect -158 -61997 -146 -61021
rect -112 -61997 -100 -61021
rect -158 -62009 -100 -61997
rect 100 -61021 158 -61009
rect 100 -61997 112 -61021
rect 146 -61997 158 -61021
rect 100 -62009 158 -61997
rect -158 -62239 -100 -62227
rect -158 -63215 -146 -62239
rect -112 -63215 -100 -62239
rect -158 -63227 -100 -63215
rect 100 -62239 158 -62227
rect 100 -63215 112 -62239
rect 146 -63215 158 -62239
rect 100 -63227 158 -63215
rect -158 -63457 -100 -63445
rect -158 -64433 -146 -63457
rect -112 -64433 -100 -63457
rect -158 -64445 -100 -64433
rect 100 -63457 158 -63445
rect 100 -64433 112 -63457
rect 146 -64433 158 -63457
rect 100 -64445 158 -64433
rect -158 -64675 -100 -64663
rect -158 -65651 -146 -64675
rect -112 -65651 -100 -64675
rect -158 -65663 -100 -65651
rect 100 -64675 158 -64663
rect 100 -65651 112 -64675
rect 146 -65651 158 -64675
rect 100 -65663 158 -65651
rect -158 -65893 -100 -65881
rect -158 -66869 -146 -65893
rect -112 -66869 -100 -65893
rect -158 -66881 -100 -66869
rect 100 -65893 158 -65881
rect 100 -66869 112 -65893
rect 146 -66869 158 -65893
rect 100 -66881 158 -66869
rect -158 -67111 -100 -67099
rect -158 -68087 -146 -67111
rect -112 -68087 -100 -67111
rect -158 -68099 -100 -68087
rect 100 -67111 158 -67099
rect 100 -68087 112 -67111
rect 146 -68087 158 -67111
rect 100 -68099 158 -68087
rect -158 -68329 -100 -68317
rect -158 -69305 -146 -68329
rect -112 -69305 -100 -68329
rect -158 -69317 -100 -69305
rect 100 -68329 158 -68317
rect 100 -69305 112 -68329
rect 146 -69305 158 -68329
rect 100 -69317 158 -69305
rect -158 -69547 -100 -69535
rect -158 -70523 -146 -69547
rect -112 -70523 -100 -69547
rect -158 -70535 -100 -70523
rect 100 -69547 158 -69535
rect 100 -70523 112 -69547
rect 146 -70523 158 -69547
rect 100 -70535 158 -70523
rect -158 -70765 -100 -70753
rect -158 -71741 -146 -70765
rect -112 -71741 -100 -70765
rect -158 -71753 -100 -71741
rect 100 -70765 158 -70753
rect 100 -71741 112 -70765
rect 146 -71741 158 -70765
rect 100 -71753 158 -71741
rect -158 -71983 -100 -71971
rect -158 -72959 -146 -71983
rect -112 -72959 -100 -71983
rect -158 -72971 -100 -72959
rect 100 -71983 158 -71971
rect 100 -72959 112 -71983
rect 146 -72959 158 -71983
rect 100 -72971 158 -72959
rect -158 -73201 -100 -73189
rect -158 -74177 -146 -73201
rect -112 -74177 -100 -73201
rect -158 -74189 -100 -74177
rect 100 -73201 158 -73189
rect 100 -74177 112 -73201
rect 146 -74177 158 -73201
rect 100 -74189 158 -74177
rect -158 -74419 -100 -74407
rect -158 -75395 -146 -74419
rect -112 -75395 -100 -74419
rect -158 -75407 -100 -75395
rect 100 -74419 158 -74407
rect 100 -75395 112 -74419
rect 146 -75395 158 -74419
rect 100 -75407 158 -75395
rect -158 -75637 -100 -75625
rect -158 -76613 -146 -75637
rect -112 -76613 -100 -75637
rect -158 -76625 -100 -76613
rect 100 -75637 158 -75625
rect 100 -76613 112 -75637
rect 146 -76613 158 -75637
rect 100 -76625 158 -76613
rect -158 -76855 -100 -76843
rect -158 -77831 -146 -76855
rect -112 -77831 -100 -76855
rect -158 -77843 -100 -77831
rect 100 -76855 158 -76843
rect 100 -77831 112 -76855
rect 146 -77831 158 -76855
rect 100 -77843 158 -77831
rect -158 -78073 -100 -78061
rect -158 -79049 -146 -78073
rect -112 -79049 -100 -78073
rect -158 -79061 -100 -79049
rect 100 -78073 158 -78061
rect 100 -79049 112 -78073
rect 146 -79049 158 -78073
rect 100 -79061 158 -79049
rect -158 -79291 -100 -79279
rect -158 -80267 -146 -79291
rect -112 -80267 -100 -79291
rect -158 -80279 -100 -80267
rect 100 -79291 158 -79279
rect 100 -80267 112 -79291
rect 146 -80267 158 -79291
rect 100 -80279 158 -80267
rect -158 -80509 -100 -80497
rect -158 -81485 -146 -80509
rect -112 -81485 -100 -80509
rect -158 -81497 -100 -81485
rect 100 -80509 158 -80497
rect 100 -81485 112 -80509
rect 146 -81485 158 -80509
rect 100 -81497 158 -81485
rect -158 -81727 -100 -81715
rect -158 -82703 -146 -81727
rect -112 -82703 -100 -81727
rect -158 -82715 -100 -82703
rect 100 -81727 158 -81715
rect 100 -82703 112 -81727
rect 146 -82703 158 -81727
rect 100 -82715 158 -82703
rect -158 -82945 -100 -82933
rect -158 -83921 -146 -82945
rect -112 -83921 -100 -82945
rect -158 -83933 -100 -83921
rect 100 -82945 158 -82933
rect 100 -83921 112 -82945
rect 146 -83921 158 -82945
rect 100 -83933 158 -83921
rect -158 -84163 -100 -84151
rect -158 -85139 -146 -84163
rect -112 -85139 -100 -84163
rect -158 -85151 -100 -85139
rect 100 -84163 158 -84151
rect 100 -85139 112 -84163
rect 146 -85139 158 -84163
rect 100 -85151 158 -85139
rect -158 -85381 -100 -85369
rect -158 -86357 -146 -85381
rect -112 -86357 -100 -85381
rect -158 -86369 -100 -86357
rect 100 -85381 158 -85369
rect 100 -86357 112 -85381
rect 146 -86357 158 -85381
rect 100 -86369 158 -86357
rect -158 -86599 -100 -86587
rect -158 -87575 -146 -86599
rect -112 -87575 -100 -86599
rect -158 -87587 -100 -87575
rect 100 -86599 158 -86587
rect 100 -87575 112 -86599
rect 146 -87575 158 -86599
rect 100 -87587 158 -87575
rect -158 -87817 -100 -87805
rect -158 -88793 -146 -87817
rect -112 -88793 -100 -87817
rect -158 -88805 -100 -88793
rect 100 -87817 158 -87805
rect 100 -88793 112 -87817
rect 146 -88793 158 -87817
rect 100 -88805 158 -88793
rect -158 -89035 -100 -89023
rect -158 -90011 -146 -89035
rect -112 -90011 -100 -89035
rect -158 -90023 -100 -90011
rect 100 -89035 158 -89023
rect 100 -90011 112 -89035
rect 146 -90011 158 -89035
rect 100 -90023 158 -90011
rect -158 -90253 -100 -90241
rect -158 -91229 -146 -90253
rect -112 -91229 -100 -90253
rect -158 -91241 -100 -91229
rect 100 -90253 158 -90241
rect 100 -91229 112 -90253
rect 146 -91229 158 -90253
rect 100 -91241 158 -91229
rect -158 -91471 -100 -91459
rect -158 -92447 -146 -91471
rect -112 -92447 -100 -91471
rect -158 -92459 -100 -92447
rect 100 -91471 158 -91459
rect 100 -92447 112 -91471
rect 146 -92447 158 -91471
rect 100 -92459 158 -92447
rect -158 -92689 -100 -92677
rect -158 -93665 -146 -92689
rect -112 -93665 -100 -92689
rect -158 -93677 -100 -93665
rect 100 -92689 158 -92677
rect 100 -93665 112 -92689
rect 146 -93665 158 -92689
rect 100 -93677 158 -93665
rect -158 -93907 -100 -93895
rect -158 -94883 -146 -93907
rect -112 -94883 -100 -93907
rect -158 -94895 -100 -94883
rect 100 -93907 158 -93895
rect 100 -94883 112 -93907
rect 146 -94883 158 -93907
rect 100 -94895 158 -94883
rect -158 -95125 -100 -95113
rect -158 -96101 -146 -95125
rect -112 -96101 -100 -95125
rect -158 -96113 -100 -96101
rect 100 -95125 158 -95113
rect 100 -96101 112 -95125
rect 146 -96101 158 -95125
rect 100 -96113 158 -96101
rect -158 -96343 -100 -96331
rect -158 -97319 -146 -96343
rect -112 -97319 -100 -96343
rect -158 -97331 -100 -97319
rect 100 -96343 158 -96331
rect 100 -97319 112 -96343
rect 146 -97319 158 -96343
rect 100 -97331 158 -97319
rect -158 -97561 -100 -97549
rect -158 -98537 -146 -97561
rect -112 -98537 -100 -97561
rect -158 -98549 -100 -98537
rect 100 -97561 158 -97549
rect 100 -98537 112 -97561
rect 146 -98537 158 -97561
rect 100 -98549 158 -98537
rect -158 -98779 -100 -98767
rect -158 -99755 -146 -98779
rect -112 -99755 -100 -98779
rect -158 -99767 -100 -99755
rect 100 -98779 158 -98767
rect 100 -99755 112 -98779
rect 146 -99755 158 -98779
rect 100 -99767 158 -99755
rect -158 -99997 -100 -99985
rect -158 -100973 -146 -99997
rect -112 -100973 -100 -99997
rect -158 -100985 -100 -100973
rect 100 -99997 158 -99985
rect 100 -100973 112 -99997
rect 146 -100973 158 -99997
rect 100 -100985 158 -100973
rect -158 -101215 -100 -101203
rect -158 -102191 -146 -101215
rect -112 -102191 -100 -101215
rect -158 -102203 -100 -102191
rect 100 -101215 158 -101203
rect 100 -102191 112 -101215
rect 146 -102191 158 -101215
rect 100 -102203 158 -102191
rect -158 -102433 -100 -102421
rect -158 -103409 -146 -102433
rect -112 -103409 -100 -102433
rect -158 -103421 -100 -103409
rect 100 -102433 158 -102421
rect 100 -103409 112 -102433
rect 146 -103409 158 -102433
rect 100 -103421 158 -103409
rect -158 -103651 -100 -103639
rect -158 -104627 -146 -103651
rect -112 -104627 -100 -103651
rect -158 -104639 -100 -104627
rect 100 -103651 158 -103639
rect 100 -104627 112 -103651
rect 146 -104627 158 -103651
rect 100 -104639 158 -104627
rect -158 -104869 -100 -104857
rect -158 -105845 -146 -104869
rect -112 -105845 -100 -104869
rect -158 -105857 -100 -105845
rect 100 -104869 158 -104857
rect 100 -105845 112 -104869
rect 146 -105845 158 -104869
rect 100 -105857 158 -105845
rect -158 -106087 -100 -106075
rect -158 -107063 -146 -106087
rect -112 -107063 -100 -106087
rect -158 -107075 -100 -107063
rect 100 -106087 158 -106075
rect 100 -107063 112 -106087
rect 146 -107063 158 -106087
rect 100 -107075 158 -107063
rect -158 -107305 -100 -107293
rect -158 -108281 -146 -107305
rect -112 -108281 -100 -107305
rect -158 -108293 -100 -108281
rect 100 -107305 158 -107293
rect 100 -108281 112 -107305
rect 146 -108281 158 -107305
rect 100 -108293 158 -108281
rect -158 -108523 -100 -108511
rect -158 -109499 -146 -108523
rect -112 -109499 -100 -108523
rect -158 -109511 -100 -109499
rect 100 -108523 158 -108511
rect 100 -109499 112 -108523
rect 146 -109499 158 -108523
rect 100 -109511 158 -109499
rect -158 -109741 -100 -109729
rect -158 -110717 -146 -109741
rect -112 -110717 -100 -109741
rect -158 -110729 -100 -110717
rect 100 -109741 158 -109729
rect 100 -110717 112 -109741
rect 146 -110717 158 -109741
rect 100 -110729 158 -110717
rect -158 -110959 -100 -110947
rect -158 -111935 -146 -110959
rect -112 -111935 -100 -110959
rect -158 -111947 -100 -111935
rect 100 -110959 158 -110947
rect 100 -111935 112 -110959
rect 146 -111935 158 -110959
rect 100 -111947 158 -111935
rect -158 -112177 -100 -112165
rect -158 -113153 -146 -112177
rect -112 -113153 -100 -112177
rect -158 -113165 -100 -113153
rect 100 -112177 158 -112165
rect 100 -113153 112 -112177
rect 146 -113153 158 -112177
rect 100 -113165 158 -113153
rect -158 -113395 -100 -113383
rect -158 -114371 -146 -113395
rect -112 -114371 -100 -113395
rect -158 -114383 -100 -114371
rect 100 -113395 158 -113383
rect 100 -114371 112 -113395
rect 146 -114371 158 -113395
rect 100 -114383 158 -114371
rect -158 -114613 -100 -114601
rect -158 -115589 -146 -114613
rect -112 -115589 -100 -114613
rect -158 -115601 -100 -115589
rect 100 -114613 158 -114601
rect 100 -115589 112 -114613
rect 146 -115589 158 -114613
rect 100 -115601 158 -115589
rect -158 -115831 -100 -115819
rect -158 -116807 -146 -115831
rect -112 -116807 -100 -115831
rect -158 -116819 -100 -116807
rect 100 -115831 158 -115819
rect 100 -116807 112 -115831
rect 146 -116807 158 -115831
rect 100 -116819 158 -116807
rect -158 -117049 -100 -117037
rect -158 -118025 -146 -117049
rect -112 -118025 -100 -117049
rect -158 -118037 -100 -118025
rect 100 -117049 158 -117037
rect 100 -118025 112 -117049
rect 146 -118025 158 -117049
rect 100 -118037 158 -118025
rect -158 -118267 -100 -118255
rect -158 -119243 -146 -118267
rect -112 -119243 -100 -118267
rect -158 -119255 -100 -119243
rect 100 -118267 158 -118255
rect 100 -119243 112 -118267
rect 146 -119243 158 -118267
rect 100 -119255 158 -119243
rect -158 -119485 -100 -119473
rect -158 -120461 -146 -119485
rect -112 -120461 -100 -119485
rect -158 -120473 -100 -120461
rect 100 -119485 158 -119473
rect 100 -120461 112 -119485
rect 146 -120461 158 -119485
rect 100 -120473 158 -120461
rect -158 -120703 -100 -120691
rect -158 -121679 -146 -120703
rect -112 -121679 -100 -120703
rect -158 -121691 -100 -121679
rect 100 -120703 158 -120691
rect 100 -121679 112 -120703
rect 146 -121679 158 -120703
rect 100 -121691 158 -121679
<< mvndiffc >>
rect -146 120703 -112 121679
rect 112 120703 146 121679
rect -146 119485 -112 120461
rect 112 119485 146 120461
rect -146 118267 -112 119243
rect 112 118267 146 119243
rect -146 117049 -112 118025
rect 112 117049 146 118025
rect -146 115831 -112 116807
rect 112 115831 146 116807
rect -146 114613 -112 115589
rect 112 114613 146 115589
rect -146 113395 -112 114371
rect 112 113395 146 114371
rect -146 112177 -112 113153
rect 112 112177 146 113153
rect -146 110959 -112 111935
rect 112 110959 146 111935
rect -146 109741 -112 110717
rect 112 109741 146 110717
rect -146 108523 -112 109499
rect 112 108523 146 109499
rect -146 107305 -112 108281
rect 112 107305 146 108281
rect -146 106087 -112 107063
rect 112 106087 146 107063
rect -146 104869 -112 105845
rect 112 104869 146 105845
rect -146 103651 -112 104627
rect 112 103651 146 104627
rect -146 102433 -112 103409
rect 112 102433 146 103409
rect -146 101215 -112 102191
rect 112 101215 146 102191
rect -146 99997 -112 100973
rect 112 99997 146 100973
rect -146 98779 -112 99755
rect 112 98779 146 99755
rect -146 97561 -112 98537
rect 112 97561 146 98537
rect -146 96343 -112 97319
rect 112 96343 146 97319
rect -146 95125 -112 96101
rect 112 95125 146 96101
rect -146 93907 -112 94883
rect 112 93907 146 94883
rect -146 92689 -112 93665
rect 112 92689 146 93665
rect -146 91471 -112 92447
rect 112 91471 146 92447
rect -146 90253 -112 91229
rect 112 90253 146 91229
rect -146 89035 -112 90011
rect 112 89035 146 90011
rect -146 87817 -112 88793
rect 112 87817 146 88793
rect -146 86599 -112 87575
rect 112 86599 146 87575
rect -146 85381 -112 86357
rect 112 85381 146 86357
rect -146 84163 -112 85139
rect 112 84163 146 85139
rect -146 82945 -112 83921
rect 112 82945 146 83921
rect -146 81727 -112 82703
rect 112 81727 146 82703
rect -146 80509 -112 81485
rect 112 80509 146 81485
rect -146 79291 -112 80267
rect 112 79291 146 80267
rect -146 78073 -112 79049
rect 112 78073 146 79049
rect -146 76855 -112 77831
rect 112 76855 146 77831
rect -146 75637 -112 76613
rect 112 75637 146 76613
rect -146 74419 -112 75395
rect 112 74419 146 75395
rect -146 73201 -112 74177
rect 112 73201 146 74177
rect -146 71983 -112 72959
rect 112 71983 146 72959
rect -146 70765 -112 71741
rect 112 70765 146 71741
rect -146 69547 -112 70523
rect 112 69547 146 70523
rect -146 68329 -112 69305
rect 112 68329 146 69305
rect -146 67111 -112 68087
rect 112 67111 146 68087
rect -146 65893 -112 66869
rect 112 65893 146 66869
rect -146 64675 -112 65651
rect 112 64675 146 65651
rect -146 63457 -112 64433
rect 112 63457 146 64433
rect -146 62239 -112 63215
rect 112 62239 146 63215
rect -146 61021 -112 61997
rect 112 61021 146 61997
rect -146 59803 -112 60779
rect 112 59803 146 60779
rect -146 58585 -112 59561
rect 112 58585 146 59561
rect -146 57367 -112 58343
rect 112 57367 146 58343
rect -146 56149 -112 57125
rect 112 56149 146 57125
rect -146 54931 -112 55907
rect 112 54931 146 55907
rect -146 53713 -112 54689
rect 112 53713 146 54689
rect -146 52495 -112 53471
rect 112 52495 146 53471
rect -146 51277 -112 52253
rect 112 51277 146 52253
rect -146 50059 -112 51035
rect 112 50059 146 51035
rect -146 48841 -112 49817
rect 112 48841 146 49817
rect -146 47623 -112 48599
rect 112 47623 146 48599
rect -146 46405 -112 47381
rect 112 46405 146 47381
rect -146 45187 -112 46163
rect 112 45187 146 46163
rect -146 43969 -112 44945
rect 112 43969 146 44945
rect -146 42751 -112 43727
rect 112 42751 146 43727
rect -146 41533 -112 42509
rect 112 41533 146 42509
rect -146 40315 -112 41291
rect 112 40315 146 41291
rect -146 39097 -112 40073
rect 112 39097 146 40073
rect -146 37879 -112 38855
rect 112 37879 146 38855
rect -146 36661 -112 37637
rect 112 36661 146 37637
rect -146 35443 -112 36419
rect 112 35443 146 36419
rect -146 34225 -112 35201
rect 112 34225 146 35201
rect -146 33007 -112 33983
rect 112 33007 146 33983
rect -146 31789 -112 32765
rect 112 31789 146 32765
rect -146 30571 -112 31547
rect 112 30571 146 31547
rect -146 29353 -112 30329
rect 112 29353 146 30329
rect -146 28135 -112 29111
rect 112 28135 146 29111
rect -146 26917 -112 27893
rect 112 26917 146 27893
rect -146 25699 -112 26675
rect 112 25699 146 26675
rect -146 24481 -112 25457
rect 112 24481 146 25457
rect -146 23263 -112 24239
rect 112 23263 146 24239
rect -146 22045 -112 23021
rect 112 22045 146 23021
rect -146 20827 -112 21803
rect 112 20827 146 21803
rect -146 19609 -112 20585
rect 112 19609 146 20585
rect -146 18391 -112 19367
rect 112 18391 146 19367
rect -146 17173 -112 18149
rect 112 17173 146 18149
rect -146 15955 -112 16931
rect 112 15955 146 16931
rect -146 14737 -112 15713
rect 112 14737 146 15713
rect -146 13519 -112 14495
rect 112 13519 146 14495
rect -146 12301 -112 13277
rect 112 12301 146 13277
rect -146 11083 -112 12059
rect 112 11083 146 12059
rect -146 9865 -112 10841
rect 112 9865 146 10841
rect -146 8647 -112 9623
rect 112 8647 146 9623
rect -146 7429 -112 8405
rect 112 7429 146 8405
rect -146 6211 -112 7187
rect 112 6211 146 7187
rect -146 4993 -112 5969
rect 112 4993 146 5969
rect -146 3775 -112 4751
rect 112 3775 146 4751
rect -146 2557 -112 3533
rect 112 2557 146 3533
rect -146 1339 -112 2315
rect 112 1339 146 2315
rect -146 121 -112 1097
rect 112 121 146 1097
rect -146 -1097 -112 -121
rect 112 -1097 146 -121
rect -146 -2315 -112 -1339
rect 112 -2315 146 -1339
rect -146 -3533 -112 -2557
rect 112 -3533 146 -2557
rect -146 -4751 -112 -3775
rect 112 -4751 146 -3775
rect -146 -5969 -112 -4993
rect 112 -5969 146 -4993
rect -146 -7187 -112 -6211
rect 112 -7187 146 -6211
rect -146 -8405 -112 -7429
rect 112 -8405 146 -7429
rect -146 -9623 -112 -8647
rect 112 -9623 146 -8647
rect -146 -10841 -112 -9865
rect 112 -10841 146 -9865
rect -146 -12059 -112 -11083
rect 112 -12059 146 -11083
rect -146 -13277 -112 -12301
rect 112 -13277 146 -12301
rect -146 -14495 -112 -13519
rect 112 -14495 146 -13519
rect -146 -15713 -112 -14737
rect 112 -15713 146 -14737
rect -146 -16931 -112 -15955
rect 112 -16931 146 -15955
rect -146 -18149 -112 -17173
rect 112 -18149 146 -17173
rect -146 -19367 -112 -18391
rect 112 -19367 146 -18391
rect -146 -20585 -112 -19609
rect 112 -20585 146 -19609
rect -146 -21803 -112 -20827
rect 112 -21803 146 -20827
rect -146 -23021 -112 -22045
rect 112 -23021 146 -22045
rect -146 -24239 -112 -23263
rect 112 -24239 146 -23263
rect -146 -25457 -112 -24481
rect 112 -25457 146 -24481
rect -146 -26675 -112 -25699
rect 112 -26675 146 -25699
rect -146 -27893 -112 -26917
rect 112 -27893 146 -26917
rect -146 -29111 -112 -28135
rect 112 -29111 146 -28135
rect -146 -30329 -112 -29353
rect 112 -30329 146 -29353
rect -146 -31547 -112 -30571
rect 112 -31547 146 -30571
rect -146 -32765 -112 -31789
rect 112 -32765 146 -31789
rect -146 -33983 -112 -33007
rect 112 -33983 146 -33007
rect -146 -35201 -112 -34225
rect 112 -35201 146 -34225
rect -146 -36419 -112 -35443
rect 112 -36419 146 -35443
rect -146 -37637 -112 -36661
rect 112 -37637 146 -36661
rect -146 -38855 -112 -37879
rect 112 -38855 146 -37879
rect -146 -40073 -112 -39097
rect 112 -40073 146 -39097
rect -146 -41291 -112 -40315
rect 112 -41291 146 -40315
rect -146 -42509 -112 -41533
rect 112 -42509 146 -41533
rect -146 -43727 -112 -42751
rect 112 -43727 146 -42751
rect -146 -44945 -112 -43969
rect 112 -44945 146 -43969
rect -146 -46163 -112 -45187
rect 112 -46163 146 -45187
rect -146 -47381 -112 -46405
rect 112 -47381 146 -46405
rect -146 -48599 -112 -47623
rect 112 -48599 146 -47623
rect -146 -49817 -112 -48841
rect 112 -49817 146 -48841
rect -146 -51035 -112 -50059
rect 112 -51035 146 -50059
rect -146 -52253 -112 -51277
rect 112 -52253 146 -51277
rect -146 -53471 -112 -52495
rect 112 -53471 146 -52495
rect -146 -54689 -112 -53713
rect 112 -54689 146 -53713
rect -146 -55907 -112 -54931
rect 112 -55907 146 -54931
rect -146 -57125 -112 -56149
rect 112 -57125 146 -56149
rect -146 -58343 -112 -57367
rect 112 -58343 146 -57367
rect -146 -59561 -112 -58585
rect 112 -59561 146 -58585
rect -146 -60779 -112 -59803
rect 112 -60779 146 -59803
rect -146 -61997 -112 -61021
rect 112 -61997 146 -61021
rect -146 -63215 -112 -62239
rect 112 -63215 146 -62239
rect -146 -64433 -112 -63457
rect 112 -64433 146 -63457
rect -146 -65651 -112 -64675
rect 112 -65651 146 -64675
rect -146 -66869 -112 -65893
rect 112 -66869 146 -65893
rect -146 -68087 -112 -67111
rect 112 -68087 146 -67111
rect -146 -69305 -112 -68329
rect 112 -69305 146 -68329
rect -146 -70523 -112 -69547
rect 112 -70523 146 -69547
rect -146 -71741 -112 -70765
rect 112 -71741 146 -70765
rect -146 -72959 -112 -71983
rect 112 -72959 146 -71983
rect -146 -74177 -112 -73201
rect 112 -74177 146 -73201
rect -146 -75395 -112 -74419
rect 112 -75395 146 -74419
rect -146 -76613 -112 -75637
rect 112 -76613 146 -75637
rect -146 -77831 -112 -76855
rect 112 -77831 146 -76855
rect -146 -79049 -112 -78073
rect 112 -79049 146 -78073
rect -146 -80267 -112 -79291
rect 112 -80267 146 -79291
rect -146 -81485 -112 -80509
rect 112 -81485 146 -80509
rect -146 -82703 -112 -81727
rect 112 -82703 146 -81727
rect -146 -83921 -112 -82945
rect 112 -83921 146 -82945
rect -146 -85139 -112 -84163
rect 112 -85139 146 -84163
rect -146 -86357 -112 -85381
rect 112 -86357 146 -85381
rect -146 -87575 -112 -86599
rect 112 -87575 146 -86599
rect -146 -88793 -112 -87817
rect 112 -88793 146 -87817
rect -146 -90011 -112 -89035
rect 112 -90011 146 -89035
rect -146 -91229 -112 -90253
rect 112 -91229 146 -90253
rect -146 -92447 -112 -91471
rect 112 -92447 146 -91471
rect -146 -93665 -112 -92689
rect 112 -93665 146 -92689
rect -146 -94883 -112 -93907
rect 112 -94883 146 -93907
rect -146 -96101 -112 -95125
rect 112 -96101 146 -95125
rect -146 -97319 -112 -96343
rect 112 -97319 146 -96343
rect -146 -98537 -112 -97561
rect 112 -98537 146 -97561
rect -146 -99755 -112 -98779
rect 112 -99755 146 -98779
rect -146 -100973 -112 -99997
rect 112 -100973 146 -99997
rect -146 -102191 -112 -101215
rect 112 -102191 146 -101215
rect -146 -103409 -112 -102433
rect 112 -103409 146 -102433
rect -146 -104627 -112 -103651
rect 112 -104627 146 -103651
rect -146 -105845 -112 -104869
rect 112 -105845 146 -104869
rect -146 -107063 -112 -106087
rect 112 -107063 146 -106087
rect -146 -108281 -112 -107305
rect 112 -108281 146 -107305
rect -146 -109499 -112 -108523
rect 112 -109499 146 -108523
rect -146 -110717 -112 -109741
rect 112 -110717 146 -109741
rect -146 -111935 -112 -110959
rect 112 -111935 146 -110959
rect -146 -113153 -112 -112177
rect 112 -113153 146 -112177
rect -146 -114371 -112 -113395
rect 112 -114371 146 -113395
rect -146 -115589 -112 -114613
rect 112 -115589 146 -114613
rect -146 -116807 -112 -115831
rect 112 -116807 146 -115831
rect -146 -118025 -112 -117049
rect 112 -118025 146 -117049
rect -146 -119243 -112 -118267
rect 112 -119243 146 -118267
rect -146 -120461 -112 -119485
rect 112 -120461 146 -119485
rect -146 -121679 -112 -120703
rect 112 -121679 146 -120703
<< mvpsubdiff >>
rect -292 121901 292 121913
rect -292 121867 -184 121901
rect 184 121867 292 121901
rect -292 121855 292 121867
rect -292 121805 -234 121855
rect -292 -121805 -280 121805
rect -246 -121805 -234 121805
rect 234 121805 292 121855
rect -292 -121855 -234 -121805
rect 234 -121805 246 121805
rect 280 -121805 292 121805
rect 234 -121855 292 -121805
rect -292 -121867 292 -121855
rect -292 -121901 -184 -121867
rect 184 -121901 292 -121867
rect -292 -121913 292 -121901
<< mvpsubdiffcont >>
rect -184 121867 184 121901
rect -280 -121805 -246 121805
rect 246 -121805 280 121805
rect -184 -121901 184 -121867
<< poly >>
rect -100 121763 100 121779
rect -100 121729 -84 121763
rect 84 121729 100 121763
rect -100 121691 100 121729
rect -100 120653 100 120691
rect -100 120619 -84 120653
rect 84 120619 100 120653
rect -100 120603 100 120619
rect -100 120545 100 120561
rect -100 120511 -84 120545
rect 84 120511 100 120545
rect -100 120473 100 120511
rect -100 119435 100 119473
rect -100 119401 -84 119435
rect 84 119401 100 119435
rect -100 119385 100 119401
rect -100 119327 100 119343
rect -100 119293 -84 119327
rect 84 119293 100 119327
rect -100 119255 100 119293
rect -100 118217 100 118255
rect -100 118183 -84 118217
rect 84 118183 100 118217
rect -100 118167 100 118183
rect -100 118109 100 118125
rect -100 118075 -84 118109
rect 84 118075 100 118109
rect -100 118037 100 118075
rect -100 116999 100 117037
rect -100 116965 -84 116999
rect 84 116965 100 116999
rect -100 116949 100 116965
rect -100 116891 100 116907
rect -100 116857 -84 116891
rect 84 116857 100 116891
rect -100 116819 100 116857
rect -100 115781 100 115819
rect -100 115747 -84 115781
rect 84 115747 100 115781
rect -100 115731 100 115747
rect -100 115673 100 115689
rect -100 115639 -84 115673
rect 84 115639 100 115673
rect -100 115601 100 115639
rect -100 114563 100 114601
rect -100 114529 -84 114563
rect 84 114529 100 114563
rect -100 114513 100 114529
rect -100 114455 100 114471
rect -100 114421 -84 114455
rect 84 114421 100 114455
rect -100 114383 100 114421
rect -100 113345 100 113383
rect -100 113311 -84 113345
rect 84 113311 100 113345
rect -100 113295 100 113311
rect -100 113237 100 113253
rect -100 113203 -84 113237
rect 84 113203 100 113237
rect -100 113165 100 113203
rect -100 112127 100 112165
rect -100 112093 -84 112127
rect 84 112093 100 112127
rect -100 112077 100 112093
rect -100 112019 100 112035
rect -100 111985 -84 112019
rect 84 111985 100 112019
rect -100 111947 100 111985
rect -100 110909 100 110947
rect -100 110875 -84 110909
rect 84 110875 100 110909
rect -100 110859 100 110875
rect -100 110801 100 110817
rect -100 110767 -84 110801
rect 84 110767 100 110801
rect -100 110729 100 110767
rect -100 109691 100 109729
rect -100 109657 -84 109691
rect 84 109657 100 109691
rect -100 109641 100 109657
rect -100 109583 100 109599
rect -100 109549 -84 109583
rect 84 109549 100 109583
rect -100 109511 100 109549
rect -100 108473 100 108511
rect -100 108439 -84 108473
rect 84 108439 100 108473
rect -100 108423 100 108439
rect -100 108365 100 108381
rect -100 108331 -84 108365
rect 84 108331 100 108365
rect -100 108293 100 108331
rect -100 107255 100 107293
rect -100 107221 -84 107255
rect 84 107221 100 107255
rect -100 107205 100 107221
rect -100 107147 100 107163
rect -100 107113 -84 107147
rect 84 107113 100 107147
rect -100 107075 100 107113
rect -100 106037 100 106075
rect -100 106003 -84 106037
rect 84 106003 100 106037
rect -100 105987 100 106003
rect -100 105929 100 105945
rect -100 105895 -84 105929
rect 84 105895 100 105929
rect -100 105857 100 105895
rect -100 104819 100 104857
rect -100 104785 -84 104819
rect 84 104785 100 104819
rect -100 104769 100 104785
rect -100 104711 100 104727
rect -100 104677 -84 104711
rect 84 104677 100 104711
rect -100 104639 100 104677
rect -100 103601 100 103639
rect -100 103567 -84 103601
rect 84 103567 100 103601
rect -100 103551 100 103567
rect -100 103493 100 103509
rect -100 103459 -84 103493
rect 84 103459 100 103493
rect -100 103421 100 103459
rect -100 102383 100 102421
rect -100 102349 -84 102383
rect 84 102349 100 102383
rect -100 102333 100 102349
rect -100 102275 100 102291
rect -100 102241 -84 102275
rect 84 102241 100 102275
rect -100 102203 100 102241
rect -100 101165 100 101203
rect -100 101131 -84 101165
rect 84 101131 100 101165
rect -100 101115 100 101131
rect -100 101057 100 101073
rect -100 101023 -84 101057
rect 84 101023 100 101057
rect -100 100985 100 101023
rect -100 99947 100 99985
rect -100 99913 -84 99947
rect 84 99913 100 99947
rect -100 99897 100 99913
rect -100 99839 100 99855
rect -100 99805 -84 99839
rect 84 99805 100 99839
rect -100 99767 100 99805
rect -100 98729 100 98767
rect -100 98695 -84 98729
rect 84 98695 100 98729
rect -100 98679 100 98695
rect -100 98621 100 98637
rect -100 98587 -84 98621
rect 84 98587 100 98621
rect -100 98549 100 98587
rect -100 97511 100 97549
rect -100 97477 -84 97511
rect 84 97477 100 97511
rect -100 97461 100 97477
rect -100 97403 100 97419
rect -100 97369 -84 97403
rect 84 97369 100 97403
rect -100 97331 100 97369
rect -100 96293 100 96331
rect -100 96259 -84 96293
rect 84 96259 100 96293
rect -100 96243 100 96259
rect -100 96185 100 96201
rect -100 96151 -84 96185
rect 84 96151 100 96185
rect -100 96113 100 96151
rect -100 95075 100 95113
rect -100 95041 -84 95075
rect 84 95041 100 95075
rect -100 95025 100 95041
rect -100 94967 100 94983
rect -100 94933 -84 94967
rect 84 94933 100 94967
rect -100 94895 100 94933
rect -100 93857 100 93895
rect -100 93823 -84 93857
rect 84 93823 100 93857
rect -100 93807 100 93823
rect -100 93749 100 93765
rect -100 93715 -84 93749
rect 84 93715 100 93749
rect -100 93677 100 93715
rect -100 92639 100 92677
rect -100 92605 -84 92639
rect 84 92605 100 92639
rect -100 92589 100 92605
rect -100 92531 100 92547
rect -100 92497 -84 92531
rect 84 92497 100 92531
rect -100 92459 100 92497
rect -100 91421 100 91459
rect -100 91387 -84 91421
rect 84 91387 100 91421
rect -100 91371 100 91387
rect -100 91313 100 91329
rect -100 91279 -84 91313
rect 84 91279 100 91313
rect -100 91241 100 91279
rect -100 90203 100 90241
rect -100 90169 -84 90203
rect 84 90169 100 90203
rect -100 90153 100 90169
rect -100 90095 100 90111
rect -100 90061 -84 90095
rect 84 90061 100 90095
rect -100 90023 100 90061
rect -100 88985 100 89023
rect -100 88951 -84 88985
rect 84 88951 100 88985
rect -100 88935 100 88951
rect -100 88877 100 88893
rect -100 88843 -84 88877
rect 84 88843 100 88877
rect -100 88805 100 88843
rect -100 87767 100 87805
rect -100 87733 -84 87767
rect 84 87733 100 87767
rect -100 87717 100 87733
rect -100 87659 100 87675
rect -100 87625 -84 87659
rect 84 87625 100 87659
rect -100 87587 100 87625
rect -100 86549 100 86587
rect -100 86515 -84 86549
rect 84 86515 100 86549
rect -100 86499 100 86515
rect -100 86441 100 86457
rect -100 86407 -84 86441
rect 84 86407 100 86441
rect -100 86369 100 86407
rect -100 85331 100 85369
rect -100 85297 -84 85331
rect 84 85297 100 85331
rect -100 85281 100 85297
rect -100 85223 100 85239
rect -100 85189 -84 85223
rect 84 85189 100 85223
rect -100 85151 100 85189
rect -100 84113 100 84151
rect -100 84079 -84 84113
rect 84 84079 100 84113
rect -100 84063 100 84079
rect -100 84005 100 84021
rect -100 83971 -84 84005
rect 84 83971 100 84005
rect -100 83933 100 83971
rect -100 82895 100 82933
rect -100 82861 -84 82895
rect 84 82861 100 82895
rect -100 82845 100 82861
rect -100 82787 100 82803
rect -100 82753 -84 82787
rect 84 82753 100 82787
rect -100 82715 100 82753
rect -100 81677 100 81715
rect -100 81643 -84 81677
rect 84 81643 100 81677
rect -100 81627 100 81643
rect -100 81569 100 81585
rect -100 81535 -84 81569
rect 84 81535 100 81569
rect -100 81497 100 81535
rect -100 80459 100 80497
rect -100 80425 -84 80459
rect 84 80425 100 80459
rect -100 80409 100 80425
rect -100 80351 100 80367
rect -100 80317 -84 80351
rect 84 80317 100 80351
rect -100 80279 100 80317
rect -100 79241 100 79279
rect -100 79207 -84 79241
rect 84 79207 100 79241
rect -100 79191 100 79207
rect -100 79133 100 79149
rect -100 79099 -84 79133
rect 84 79099 100 79133
rect -100 79061 100 79099
rect -100 78023 100 78061
rect -100 77989 -84 78023
rect 84 77989 100 78023
rect -100 77973 100 77989
rect -100 77915 100 77931
rect -100 77881 -84 77915
rect 84 77881 100 77915
rect -100 77843 100 77881
rect -100 76805 100 76843
rect -100 76771 -84 76805
rect 84 76771 100 76805
rect -100 76755 100 76771
rect -100 76697 100 76713
rect -100 76663 -84 76697
rect 84 76663 100 76697
rect -100 76625 100 76663
rect -100 75587 100 75625
rect -100 75553 -84 75587
rect 84 75553 100 75587
rect -100 75537 100 75553
rect -100 75479 100 75495
rect -100 75445 -84 75479
rect 84 75445 100 75479
rect -100 75407 100 75445
rect -100 74369 100 74407
rect -100 74335 -84 74369
rect 84 74335 100 74369
rect -100 74319 100 74335
rect -100 74261 100 74277
rect -100 74227 -84 74261
rect 84 74227 100 74261
rect -100 74189 100 74227
rect -100 73151 100 73189
rect -100 73117 -84 73151
rect 84 73117 100 73151
rect -100 73101 100 73117
rect -100 73043 100 73059
rect -100 73009 -84 73043
rect 84 73009 100 73043
rect -100 72971 100 73009
rect -100 71933 100 71971
rect -100 71899 -84 71933
rect 84 71899 100 71933
rect -100 71883 100 71899
rect -100 71825 100 71841
rect -100 71791 -84 71825
rect 84 71791 100 71825
rect -100 71753 100 71791
rect -100 70715 100 70753
rect -100 70681 -84 70715
rect 84 70681 100 70715
rect -100 70665 100 70681
rect -100 70607 100 70623
rect -100 70573 -84 70607
rect 84 70573 100 70607
rect -100 70535 100 70573
rect -100 69497 100 69535
rect -100 69463 -84 69497
rect 84 69463 100 69497
rect -100 69447 100 69463
rect -100 69389 100 69405
rect -100 69355 -84 69389
rect 84 69355 100 69389
rect -100 69317 100 69355
rect -100 68279 100 68317
rect -100 68245 -84 68279
rect 84 68245 100 68279
rect -100 68229 100 68245
rect -100 68171 100 68187
rect -100 68137 -84 68171
rect 84 68137 100 68171
rect -100 68099 100 68137
rect -100 67061 100 67099
rect -100 67027 -84 67061
rect 84 67027 100 67061
rect -100 67011 100 67027
rect -100 66953 100 66969
rect -100 66919 -84 66953
rect 84 66919 100 66953
rect -100 66881 100 66919
rect -100 65843 100 65881
rect -100 65809 -84 65843
rect 84 65809 100 65843
rect -100 65793 100 65809
rect -100 65735 100 65751
rect -100 65701 -84 65735
rect 84 65701 100 65735
rect -100 65663 100 65701
rect -100 64625 100 64663
rect -100 64591 -84 64625
rect 84 64591 100 64625
rect -100 64575 100 64591
rect -100 64517 100 64533
rect -100 64483 -84 64517
rect 84 64483 100 64517
rect -100 64445 100 64483
rect -100 63407 100 63445
rect -100 63373 -84 63407
rect 84 63373 100 63407
rect -100 63357 100 63373
rect -100 63299 100 63315
rect -100 63265 -84 63299
rect 84 63265 100 63299
rect -100 63227 100 63265
rect -100 62189 100 62227
rect -100 62155 -84 62189
rect 84 62155 100 62189
rect -100 62139 100 62155
rect -100 62081 100 62097
rect -100 62047 -84 62081
rect 84 62047 100 62081
rect -100 62009 100 62047
rect -100 60971 100 61009
rect -100 60937 -84 60971
rect 84 60937 100 60971
rect -100 60921 100 60937
rect -100 60863 100 60879
rect -100 60829 -84 60863
rect 84 60829 100 60863
rect -100 60791 100 60829
rect -100 59753 100 59791
rect -100 59719 -84 59753
rect 84 59719 100 59753
rect -100 59703 100 59719
rect -100 59645 100 59661
rect -100 59611 -84 59645
rect 84 59611 100 59645
rect -100 59573 100 59611
rect -100 58535 100 58573
rect -100 58501 -84 58535
rect 84 58501 100 58535
rect -100 58485 100 58501
rect -100 58427 100 58443
rect -100 58393 -84 58427
rect 84 58393 100 58427
rect -100 58355 100 58393
rect -100 57317 100 57355
rect -100 57283 -84 57317
rect 84 57283 100 57317
rect -100 57267 100 57283
rect -100 57209 100 57225
rect -100 57175 -84 57209
rect 84 57175 100 57209
rect -100 57137 100 57175
rect -100 56099 100 56137
rect -100 56065 -84 56099
rect 84 56065 100 56099
rect -100 56049 100 56065
rect -100 55991 100 56007
rect -100 55957 -84 55991
rect 84 55957 100 55991
rect -100 55919 100 55957
rect -100 54881 100 54919
rect -100 54847 -84 54881
rect 84 54847 100 54881
rect -100 54831 100 54847
rect -100 54773 100 54789
rect -100 54739 -84 54773
rect 84 54739 100 54773
rect -100 54701 100 54739
rect -100 53663 100 53701
rect -100 53629 -84 53663
rect 84 53629 100 53663
rect -100 53613 100 53629
rect -100 53555 100 53571
rect -100 53521 -84 53555
rect 84 53521 100 53555
rect -100 53483 100 53521
rect -100 52445 100 52483
rect -100 52411 -84 52445
rect 84 52411 100 52445
rect -100 52395 100 52411
rect -100 52337 100 52353
rect -100 52303 -84 52337
rect 84 52303 100 52337
rect -100 52265 100 52303
rect -100 51227 100 51265
rect -100 51193 -84 51227
rect 84 51193 100 51227
rect -100 51177 100 51193
rect -100 51119 100 51135
rect -100 51085 -84 51119
rect 84 51085 100 51119
rect -100 51047 100 51085
rect -100 50009 100 50047
rect -100 49975 -84 50009
rect 84 49975 100 50009
rect -100 49959 100 49975
rect -100 49901 100 49917
rect -100 49867 -84 49901
rect 84 49867 100 49901
rect -100 49829 100 49867
rect -100 48791 100 48829
rect -100 48757 -84 48791
rect 84 48757 100 48791
rect -100 48741 100 48757
rect -100 48683 100 48699
rect -100 48649 -84 48683
rect 84 48649 100 48683
rect -100 48611 100 48649
rect -100 47573 100 47611
rect -100 47539 -84 47573
rect 84 47539 100 47573
rect -100 47523 100 47539
rect -100 47465 100 47481
rect -100 47431 -84 47465
rect 84 47431 100 47465
rect -100 47393 100 47431
rect -100 46355 100 46393
rect -100 46321 -84 46355
rect 84 46321 100 46355
rect -100 46305 100 46321
rect -100 46247 100 46263
rect -100 46213 -84 46247
rect 84 46213 100 46247
rect -100 46175 100 46213
rect -100 45137 100 45175
rect -100 45103 -84 45137
rect 84 45103 100 45137
rect -100 45087 100 45103
rect -100 45029 100 45045
rect -100 44995 -84 45029
rect 84 44995 100 45029
rect -100 44957 100 44995
rect -100 43919 100 43957
rect -100 43885 -84 43919
rect 84 43885 100 43919
rect -100 43869 100 43885
rect -100 43811 100 43827
rect -100 43777 -84 43811
rect 84 43777 100 43811
rect -100 43739 100 43777
rect -100 42701 100 42739
rect -100 42667 -84 42701
rect 84 42667 100 42701
rect -100 42651 100 42667
rect -100 42593 100 42609
rect -100 42559 -84 42593
rect 84 42559 100 42593
rect -100 42521 100 42559
rect -100 41483 100 41521
rect -100 41449 -84 41483
rect 84 41449 100 41483
rect -100 41433 100 41449
rect -100 41375 100 41391
rect -100 41341 -84 41375
rect 84 41341 100 41375
rect -100 41303 100 41341
rect -100 40265 100 40303
rect -100 40231 -84 40265
rect 84 40231 100 40265
rect -100 40215 100 40231
rect -100 40157 100 40173
rect -100 40123 -84 40157
rect 84 40123 100 40157
rect -100 40085 100 40123
rect -100 39047 100 39085
rect -100 39013 -84 39047
rect 84 39013 100 39047
rect -100 38997 100 39013
rect -100 38939 100 38955
rect -100 38905 -84 38939
rect 84 38905 100 38939
rect -100 38867 100 38905
rect -100 37829 100 37867
rect -100 37795 -84 37829
rect 84 37795 100 37829
rect -100 37779 100 37795
rect -100 37721 100 37737
rect -100 37687 -84 37721
rect 84 37687 100 37721
rect -100 37649 100 37687
rect -100 36611 100 36649
rect -100 36577 -84 36611
rect 84 36577 100 36611
rect -100 36561 100 36577
rect -100 36503 100 36519
rect -100 36469 -84 36503
rect 84 36469 100 36503
rect -100 36431 100 36469
rect -100 35393 100 35431
rect -100 35359 -84 35393
rect 84 35359 100 35393
rect -100 35343 100 35359
rect -100 35285 100 35301
rect -100 35251 -84 35285
rect 84 35251 100 35285
rect -100 35213 100 35251
rect -100 34175 100 34213
rect -100 34141 -84 34175
rect 84 34141 100 34175
rect -100 34125 100 34141
rect -100 34067 100 34083
rect -100 34033 -84 34067
rect 84 34033 100 34067
rect -100 33995 100 34033
rect -100 32957 100 32995
rect -100 32923 -84 32957
rect 84 32923 100 32957
rect -100 32907 100 32923
rect -100 32849 100 32865
rect -100 32815 -84 32849
rect 84 32815 100 32849
rect -100 32777 100 32815
rect -100 31739 100 31777
rect -100 31705 -84 31739
rect 84 31705 100 31739
rect -100 31689 100 31705
rect -100 31631 100 31647
rect -100 31597 -84 31631
rect 84 31597 100 31631
rect -100 31559 100 31597
rect -100 30521 100 30559
rect -100 30487 -84 30521
rect 84 30487 100 30521
rect -100 30471 100 30487
rect -100 30413 100 30429
rect -100 30379 -84 30413
rect 84 30379 100 30413
rect -100 30341 100 30379
rect -100 29303 100 29341
rect -100 29269 -84 29303
rect 84 29269 100 29303
rect -100 29253 100 29269
rect -100 29195 100 29211
rect -100 29161 -84 29195
rect 84 29161 100 29195
rect -100 29123 100 29161
rect -100 28085 100 28123
rect -100 28051 -84 28085
rect 84 28051 100 28085
rect -100 28035 100 28051
rect -100 27977 100 27993
rect -100 27943 -84 27977
rect 84 27943 100 27977
rect -100 27905 100 27943
rect -100 26867 100 26905
rect -100 26833 -84 26867
rect 84 26833 100 26867
rect -100 26817 100 26833
rect -100 26759 100 26775
rect -100 26725 -84 26759
rect 84 26725 100 26759
rect -100 26687 100 26725
rect -100 25649 100 25687
rect -100 25615 -84 25649
rect 84 25615 100 25649
rect -100 25599 100 25615
rect -100 25541 100 25557
rect -100 25507 -84 25541
rect 84 25507 100 25541
rect -100 25469 100 25507
rect -100 24431 100 24469
rect -100 24397 -84 24431
rect 84 24397 100 24431
rect -100 24381 100 24397
rect -100 24323 100 24339
rect -100 24289 -84 24323
rect 84 24289 100 24323
rect -100 24251 100 24289
rect -100 23213 100 23251
rect -100 23179 -84 23213
rect 84 23179 100 23213
rect -100 23163 100 23179
rect -100 23105 100 23121
rect -100 23071 -84 23105
rect 84 23071 100 23105
rect -100 23033 100 23071
rect -100 21995 100 22033
rect -100 21961 -84 21995
rect 84 21961 100 21995
rect -100 21945 100 21961
rect -100 21887 100 21903
rect -100 21853 -84 21887
rect 84 21853 100 21887
rect -100 21815 100 21853
rect -100 20777 100 20815
rect -100 20743 -84 20777
rect 84 20743 100 20777
rect -100 20727 100 20743
rect -100 20669 100 20685
rect -100 20635 -84 20669
rect 84 20635 100 20669
rect -100 20597 100 20635
rect -100 19559 100 19597
rect -100 19525 -84 19559
rect 84 19525 100 19559
rect -100 19509 100 19525
rect -100 19451 100 19467
rect -100 19417 -84 19451
rect 84 19417 100 19451
rect -100 19379 100 19417
rect -100 18341 100 18379
rect -100 18307 -84 18341
rect 84 18307 100 18341
rect -100 18291 100 18307
rect -100 18233 100 18249
rect -100 18199 -84 18233
rect 84 18199 100 18233
rect -100 18161 100 18199
rect -100 17123 100 17161
rect -100 17089 -84 17123
rect 84 17089 100 17123
rect -100 17073 100 17089
rect -100 17015 100 17031
rect -100 16981 -84 17015
rect 84 16981 100 17015
rect -100 16943 100 16981
rect -100 15905 100 15943
rect -100 15871 -84 15905
rect 84 15871 100 15905
rect -100 15855 100 15871
rect -100 15797 100 15813
rect -100 15763 -84 15797
rect 84 15763 100 15797
rect -100 15725 100 15763
rect -100 14687 100 14725
rect -100 14653 -84 14687
rect 84 14653 100 14687
rect -100 14637 100 14653
rect -100 14579 100 14595
rect -100 14545 -84 14579
rect 84 14545 100 14579
rect -100 14507 100 14545
rect -100 13469 100 13507
rect -100 13435 -84 13469
rect 84 13435 100 13469
rect -100 13419 100 13435
rect -100 13361 100 13377
rect -100 13327 -84 13361
rect 84 13327 100 13361
rect -100 13289 100 13327
rect -100 12251 100 12289
rect -100 12217 -84 12251
rect 84 12217 100 12251
rect -100 12201 100 12217
rect -100 12143 100 12159
rect -100 12109 -84 12143
rect 84 12109 100 12143
rect -100 12071 100 12109
rect -100 11033 100 11071
rect -100 10999 -84 11033
rect 84 10999 100 11033
rect -100 10983 100 10999
rect -100 10925 100 10941
rect -100 10891 -84 10925
rect 84 10891 100 10925
rect -100 10853 100 10891
rect -100 9815 100 9853
rect -100 9781 -84 9815
rect 84 9781 100 9815
rect -100 9765 100 9781
rect -100 9707 100 9723
rect -100 9673 -84 9707
rect 84 9673 100 9707
rect -100 9635 100 9673
rect -100 8597 100 8635
rect -100 8563 -84 8597
rect 84 8563 100 8597
rect -100 8547 100 8563
rect -100 8489 100 8505
rect -100 8455 -84 8489
rect 84 8455 100 8489
rect -100 8417 100 8455
rect -100 7379 100 7417
rect -100 7345 -84 7379
rect 84 7345 100 7379
rect -100 7329 100 7345
rect -100 7271 100 7287
rect -100 7237 -84 7271
rect 84 7237 100 7271
rect -100 7199 100 7237
rect -100 6161 100 6199
rect -100 6127 -84 6161
rect 84 6127 100 6161
rect -100 6111 100 6127
rect -100 6053 100 6069
rect -100 6019 -84 6053
rect 84 6019 100 6053
rect -100 5981 100 6019
rect -100 4943 100 4981
rect -100 4909 -84 4943
rect 84 4909 100 4943
rect -100 4893 100 4909
rect -100 4835 100 4851
rect -100 4801 -84 4835
rect 84 4801 100 4835
rect -100 4763 100 4801
rect -100 3725 100 3763
rect -100 3691 -84 3725
rect 84 3691 100 3725
rect -100 3675 100 3691
rect -100 3617 100 3633
rect -100 3583 -84 3617
rect 84 3583 100 3617
rect -100 3545 100 3583
rect -100 2507 100 2545
rect -100 2473 -84 2507
rect 84 2473 100 2507
rect -100 2457 100 2473
rect -100 2399 100 2415
rect -100 2365 -84 2399
rect 84 2365 100 2399
rect -100 2327 100 2365
rect -100 1289 100 1327
rect -100 1255 -84 1289
rect 84 1255 100 1289
rect -100 1239 100 1255
rect -100 1181 100 1197
rect -100 1147 -84 1181
rect 84 1147 100 1181
rect -100 1109 100 1147
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect -100 -1147 100 -1109
rect -100 -1181 -84 -1147
rect 84 -1181 100 -1147
rect -100 -1197 100 -1181
rect -100 -1255 100 -1239
rect -100 -1289 -84 -1255
rect 84 -1289 100 -1255
rect -100 -1327 100 -1289
rect -100 -2365 100 -2327
rect -100 -2399 -84 -2365
rect 84 -2399 100 -2365
rect -100 -2415 100 -2399
rect -100 -2473 100 -2457
rect -100 -2507 -84 -2473
rect 84 -2507 100 -2473
rect -100 -2545 100 -2507
rect -100 -3583 100 -3545
rect -100 -3617 -84 -3583
rect 84 -3617 100 -3583
rect -100 -3633 100 -3617
rect -100 -3691 100 -3675
rect -100 -3725 -84 -3691
rect 84 -3725 100 -3691
rect -100 -3763 100 -3725
rect -100 -4801 100 -4763
rect -100 -4835 -84 -4801
rect 84 -4835 100 -4801
rect -100 -4851 100 -4835
rect -100 -4909 100 -4893
rect -100 -4943 -84 -4909
rect 84 -4943 100 -4909
rect -100 -4981 100 -4943
rect -100 -6019 100 -5981
rect -100 -6053 -84 -6019
rect 84 -6053 100 -6019
rect -100 -6069 100 -6053
rect -100 -6127 100 -6111
rect -100 -6161 -84 -6127
rect 84 -6161 100 -6127
rect -100 -6199 100 -6161
rect -100 -7237 100 -7199
rect -100 -7271 -84 -7237
rect 84 -7271 100 -7237
rect -100 -7287 100 -7271
rect -100 -7345 100 -7329
rect -100 -7379 -84 -7345
rect 84 -7379 100 -7345
rect -100 -7417 100 -7379
rect -100 -8455 100 -8417
rect -100 -8489 -84 -8455
rect 84 -8489 100 -8455
rect -100 -8505 100 -8489
rect -100 -8563 100 -8547
rect -100 -8597 -84 -8563
rect 84 -8597 100 -8563
rect -100 -8635 100 -8597
rect -100 -9673 100 -9635
rect -100 -9707 -84 -9673
rect 84 -9707 100 -9673
rect -100 -9723 100 -9707
rect -100 -9781 100 -9765
rect -100 -9815 -84 -9781
rect 84 -9815 100 -9781
rect -100 -9853 100 -9815
rect -100 -10891 100 -10853
rect -100 -10925 -84 -10891
rect 84 -10925 100 -10891
rect -100 -10941 100 -10925
rect -100 -10999 100 -10983
rect -100 -11033 -84 -10999
rect 84 -11033 100 -10999
rect -100 -11071 100 -11033
rect -100 -12109 100 -12071
rect -100 -12143 -84 -12109
rect 84 -12143 100 -12109
rect -100 -12159 100 -12143
rect -100 -12217 100 -12201
rect -100 -12251 -84 -12217
rect 84 -12251 100 -12217
rect -100 -12289 100 -12251
rect -100 -13327 100 -13289
rect -100 -13361 -84 -13327
rect 84 -13361 100 -13327
rect -100 -13377 100 -13361
rect -100 -13435 100 -13419
rect -100 -13469 -84 -13435
rect 84 -13469 100 -13435
rect -100 -13507 100 -13469
rect -100 -14545 100 -14507
rect -100 -14579 -84 -14545
rect 84 -14579 100 -14545
rect -100 -14595 100 -14579
rect -100 -14653 100 -14637
rect -100 -14687 -84 -14653
rect 84 -14687 100 -14653
rect -100 -14725 100 -14687
rect -100 -15763 100 -15725
rect -100 -15797 -84 -15763
rect 84 -15797 100 -15763
rect -100 -15813 100 -15797
rect -100 -15871 100 -15855
rect -100 -15905 -84 -15871
rect 84 -15905 100 -15871
rect -100 -15943 100 -15905
rect -100 -16981 100 -16943
rect -100 -17015 -84 -16981
rect 84 -17015 100 -16981
rect -100 -17031 100 -17015
rect -100 -17089 100 -17073
rect -100 -17123 -84 -17089
rect 84 -17123 100 -17089
rect -100 -17161 100 -17123
rect -100 -18199 100 -18161
rect -100 -18233 -84 -18199
rect 84 -18233 100 -18199
rect -100 -18249 100 -18233
rect -100 -18307 100 -18291
rect -100 -18341 -84 -18307
rect 84 -18341 100 -18307
rect -100 -18379 100 -18341
rect -100 -19417 100 -19379
rect -100 -19451 -84 -19417
rect 84 -19451 100 -19417
rect -100 -19467 100 -19451
rect -100 -19525 100 -19509
rect -100 -19559 -84 -19525
rect 84 -19559 100 -19525
rect -100 -19597 100 -19559
rect -100 -20635 100 -20597
rect -100 -20669 -84 -20635
rect 84 -20669 100 -20635
rect -100 -20685 100 -20669
rect -100 -20743 100 -20727
rect -100 -20777 -84 -20743
rect 84 -20777 100 -20743
rect -100 -20815 100 -20777
rect -100 -21853 100 -21815
rect -100 -21887 -84 -21853
rect 84 -21887 100 -21853
rect -100 -21903 100 -21887
rect -100 -21961 100 -21945
rect -100 -21995 -84 -21961
rect 84 -21995 100 -21961
rect -100 -22033 100 -21995
rect -100 -23071 100 -23033
rect -100 -23105 -84 -23071
rect 84 -23105 100 -23071
rect -100 -23121 100 -23105
rect -100 -23179 100 -23163
rect -100 -23213 -84 -23179
rect 84 -23213 100 -23179
rect -100 -23251 100 -23213
rect -100 -24289 100 -24251
rect -100 -24323 -84 -24289
rect 84 -24323 100 -24289
rect -100 -24339 100 -24323
rect -100 -24397 100 -24381
rect -100 -24431 -84 -24397
rect 84 -24431 100 -24397
rect -100 -24469 100 -24431
rect -100 -25507 100 -25469
rect -100 -25541 -84 -25507
rect 84 -25541 100 -25507
rect -100 -25557 100 -25541
rect -100 -25615 100 -25599
rect -100 -25649 -84 -25615
rect 84 -25649 100 -25615
rect -100 -25687 100 -25649
rect -100 -26725 100 -26687
rect -100 -26759 -84 -26725
rect 84 -26759 100 -26725
rect -100 -26775 100 -26759
rect -100 -26833 100 -26817
rect -100 -26867 -84 -26833
rect 84 -26867 100 -26833
rect -100 -26905 100 -26867
rect -100 -27943 100 -27905
rect -100 -27977 -84 -27943
rect 84 -27977 100 -27943
rect -100 -27993 100 -27977
rect -100 -28051 100 -28035
rect -100 -28085 -84 -28051
rect 84 -28085 100 -28051
rect -100 -28123 100 -28085
rect -100 -29161 100 -29123
rect -100 -29195 -84 -29161
rect 84 -29195 100 -29161
rect -100 -29211 100 -29195
rect -100 -29269 100 -29253
rect -100 -29303 -84 -29269
rect 84 -29303 100 -29269
rect -100 -29341 100 -29303
rect -100 -30379 100 -30341
rect -100 -30413 -84 -30379
rect 84 -30413 100 -30379
rect -100 -30429 100 -30413
rect -100 -30487 100 -30471
rect -100 -30521 -84 -30487
rect 84 -30521 100 -30487
rect -100 -30559 100 -30521
rect -100 -31597 100 -31559
rect -100 -31631 -84 -31597
rect 84 -31631 100 -31597
rect -100 -31647 100 -31631
rect -100 -31705 100 -31689
rect -100 -31739 -84 -31705
rect 84 -31739 100 -31705
rect -100 -31777 100 -31739
rect -100 -32815 100 -32777
rect -100 -32849 -84 -32815
rect 84 -32849 100 -32815
rect -100 -32865 100 -32849
rect -100 -32923 100 -32907
rect -100 -32957 -84 -32923
rect 84 -32957 100 -32923
rect -100 -32995 100 -32957
rect -100 -34033 100 -33995
rect -100 -34067 -84 -34033
rect 84 -34067 100 -34033
rect -100 -34083 100 -34067
rect -100 -34141 100 -34125
rect -100 -34175 -84 -34141
rect 84 -34175 100 -34141
rect -100 -34213 100 -34175
rect -100 -35251 100 -35213
rect -100 -35285 -84 -35251
rect 84 -35285 100 -35251
rect -100 -35301 100 -35285
rect -100 -35359 100 -35343
rect -100 -35393 -84 -35359
rect 84 -35393 100 -35359
rect -100 -35431 100 -35393
rect -100 -36469 100 -36431
rect -100 -36503 -84 -36469
rect 84 -36503 100 -36469
rect -100 -36519 100 -36503
rect -100 -36577 100 -36561
rect -100 -36611 -84 -36577
rect 84 -36611 100 -36577
rect -100 -36649 100 -36611
rect -100 -37687 100 -37649
rect -100 -37721 -84 -37687
rect 84 -37721 100 -37687
rect -100 -37737 100 -37721
rect -100 -37795 100 -37779
rect -100 -37829 -84 -37795
rect 84 -37829 100 -37795
rect -100 -37867 100 -37829
rect -100 -38905 100 -38867
rect -100 -38939 -84 -38905
rect 84 -38939 100 -38905
rect -100 -38955 100 -38939
rect -100 -39013 100 -38997
rect -100 -39047 -84 -39013
rect 84 -39047 100 -39013
rect -100 -39085 100 -39047
rect -100 -40123 100 -40085
rect -100 -40157 -84 -40123
rect 84 -40157 100 -40123
rect -100 -40173 100 -40157
rect -100 -40231 100 -40215
rect -100 -40265 -84 -40231
rect 84 -40265 100 -40231
rect -100 -40303 100 -40265
rect -100 -41341 100 -41303
rect -100 -41375 -84 -41341
rect 84 -41375 100 -41341
rect -100 -41391 100 -41375
rect -100 -41449 100 -41433
rect -100 -41483 -84 -41449
rect 84 -41483 100 -41449
rect -100 -41521 100 -41483
rect -100 -42559 100 -42521
rect -100 -42593 -84 -42559
rect 84 -42593 100 -42559
rect -100 -42609 100 -42593
rect -100 -42667 100 -42651
rect -100 -42701 -84 -42667
rect 84 -42701 100 -42667
rect -100 -42739 100 -42701
rect -100 -43777 100 -43739
rect -100 -43811 -84 -43777
rect 84 -43811 100 -43777
rect -100 -43827 100 -43811
rect -100 -43885 100 -43869
rect -100 -43919 -84 -43885
rect 84 -43919 100 -43885
rect -100 -43957 100 -43919
rect -100 -44995 100 -44957
rect -100 -45029 -84 -44995
rect 84 -45029 100 -44995
rect -100 -45045 100 -45029
rect -100 -45103 100 -45087
rect -100 -45137 -84 -45103
rect 84 -45137 100 -45103
rect -100 -45175 100 -45137
rect -100 -46213 100 -46175
rect -100 -46247 -84 -46213
rect 84 -46247 100 -46213
rect -100 -46263 100 -46247
rect -100 -46321 100 -46305
rect -100 -46355 -84 -46321
rect 84 -46355 100 -46321
rect -100 -46393 100 -46355
rect -100 -47431 100 -47393
rect -100 -47465 -84 -47431
rect 84 -47465 100 -47431
rect -100 -47481 100 -47465
rect -100 -47539 100 -47523
rect -100 -47573 -84 -47539
rect 84 -47573 100 -47539
rect -100 -47611 100 -47573
rect -100 -48649 100 -48611
rect -100 -48683 -84 -48649
rect 84 -48683 100 -48649
rect -100 -48699 100 -48683
rect -100 -48757 100 -48741
rect -100 -48791 -84 -48757
rect 84 -48791 100 -48757
rect -100 -48829 100 -48791
rect -100 -49867 100 -49829
rect -100 -49901 -84 -49867
rect 84 -49901 100 -49867
rect -100 -49917 100 -49901
rect -100 -49975 100 -49959
rect -100 -50009 -84 -49975
rect 84 -50009 100 -49975
rect -100 -50047 100 -50009
rect -100 -51085 100 -51047
rect -100 -51119 -84 -51085
rect 84 -51119 100 -51085
rect -100 -51135 100 -51119
rect -100 -51193 100 -51177
rect -100 -51227 -84 -51193
rect 84 -51227 100 -51193
rect -100 -51265 100 -51227
rect -100 -52303 100 -52265
rect -100 -52337 -84 -52303
rect 84 -52337 100 -52303
rect -100 -52353 100 -52337
rect -100 -52411 100 -52395
rect -100 -52445 -84 -52411
rect 84 -52445 100 -52411
rect -100 -52483 100 -52445
rect -100 -53521 100 -53483
rect -100 -53555 -84 -53521
rect 84 -53555 100 -53521
rect -100 -53571 100 -53555
rect -100 -53629 100 -53613
rect -100 -53663 -84 -53629
rect 84 -53663 100 -53629
rect -100 -53701 100 -53663
rect -100 -54739 100 -54701
rect -100 -54773 -84 -54739
rect 84 -54773 100 -54739
rect -100 -54789 100 -54773
rect -100 -54847 100 -54831
rect -100 -54881 -84 -54847
rect 84 -54881 100 -54847
rect -100 -54919 100 -54881
rect -100 -55957 100 -55919
rect -100 -55991 -84 -55957
rect 84 -55991 100 -55957
rect -100 -56007 100 -55991
rect -100 -56065 100 -56049
rect -100 -56099 -84 -56065
rect 84 -56099 100 -56065
rect -100 -56137 100 -56099
rect -100 -57175 100 -57137
rect -100 -57209 -84 -57175
rect 84 -57209 100 -57175
rect -100 -57225 100 -57209
rect -100 -57283 100 -57267
rect -100 -57317 -84 -57283
rect 84 -57317 100 -57283
rect -100 -57355 100 -57317
rect -100 -58393 100 -58355
rect -100 -58427 -84 -58393
rect 84 -58427 100 -58393
rect -100 -58443 100 -58427
rect -100 -58501 100 -58485
rect -100 -58535 -84 -58501
rect 84 -58535 100 -58501
rect -100 -58573 100 -58535
rect -100 -59611 100 -59573
rect -100 -59645 -84 -59611
rect 84 -59645 100 -59611
rect -100 -59661 100 -59645
rect -100 -59719 100 -59703
rect -100 -59753 -84 -59719
rect 84 -59753 100 -59719
rect -100 -59791 100 -59753
rect -100 -60829 100 -60791
rect -100 -60863 -84 -60829
rect 84 -60863 100 -60829
rect -100 -60879 100 -60863
rect -100 -60937 100 -60921
rect -100 -60971 -84 -60937
rect 84 -60971 100 -60937
rect -100 -61009 100 -60971
rect -100 -62047 100 -62009
rect -100 -62081 -84 -62047
rect 84 -62081 100 -62047
rect -100 -62097 100 -62081
rect -100 -62155 100 -62139
rect -100 -62189 -84 -62155
rect 84 -62189 100 -62155
rect -100 -62227 100 -62189
rect -100 -63265 100 -63227
rect -100 -63299 -84 -63265
rect 84 -63299 100 -63265
rect -100 -63315 100 -63299
rect -100 -63373 100 -63357
rect -100 -63407 -84 -63373
rect 84 -63407 100 -63373
rect -100 -63445 100 -63407
rect -100 -64483 100 -64445
rect -100 -64517 -84 -64483
rect 84 -64517 100 -64483
rect -100 -64533 100 -64517
rect -100 -64591 100 -64575
rect -100 -64625 -84 -64591
rect 84 -64625 100 -64591
rect -100 -64663 100 -64625
rect -100 -65701 100 -65663
rect -100 -65735 -84 -65701
rect 84 -65735 100 -65701
rect -100 -65751 100 -65735
rect -100 -65809 100 -65793
rect -100 -65843 -84 -65809
rect 84 -65843 100 -65809
rect -100 -65881 100 -65843
rect -100 -66919 100 -66881
rect -100 -66953 -84 -66919
rect 84 -66953 100 -66919
rect -100 -66969 100 -66953
rect -100 -67027 100 -67011
rect -100 -67061 -84 -67027
rect 84 -67061 100 -67027
rect -100 -67099 100 -67061
rect -100 -68137 100 -68099
rect -100 -68171 -84 -68137
rect 84 -68171 100 -68137
rect -100 -68187 100 -68171
rect -100 -68245 100 -68229
rect -100 -68279 -84 -68245
rect 84 -68279 100 -68245
rect -100 -68317 100 -68279
rect -100 -69355 100 -69317
rect -100 -69389 -84 -69355
rect 84 -69389 100 -69355
rect -100 -69405 100 -69389
rect -100 -69463 100 -69447
rect -100 -69497 -84 -69463
rect 84 -69497 100 -69463
rect -100 -69535 100 -69497
rect -100 -70573 100 -70535
rect -100 -70607 -84 -70573
rect 84 -70607 100 -70573
rect -100 -70623 100 -70607
rect -100 -70681 100 -70665
rect -100 -70715 -84 -70681
rect 84 -70715 100 -70681
rect -100 -70753 100 -70715
rect -100 -71791 100 -71753
rect -100 -71825 -84 -71791
rect 84 -71825 100 -71791
rect -100 -71841 100 -71825
rect -100 -71899 100 -71883
rect -100 -71933 -84 -71899
rect 84 -71933 100 -71899
rect -100 -71971 100 -71933
rect -100 -73009 100 -72971
rect -100 -73043 -84 -73009
rect 84 -73043 100 -73009
rect -100 -73059 100 -73043
rect -100 -73117 100 -73101
rect -100 -73151 -84 -73117
rect 84 -73151 100 -73117
rect -100 -73189 100 -73151
rect -100 -74227 100 -74189
rect -100 -74261 -84 -74227
rect 84 -74261 100 -74227
rect -100 -74277 100 -74261
rect -100 -74335 100 -74319
rect -100 -74369 -84 -74335
rect 84 -74369 100 -74335
rect -100 -74407 100 -74369
rect -100 -75445 100 -75407
rect -100 -75479 -84 -75445
rect 84 -75479 100 -75445
rect -100 -75495 100 -75479
rect -100 -75553 100 -75537
rect -100 -75587 -84 -75553
rect 84 -75587 100 -75553
rect -100 -75625 100 -75587
rect -100 -76663 100 -76625
rect -100 -76697 -84 -76663
rect 84 -76697 100 -76663
rect -100 -76713 100 -76697
rect -100 -76771 100 -76755
rect -100 -76805 -84 -76771
rect 84 -76805 100 -76771
rect -100 -76843 100 -76805
rect -100 -77881 100 -77843
rect -100 -77915 -84 -77881
rect 84 -77915 100 -77881
rect -100 -77931 100 -77915
rect -100 -77989 100 -77973
rect -100 -78023 -84 -77989
rect 84 -78023 100 -77989
rect -100 -78061 100 -78023
rect -100 -79099 100 -79061
rect -100 -79133 -84 -79099
rect 84 -79133 100 -79099
rect -100 -79149 100 -79133
rect -100 -79207 100 -79191
rect -100 -79241 -84 -79207
rect 84 -79241 100 -79207
rect -100 -79279 100 -79241
rect -100 -80317 100 -80279
rect -100 -80351 -84 -80317
rect 84 -80351 100 -80317
rect -100 -80367 100 -80351
rect -100 -80425 100 -80409
rect -100 -80459 -84 -80425
rect 84 -80459 100 -80425
rect -100 -80497 100 -80459
rect -100 -81535 100 -81497
rect -100 -81569 -84 -81535
rect 84 -81569 100 -81535
rect -100 -81585 100 -81569
rect -100 -81643 100 -81627
rect -100 -81677 -84 -81643
rect 84 -81677 100 -81643
rect -100 -81715 100 -81677
rect -100 -82753 100 -82715
rect -100 -82787 -84 -82753
rect 84 -82787 100 -82753
rect -100 -82803 100 -82787
rect -100 -82861 100 -82845
rect -100 -82895 -84 -82861
rect 84 -82895 100 -82861
rect -100 -82933 100 -82895
rect -100 -83971 100 -83933
rect -100 -84005 -84 -83971
rect 84 -84005 100 -83971
rect -100 -84021 100 -84005
rect -100 -84079 100 -84063
rect -100 -84113 -84 -84079
rect 84 -84113 100 -84079
rect -100 -84151 100 -84113
rect -100 -85189 100 -85151
rect -100 -85223 -84 -85189
rect 84 -85223 100 -85189
rect -100 -85239 100 -85223
rect -100 -85297 100 -85281
rect -100 -85331 -84 -85297
rect 84 -85331 100 -85297
rect -100 -85369 100 -85331
rect -100 -86407 100 -86369
rect -100 -86441 -84 -86407
rect 84 -86441 100 -86407
rect -100 -86457 100 -86441
rect -100 -86515 100 -86499
rect -100 -86549 -84 -86515
rect 84 -86549 100 -86515
rect -100 -86587 100 -86549
rect -100 -87625 100 -87587
rect -100 -87659 -84 -87625
rect 84 -87659 100 -87625
rect -100 -87675 100 -87659
rect -100 -87733 100 -87717
rect -100 -87767 -84 -87733
rect 84 -87767 100 -87733
rect -100 -87805 100 -87767
rect -100 -88843 100 -88805
rect -100 -88877 -84 -88843
rect 84 -88877 100 -88843
rect -100 -88893 100 -88877
rect -100 -88951 100 -88935
rect -100 -88985 -84 -88951
rect 84 -88985 100 -88951
rect -100 -89023 100 -88985
rect -100 -90061 100 -90023
rect -100 -90095 -84 -90061
rect 84 -90095 100 -90061
rect -100 -90111 100 -90095
rect -100 -90169 100 -90153
rect -100 -90203 -84 -90169
rect 84 -90203 100 -90169
rect -100 -90241 100 -90203
rect -100 -91279 100 -91241
rect -100 -91313 -84 -91279
rect 84 -91313 100 -91279
rect -100 -91329 100 -91313
rect -100 -91387 100 -91371
rect -100 -91421 -84 -91387
rect 84 -91421 100 -91387
rect -100 -91459 100 -91421
rect -100 -92497 100 -92459
rect -100 -92531 -84 -92497
rect 84 -92531 100 -92497
rect -100 -92547 100 -92531
rect -100 -92605 100 -92589
rect -100 -92639 -84 -92605
rect 84 -92639 100 -92605
rect -100 -92677 100 -92639
rect -100 -93715 100 -93677
rect -100 -93749 -84 -93715
rect 84 -93749 100 -93715
rect -100 -93765 100 -93749
rect -100 -93823 100 -93807
rect -100 -93857 -84 -93823
rect 84 -93857 100 -93823
rect -100 -93895 100 -93857
rect -100 -94933 100 -94895
rect -100 -94967 -84 -94933
rect 84 -94967 100 -94933
rect -100 -94983 100 -94967
rect -100 -95041 100 -95025
rect -100 -95075 -84 -95041
rect 84 -95075 100 -95041
rect -100 -95113 100 -95075
rect -100 -96151 100 -96113
rect -100 -96185 -84 -96151
rect 84 -96185 100 -96151
rect -100 -96201 100 -96185
rect -100 -96259 100 -96243
rect -100 -96293 -84 -96259
rect 84 -96293 100 -96259
rect -100 -96331 100 -96293
rect -100 -97369 100 -97331
rect -100 -97403 -84 -97369
rect 84 -97403 100 -97369
rect -100 -97419 100 -97403
rect -100 -97477 100 -97461
rect -100 -97511 -84 -97477
rect 84 -97511 100 -97477
rect -100 -97549 100 -97511
rect -100 -98587 100 -98549
rect -100 -98621 -84 -98587
rect 84 -98621 100 -98587
rect -100 -98637 100 -98621
rect -100 -98695 100 -98679
rect -100 -98729 -84 -98695
rect 84 -98729 100 -98695
rect -100 -98767 100 -98729
rect -100 -99805 100 -99767
rect -100 -99839 -84 -99805
rect 84 -99839 100 -99805
rect -100 -99855 100 -99839
rect -100 -99913 100 -99897
rect -100 -99947 -84 -99913
rect 84 -99947 100 -99913
rect -100 -99985 100 -99947
rect -100 -101023 100 -100985
rect -100 -101057 -84 -101023
rect 84 -101057 100 -101023
rect -100 -101073 100 -101057
rect -100 -101131 100 -101115
rect -100 -101165 -84 -101131
rect 84 -101165 100 -101131
rect -100 -101203 100 -101165
rect -100 -102241 100 -102203
rect -100 -102275 -84 -102241
rect 84 -102275 100 -102241
rect -100 -102291 100 -102275
rect -100 -102349 100 -102333
rect -100 -102383 -84 -102349
rect 84 -102383 100 -102349
rect -100 -102421 100 -102383
rect -100 -103459 100 -103421
rect -100 -103493 -84 -103459
rect 84 -103493 100 -103459
rect -100 -103509 100 -103493
rect -100 -103567 100 -103551
rect -100 -103601 -84 -103567
rect 84 -103601 100 -103567
rect -100 -103639 100 -103601
rect -100 -104677 100 -104639
rect -100 -104711 -84 -104677
rect 84 -104711 100 -104677
rect -100 -104727 100 -104711
rect -100 -104785 100 -104769
rect -100 -104819 -84 -104785
rect 84 -104819 100 -104785
rect -100 -104857 100 -104819
rect -100 -105895 100 -105857
rect -100 -105929 -84 -105895
rect 84 -105929 100 -105895
rect -100 -105945 100 -105929
rect -100 -106003 100 -105987
rect -100 -106037 -84 -106003
rect 84 -106037 100 -106003
rect -100 -106075 100 -106037
rect -100 -107113 100 -107075
rect -100 -107147 -84 -107113
rect 84 -107147 100 -107113
rect -100 -107163 100 -107147
rect -100 -107221 100 -107205
rect -100 -107255 -84 -107221
rect 84 -107255 100 -107221
rect -100 -107293 100 -107255
rect -100 -108331 100 -108293
rect -100 -108365 -84 -108331
rect 84 -108365 100 -108331
rect -100 -108381 100 -108365
rect -100 -108439 100 -108423
rect -100 -108473 -84 -108439
rect 84 -108473 100 -108439
rect -100 -108511 100 -108473
rect -100 -109549 100 -109511
rect -100 -109583 -84 -109549
rect 84 -109583 100 -109549
rect -100 -109599 100 -109583
rect -100 -109657 100 -109641
rect -100 -109691 -84 -109657
rect 84 -109691 100 -109657
rect -100 -109729 100 -109691
rect -100 -110767 100 -110729
rect -100 -110801 -84 -110767
rect 84 -110801 100 -110767
rect -100 -110817 100 -110801
rect -100 -110875 100 -110859
rect -100 -110909 -84 -110875
rect 84 -110909 100 -110875
rect -100 -110947 100 -110909
rect -100 -111985 100 -111947
rect -100 -112019 -84 -111985
rect 84 -112019 100 -111985
rect -100 -112035 100 -112019
rect -100 -112093 100 -112077
rect -100 -112127 -84 -112093
rect 84 -112127 100 -112093
rect -100 -112165 100 -112127
rect -100 -113203 100 -113165
rect -100 -113237 -84 -113203
rect 84 -113237 100 -113203
rect -100 -113253 100 -113237
rect -100 -113311 100 -113295
rect -100 -113345 -84 -113311
rect 84 -113345 100 -113311
rect -100 -113383 100 -113345
rect -100 -114421 100 -114383
rect -100 -114455 -84 -114421
rect 84 -114455 100 -114421
rect -100 -114471 100 -114455
rect -100 -114529 100 -114513
rect -100 -114563 -84 -114529
rect 84 -114563 100 -114529
rect -100 -114601 100 -114563
rect -100 -115639 100 -115601
rect -100 -115673 -84 -115639
rect 84 -115673 100 -115639
rect -100 -115689 100 -115673
rect -100 -115747 100 -115731
rect -100 -115781 -84 -115747
rect 84 -115781 100 -115747
rect -100 -115819 100 -115781
rect -100 -116857 100 -116819
rect -100 -116891 -84 -116857
rect 84 -116891 100 -116857
rect -100 -116907 100 -116891
rect -100 -116965 100 -116949
rect -100 -116999 -84 -116965
rect 84 -116999 100 -116965
rect -100 -117037 100 -116999
rect -100 -118075 100 -118037
rect -100 -118109 -84 -118075
rect 84 -118109 100 -118075
rect -100 -118125 100 -118109
rect -100 -118183 100 -118167
rect -100 -118217 -84 -118183
rect 84 -118217 100 -118183
rect -100 -118255 100 -118217
rect -100 -119293 100 -119255
rect -100 -119327 -84 -119293
rect 84 -119327 100 -119293
rect -100 -119343 100 -119327
rect -100 -119401 100 -119385
rect -100 -119435 -84 -119401
rect 84 -119435 100 -119401
rect -100 -119473 100 -119435
rect -100 -120511 100 -120473
rect -100 -120545 -84 -120511
rect 84 -120545 100 -120511
rect -100 -120561 100 -120545
rect -100 -120619 100 -120603
rect -100 -120653 -84 -120619
rect 84 -120653 100 -120619
rect -100 -120691 100 -120653
rect -100 -121729 100 -121691
rect -100 -121763 -84 -121729
rect 84 -121763 100 -121729
rect -100 -121779 100 -121763
<< polycont >>
rect -84 121729 84 121763
rect -84 120619 84 120653
rect -84 120511 84 120545
rect -84 119401 84 119435
rect -84 119293 84 119327
rect -84 118183 84 118217
rect -84 118075 84 118109
rect -84 116965 84 116999
rect -84 116857 84 116891
rect -84 115747 84 115781
rect -84 115639 84 115673
rect -84 114529 84 114563
rect -84 114421 84 114455
rect -84 113311 84 113345
rect -84 113203 84 113237
rect -84 112093 84 112127
rect -84 111985 84 112019
rect -84 110875 84 110909
rect -84 110767 84 110801
rect -84 109657 84 109691
rect -84 109549 84 109583
rect -84 108439 84 108473
rect -84 108331 84 108365
rect -84 107221 84 107255
rect -84 107113 84 107147
rect -84 106003 84 106037
rect -84 105895 84 105929
rect -84 104785 84 104819
rect -84 104677 84 104711
rect -84 103567 84 103601
rect -84 103459 84 103493
rect -84 102349 84 102383
rect -84 102241 84 102275
rect -84 101131 84 101165
rect -84 101023 84 101057
rect -84 99913 84 99947
rect -84 99805 84 99839
rect -84 98695 84 98729
rect -84 98587 84 98621
rect -84 97477 84 97511
rect -84 97369 84 97403
rect -84 96259 84 96293
rect -84 96151 84 96185
rect -84 95041 84 95075
rect -84 94933 84 94967
rect -84 93823 84 93857
rect -84 93715 84 93749
rect -84 92605 84 92639
rect -84 92497 84 92531
rect -84 91387 84 91421
rect -84 91279 84 91313
rect -84 90169 84 90203
rect -84 90061 84 90095
rect -84 88951 84 88985
rect -84 88843 84 88877
rect -84 87733 84 87767
rect -84 87625 84 87659
rect -84 86515 84 86549
rect -84 86407 84 86441
rect -84 85297 84 85331
rect -84 85189 84 85223
rect -84 84079 84 84113
rect -84 83971 84 84005
rect -84 82861 84 82895
rect -84 82753 84 82787
rect -84 81643 84 81677
rect -84 81535 84 81569
rect -84 80425 84 80459
rect -84 80317 84 80351
rect -84 79207 84 79241
rect -84 79099 84 79133
rect -84 77989 84 78023
rect -84 77881 84 77915
rect -84 76771 84 76805
rect -84 76663 84 76697
rect -84 75553 84 75587
rect -84 75445 84 75479
rect -84 74335 84 74369
rect -84 74227 84 74261
rect -84 73117 84 73151
rect -84 73009 84 73043
rect -84 71899 84 71933
rect -84 71791 84 71825
rect -84 70681 84 70715
rect -84 70573 84 70607
rect -84 69463 84 69497
rect -84 69355 84 69389
rect -84 68245 84 68279
rect -84 68137 84 68171
rect -84 67027 84 67061
rect -84 66919 84 66953
rect -84 65809 84 65843
rect -84 65701 84 65735
rect -84 64591 84 64625
rect -84 64483 84 64517
rect -84 63373 84 63407
rect -84 63265 84 63299
rect -84 62155 84 62189
rect -84 62047 84 62081
rect -84 60937 84 60971
rect -84 60829 84 60863
rect -84 59719 84 59753
rect -84 59611 84 59645
rect -84 58501 84 58535
rect -84 58393 84 58427
rect -84 57283 84 57317
rect -84 57175 84 57209
rect -84 56065 84 56099
rect -84 55957 84 55991
rect -84 54847 84 54881
rect -84 54739 84 54773
rect -84 53629 84 53663
rect -84 53521 84 53555
rect -84 52411 84 52445
rect -84 52303 84 52337
rect -84 51193 84 51227
rect -84 51085 84 51119
rect -84 49975 84 50009
rect -84 49867 84 49901
rect -84 48757 84 48791
rect -84 48649 84 48683
rect -84 47539 84 47573
rect -84 47431 84 47465
rect -84 46321 84 46355
rect -84 46213 84 46247
rect -84 45103 84 45137
rect -84 44995 84 45029
rect -84 43885 84 43919
rect -84 43777 84 43811
rect -84 42667 84 42701
rect -84 42559 84 42593
rect -84 41449 84 41483
rect -84 41341 84 41375
rect -84 40231 84 40265
rect -84 40123 84 40157
rect -84 39013 84 39047
rect -84 38905 84 38939
rect -84 37795 84 37829
rect -84 37687 84 37721
rect -84 36577 84 36611
rect -84 36469 84 36503
rect -84 35359 84 35393
rect -84 35251 84 35285
rect -84 34141 84 34175
rect -84 34033 84 34067
rect -84 32923 84 32957
rect -84 32815 84 32849
rect -84 31705 84 31739
rect -84 31597 84 31631
rect -84 30487 84 30521
rect -84 30379 84 30413
rect -84 29269 84 29303
rect -84 29161 84 29195
rect -84 28051 84 28085
rect -84 27943 84 27977
rect -84 26833 84 26867
rect -84 26725 84 26759
rect -84 25615 84 25649
rect -84 25507 84 25541
rect -84 24397 84 24431
rect -84 24289 84 24323
rect -84 23179 84 23213
rect -84 23071 84 23105
rect -84 21961 84 21995
rect -84 21853 84 21887
rect -84 20743 84 20777
rect -84 20635 84 20669
rect -84 19525 84 19559
rect -84 19417 84 19451
rect -84 18307 84 18341
rect -84 18199 84 18233
rect -84 17089 84 17123
rect -84 16981 84 17015
rect -84 15871 84 15905
rect -84 15763 84 15797
rect -84 14653 84 14687
rect -84 14545 84 14579
rect -84 13435 84 13469
rect -84 13327 84 13361
rect -84 12217 84 12251
rect -84 12109 84 12143
rect -84 10999 84 11033
rect -84 10891 84 10925
rect -84 9781 84 9815
rect -84 9673 84 9707
rect -84 8563 84 8597
rect -84 8455 84 8489
rect -84 7345 84 7379
rect -84 7237 84 7271
rect -84 6127 84 6161
rect -84 6019 84 6053
rect -84 4909 84 4943
rect -84 4801 84 4835
rect -84 3691 84 3725
rect -84 3583 84 3617
rect -84 2473 84 2507
rect -84 2365 84 2399
rect -84 1255 84 1289
rect -84 1147 84 1181
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -1181 84 -1147
rect -84 -1289 84 -1255
rect -84 -2399 84 -2365
rect -84 -2507 84 -2473
rect -84 -3617 84 -3583
rect -84 -3725 84 -3691
rect -84 -4835 84 -4801
rect -84 -4943 84 -4909
rect -84 -6053 84 -6019
rect -84 -6161 84 -6127
rect -84 -7271 84 -7237
rect -84 -7379 84 -7345
rect -84 -8489 84 -8455
rect -84 -8597 84 -8563
rect -84 -9707 84 -9673
rect -84 -9815 84 -9781
rect -84 -10925 84 -10891
rect -84 -11033 84 -10999
rect -84 -12143 84 -12109
rect -84 -12251 84 -12217
rect -84 -13361 84 -13327
rect -84 -13469 84 -13435
rect -84 -14579 84 -14545
rect -84 -14687 84 -14653
rect -84 -15797 84 -15763
rect -84 -15905 84 -15871
rect -84 -17015 84 -16981
rect -84 -17123 84 -17089
rect -84 -18233 84 -18199
rect -84 -18341 84 -18307
rect -84 -19451 84 -19417
rect -84 -19559 84 -19525
rect -84 -20669 84 -20635
rect -84 -20777 84 -20743
rect -84 -21887 84 -21853
rect -84 -21995 84 -21961
rect -84 -23105 84 -23071
rect -84 -23213 84 -23179
rect -84 -24323 84 -24289
rect -84 -24431 84 -24397
rect -84 -25541 84 -25507
rect -84 -25649 84 -25615
rect -84 -26759 84 -26725
rect -84 -26867 84 -26833
rect -84 -27977 84 -27943
rect -84 -28085 84 -28051
rect -84 -29195 84 -29161
rect -84 -29303 84 -29269
rect -84 -30413 84 -30379
rect -84 -30521 84 -30487
rect -84 -31631 84 -31597
rect -84 -31739 84 -31705
rect -84 -32849 84 -32815
rect -84 -32957 84 -32923
rect -84 -34067 84 -34033
rect -84 -34175 84 -34141
rect -84 -35285 84 -35251
rect -84 -35393 84 -35359
rect -84 -36503 84 -36469
rect -84 -36611 84 -36577
rect -84 -37721 84 -37687
rect -84 -37829 84 -37795
rect -84 -38939 84 -38905
rect -84 -39047 84 -39013
rect -84 -40157 84 -40123
rect -84 -40265 84 -40231
rect -84 -41375 84 -41341
rect -84 -41483 84 -41449
rect -84 -42593 84 -42559
rect -84 -42701 84 -42667
rect -84 -43811 84 -43777
rect -84 -43919 84 -43885
rect -84 -45029 84 -44995
rect -84 -45137 84 -45103
rect -84 -46247 84 -46213
rect -84 -46355 84 -46321
rect -84 -47465 84 -47431
rect -84 -47573 84 -47539
rect -84 -48683 84 -48649
rect -84 -48791 84 -48757
rect -84 -49901 84 -49867
rect -84 -50009 84 -49975
rect -84 -51119 84 -51085
rect -84 -51227 84 -51193
rect -84 -52337 84 -52303
rect -84 -52445 84 -52411
rect -84 -53555 84 -53521
rect -84 -53663 84 -53629
rect -84 -54773 84 -54739
rect -84 -54881 84 -54847
rect -84 -55991 84 -55957
rect -84 -56099 84 -56065
rect -84 -57209 84 -57175
rect -84 -57317 84 -57283
rect -84 -58427 84 -58393
rect -84 -58535 84 -58501
rect -84 -59645 84 -59611
rect -84 -59753 84 -59719
rect -84 -60863 84 -60829
rect -84 -60971 84 -60937
rect -84 -62081 84 -62047
rect -84 -62189 84 -62155
rect -84 -63299 84 -63265
rect -84 -63407 84 -63373
rect -84 -64517 84 -64483
rect -84 -64625 84 -64591
rect -84 -65735 84 -65701
rect -84 -65843 84 -65809
rect -84 -66953 84 -66919
rect -84 -67061 84 -67027
rect -84 -68171 84 -68137
rect -84 -68279 84 -68245
rect -84 -69389 84 -69355
rect -84 -69497 84 -69463
rect -84 -70607 84 -70573
rect -84 -70715 84 -70681
rect -84 -71825 84 -71791
rect -84 -71933 84 -71899
rect -84 -73043 84 -73009
rect -84 -73151 84 -73117
rect -84 -74261 84 -74227
rect -84 -74369 84 -74335
rect -84 -75479 84 -75445
rect -84 -75587 84 -75553
rect -84 -76697 84 -76663
rect -84 -76805 84 -76771
rect -84 -77915 84 -77881
rect -84 -78023 84 -77989
rect -84 -79133 84 -79099
rect -84 -79241 84 -79207
rect -84 -80351 84 -80317
rect -84 -80459 84 -80425
rect -84 -81569 84 -81535
rect -84 -81677 84 -81643
rect -84 -82787 84 -82753
rect -84 -82895 84 -82861
rect -84 -84005 84 -83971
rect -84 -84113 84 -84079
rect -84 -85223 84 -85189
rect -84 -85331 84 -85297
rect -84 -86441 84 -86407
rect -84 -86549 84 -86515
rect -84 -87659 84 -87625
rect -84 -87767 84 -87733
rect -84 -88877 84 -88843
rect -84 -88985 84 -88951
rect -84 -90095 84 -90061
rect -84 -90203 84 -90169
rect -84 -91313 84 -91279
rect -84 -91421 84 -91387
rect -84 -92531 84 -92497
rect -84 -92639 84 -92605
rect -84 -93749 84 -93715
rect -84 -93857 84 -93823
rect -84 -94967 84 -94933
rect -84 -95075 84 -95041
rect -84 -96185 84 -96151
rect -84 -96293 84 -96259
rect -84 -97403 84 -97369
rect -84 -97511 84 -97477
rect -84 -98621 84 -98587
rect -84 -98729 84 -98695
rect -84 -99839 84 -99805
rect -84 -99947 84 -99913
rect -84 -101057 84 -101023
rect -84 -101165 84 -101131
rect -84 -102275 84 -102241
rect -84 -102383 84 -102349
rect -84 -103493 84 -103459
rect -84 -103601 84 -103567
rect -84 -104711 84 -104677
rect -84 -104819 84 -104785
rect -84 -105929 84 -105895
rect -84 -106037 84 -106003
rect -84 -107147 84 -107113
rect -84 -107255 84 -107221
rect -84 -108365 84 -108331
rect -84 -108473 84 -108439
rect -84 -109583 84 -109549
rect -84 -109691 84 -109657
rect -84 -110801 84 -110767
rect -84 -110909 84 -110875
rect -84 -112019 84 -111985
rect -84 -112127 84 -112093
rect -84 -113237 84 -113203
rect -84 -113345 84 -113311
rect -84 -114455 84 -114421
rect -84 -114563 84 -114529
rect -84 -115673 84 -115639
rect -84 -115781 84 -115747
rect -84 -116891 84 -116857
rect -84 -116999 84 -116965
rect -84 -118109 84 -118075
rect -84 -118217 84 -118183
rect -84 -119327 84 -119293
rect -84 -119435 84 -119401
rect -84 -120545 84 -120511
rect -84 -120653 84 -120619
rect -84 -121763 84 -121729
<< locali >>
rect -280 121867 -184 121901
rect 184 121867 280 121901
rect -280 121805 -246 121867
rect 246 121805 280 121867
rect -100 121729 -84 121763
rect 84 121729 100 121763
rect -146 121679 -112 121695
rect -146 120687 -112 120703
rect 112 121679 146 121695
rect 112 120687 146 120703
rect -100 120619 -84 120653
rect 84 120619 100 120653
rect -100 120511 -84 120545
rect 84 120511 100 120545
rect -146 120461 -112 120477
rect -146 119469 -112 119485
rect 112 120461 146 120477
rect 112 119469 146 119485
rect -100 119401 -84 119435
rect 84 119401 100 119435
rect -100 119293 -84 119327
rect 84 119293 100 119327
rect -146 119243 -112 119259
rect -146 118251 -112 118267
rect 112 119243 146 119259
rect 112 118251 146 118267
rect -100 118183 -84 118217
rect 84 118183 100 118217
rect -100 118075 -84 118109
rect 84 118075 100 118109
rect -146 118025 -112 118041
rect -146 117033 -112 117049
rect 112 118025 146 118041
rect 112 117033 146 117049
rect -100 116965 -84 116999
rect 84 116965 100 116999
rect -100 116857 -84 116891
rect 84 116857 100 116891
rect -146 116807 -112 116823
rect -146 115815 -112 115831
rect 112 116807 146 116823
rect 112 115815 146 115831
rect -100 115747 -84 115781
rect 84 115747 100 115781
rect -100 115639 -84 115673
rect 84 115639 100 115673
rect -146 115589 -112 115605
rect -146 114597 -112 114613
rect 112 115589 146 115605
rect 112 114597 146 114613
rect -100 114529 -84 114563
rect 84 114529 100 114563
rect -100 114421 -84 114455
rect 84 114421 100 114455
rect -146 114371 -112 114387
rect -146 113379 -112 113395
rect 112 114371 146 114387
rect 112 113379 146 113395
rect -100 113311 -84 113345
rect 84 113311 100 113345
rect -100 113203 -84 113237
rect 84 113203 100 113237
rect -146 113153 -112 113169
rect -146 112161 -112 112177
rect 112 113153 146 113169
rect 112 112161 146 112177
rect -100 112093 -84 112127
rect 84 112093 100 112127
rect -100 111985 -84 112019
rect 84 111985 100 112019
rect -146 111935 -112 111951
rect -146 110943 -112 110959
rect 112 111935 146 111951
rect 112 110943 146 110959
rect -100 110875 -84 110909
rect 84 110875 100 110909
rect -100 110767 -84 110801
rect 84 110767 100 110801
rect -146 110717 -112 110733
rect -146 109725 -112 109741
rect 112 110717 146 110733
rect 112 109725 146 109741
rect -100 109657 -84 109691
rect 84 109657 100 109691
rect -100 109549 -84 109583
rect 84 109549 100 109583
rect -146 109499 -112 109515
rect -146 108507 -112 108523
rect 112 109499 146 109515
rect 112 108507 146 108523
rect -100 108439 -84 108473
rect 84 108439 100 108473
rect -100 108331 -84 108365
rect 84 108331 100 108365
rect -146 108281 -112 108297
rect -146 107289 -112 107305
rect 112 108281 146 108297
rect 112 107289 146 107305
rect -100 107221 -84 107255
rect 84 107221 100 107255
rect -100 107113 -84 107147
rect 84 107113 100 107147
rect -146 107063 -112 107079
rect -146 106071 -112 106087
rect 112 107063 146 107079
rect 112 106071 146 106087
rect -100 106003 -84 106037
rect 84 106003 100 106037
rect -100 105895 -84 105929
rect 84 105895 100 105929
rect -146 105845 -112 105861
rect -146 104853 -112 104869
rect 112 105845 146 105861
rect 112 104853 146 104869
rect -100 104785 -84 104819
rect 84 104785 100 104819
rect -100 104677 -84 104711
rect 84 104677 100 104711
rect -146 104627 -112 104643
rect -146 103635 -112 103651
rect 112 104627 146 104643
rect 112 103635 146 103651
rect -100 103567 -84 103601
rect 84 103567 100 103601
rect -100 103459 -84 103493
rect 84 103459 100 103493
rect -146 103409 -112 103425
rect -146 102417 -112 102433
rect 112 103409 146 103425
rect 112 102417 146 102433
rect -100 102349 -84 102383
rect 84 102349 100 102383
rect -100 102241 -84 102275
rect 84 102241 100 102275
rect -146 102191 -112 102207
rect -146 101199 -112 101215
rect 112 102191 146 102207
rect 112 101199 146 101215
rect -100 101131 -84 101165
rect 84 101131 100 101165
rect -100 101023 -84 101057
rect 84 101023 100 101057
rect -146 100973 -112 100989
rect -146 99981 -112 99997
rect 112 100973 146 100989
rect 112 99981 146 99997
rect -100 99913 -84 99947
rect 84 99913 100 99947
rect -100 99805 -84 99839
rect 84 99805 100 99839
rect -146 99755 -112 99771
rect -146 98763 -112 98779
rect 112 99755 146 99771
rect 112 98763 146 98779
rect -100 98695 -84 98729
rect 84 98695 100 98729
rect -100 98587 -84 98621
rect 84 98587 100 98621
rect -146 98537 -112 98553
rect -146 97545 -112 97561
rect 112 98537 146 98553
rect 112 97545 146 97561
rect -100 97477 -84 97511
rect 84 97477 100 97511
rect -100 97369 -84 97403
rect 84 97369 100 97403
rect -146 97319 -112 97335
rect -146 96327 -112 96343
rect 112 97319 146 97335
rect 112 96327 146 96343
rect -100 96259 -84 96293
rect 84 96259 100 96293
rect -100 96151 -84 96185
rect 84 96151 100 96185
rect -146 96101 -112 96117
rect -146 95109 -112 95125
rect 112 96101 146 96117
rect 112 95109 146 95125
rect -100 95041 -84 95075
rect 84 95041 100 95075
rect -100 94933 -84 94967
rect 84 94933 100 94967
rect -146 94883 -112 94899
rect -146 93891 -112 93907
rect 112 94883 146 94899
rect 112 93891 146 93907
rect -100 93823 -84 93857
rect 84 93823 100 93857
rect -100 93715 -84 93749
rect 84 93715 100 93749
rect -146 93665 -112 93681
rect -146 92673 -112 92689
rect 112 93665 146 93681
rect 112 92673 146 92689
rect -100 92605 -84 92639
rect 84 92605 100 92639
rect -100 92497 -84 92531
rect 84 92497 100 92531
rect -146 92447 -112 92463
rect -146 91455 -112 91471
rect 112 92447 146 92463
rect 112 91455 146 91471
rect -100 91387 -84 91421
rect 84 91387 100 91421
rect -100 91279 -84 91313
rect 84 91279 100 91313
rect -146 91229 -112 91245
rect -146 90237 -112 90253
rect 112 91229 146 91245
rect 112 90237 146 90253
rect -100 90169 -84 90203
rect 84 90169 100 90203
rect -100 90061 -84 90095
rect 84 90061 100 90095
rect -146 90011 -112 90027
rect -146 89019 -112 89035
rect 112 90011 146 90027
rect 112 89019 146 89035
rect -100 88951 -84 88985
rect 84 88951 100 88985
rect -100 88843 -84 88877
rect 84 88843 100 88877
rect -146 88793 -112 88809
rect -146 87801 -112 87817
rect 112 88793 146 88809
rect 112 87801 146 87817
rect -100 87733 -84 87767
rect 84 87733 100 87767
rect -100 87625 -84 87659
rect 84 87625 100 87659
rect -146 87575 -112 87591
rect -146 86583 -112 86599
rect 112 87575 146 87591
rect 112 86583 146 86599
rect -100 86515 -84 86549
rect 84 86515 100 86549
rect -100 86407 -84 86441
rect 84 86407 100 86441
rect -146 86357 -112 86373
rect -146 85365 -112 85381
rect 112 86357 146 86373
rect 112 85365 146 85381
rect -100 85297 -84 85331
rect 84 85297 100 85331
rect -100 85189 -84 85223
rect 84 85189 100 85223
rect -146 85139 -112 85155
rect -146 84147 -112 84163
rect 112 85139 146 85155
rect 112 84147 146 84163
rect -100 84079 -84 84113
rect 84 84079 100 84113
rect -100 83971 -84 84005
rect 84 83971 100 84005
rect -146 83921 -112 83937
rect -146 82929 -112 82945
rect 112 83921 146 83937
rect 112 82929 146 82945
rect -100 82861 -84 82895
rect 84 82861 100 82895
rect -100 82753 -84 82787
rect 84 82753 100 82787
rect -146 82703 -112 82719
rect -146 81711 -112 81727
rect 112 82703 146 82719
rect 112 81711 146 81727
rect -100 81643 -84 81677
rect 84 81643 100 81677
rect -100 81535 -84 81569
rect 84 81535 100 81569
rect -146 81485 -112 81501
rect -146 80493 -112 80509
rect 112 81485 146 81501
rect 112 80493 146 80509
rect -100 80425 -84 80459
rect 84 80425 100 80459
rect -100 80317 -84 80351
rect 84 80317 100 80351
rect -146 80267 -112 80283
rect -146 79275 -112 79291
rect 112 80267 146 80283
rect 112 79275 146 79291
rect -100 79207 -84 79241
rect 84 79207 100 79241
rect -100 79099 -84 79133
rect 84 79099 100 79133
rect -146 79049 -112 79065
rect -146 78057 -112 78073
rect 112 79049 146 79065
rect 112 78057 146 78073
rect -100 77989 -84 78023
rect 84 77989 100 78023
rect -100 77881 -84 77915
rect 84 77881 100 77915
rect -146 77831 -112 77847
rect -146 76839 -112 76855
rect 112 77831 146 77847
rect 112 76839 146 76855
rect -100 76771 -84 76805
rect 84 76771 100 76805
rect -100 76663 -84 76697
rect 84 76663 100 76697
rect -146 76613 -112 76629
rect -146 75621 -112 75637
rect 112 76613 146 76629
rect 112 75621 146 75637
rect -100 75553 -84 75587
rect 84 75553 100 75587
rect -100 75445 -84 75479
rect 84 75445 100 75479
rect -146 75395 -112 75411
rect -146 74403 -112 74419
rect 112 75395 146 75411
rect 112 74403 146 74419
rect -100 74335 -84 74369
rect 84 74335 100 74369
rect -100 74227 -84 74261
rect 84 74227 100 74261
rect -146 74177 -112 74193
rect -146 73185 -112 73201
rect 112 74177 146 74193
rect 112 73185 146 73201
rect -100 73117 -84 73151
rect 84 73117 100 73151
rect -100 73009 -84 73043
rect 84 73009 100 73043
rect -146 72959 -112 72975
rect -146 71967 -112 71983
rect 112 72959 146 72975
rect 112 71967 146 71983
rect -100 71899 -84 71933
rect 84 71899 100 71933
rect -100 71791 -84 71825
rect 84 71791 100 71825
rect -146 71741 -112 71757
rect -146 70749 -112 70765
rect 112 71741 146 71757
rect 112 70749 146 70765
rect -100 70681 -84 70715
rect 84 70681 100 70715
rect -100 70573 -84 70607
rect 84 70573 100 70607
rect -146 70523 -112 70539
rect -146 69531 -112 69547
rect 112 70523 146 70539
rect 112 69531 146 69547
rect -100 69463 -84 69497
rect 84 69463 100 69497
rect -100 69355 -84 69389
rect 84 69355 100 69389
rect -146 69305 -112 69321
rect -146 68313 -112 68329
rect 112 69305 146 69321
rect 112 68313 146 68329
rect -100 68245 -84 68279
rect 84 68245 100 68279
rect -100 68137 -84 68171
rect 84 68137 100 68171
rect -146 68087 -112 68103
rect -146 67095 -112 67111
rect 112 68087 146 68103
rect 112 67095 146 67111
rect -100 67027 -84 67061
rect 84 67027 100 67061
rect -100 66919 -84 66953
rect 84 66919 100 66953
rect -146 66869 -112 66885
rect -146 65877 -112 65893
rect 112 66869 146 66885
rect 112 65877 146 65893
rect -100 65809 -84 65843
rect 84 65809 100 65843
rect -100 65701 -84 65735
rect 84 65701 100 65735
rect -146 65651 -112 65667
rect -146 64659 -112 64675
rect 112 65651 146 65667
rect 112 64659 146 64675
rect -100 64591 -84 64625
rect 84 64591 100 64625
rect -100 64483 -84 64517
rect 84 64483 100 64517
rect -146 64433 -112 64449
rect -146 63441 -112 63457
rect 112 64433 146 64449
rect 112 63441 146 63457
rect -100 63373 -84 63407
rect 84 63373 100 63407
rect -100 63265 -84 63299
rect 84 63265 100 63299
rect -146 63215 -112 63231
rect -146 62223 -112 62239
rect 112 63215 146 63231
rect 112 62223 146 62239
rect -100 62155 -84 62189
rect 84 62155 100 62189
rect -100 62047 -84 62081
rect 84 62047 100 62081
rect -146 61997 -112 62013
rect -146 61005 -112 61021
rect 112 61997 146 62013
rect 112 61005 146 61021
rect -100 60937 -84 60971
rect 84 60937 100 60971
rect -100 60829 -84 60863
rect 84 60829 100 60863
rect -146 60779 -112 60795
rect -146 59787 -112 59803
rect 112 60779 146 60795
rect 112 59787 146 59803
rect -100 59719 -84 59753
rect 84 59719 100 59753
rect -100 59611 -84 59645
rect 84 59611 100 59645
rect -146 59561 -112 59577
rect -146 58569 -112 58585
rect 112 59561 146 59577
rect 112 58569 146 58585
rect -100 58501 -84 58535
rect 84 58501 100 58535
rect -100 58393 -84 58427
rect 84 58393 100 58427
rect -146 58343 -112 58359
rect -146 57351 -112 57367
rect 112 58343 146 58359
rect 112 57351 146 57367
rect -100 57283 -84 57317
rect 84 57283 100 57317
rect -100 57175 -84 57209
rect 84 57175 100 57209
rect -146 57125 -112 57141
rect -146 56133 -112 56149
rect 112 57125 146 57141
rect 112 56133 146 56149
rect -100 56065 -84 56099
rect 84 56065 100 56099
rect -100 55957 -84 55991
rect 84 55957 100 55991
rect -146 55907 -112 55923
rect -146 54915 -112 54931
rect 112 55907 146 55923
rect 112 54915 146 54931
rect -100 54847 -84 54881
rect 84 54847 100 54881
rect -100 54739 -84 54773
rect 84 54739 100 54773
rect -146 54689 -112 54705
rect -146 53697 -112 53713
rect 112 54689 146 54705
rect 112 53697 146 53713
rect -100 53629 -84 53663
rect 84 53629 100 53663
rect -100 53521 -84 53555
rect 84 53521 100 53555
rect -146 53471 -112 53487
rect -146 52479 -112 52495
rect 112 53471 146 53487
rect 112 52479 146 52495
rect -100 52411 -84 52445
rect 84 52411 100 52445
rect -100 52303 -84 52337
rect 84 52303 100 52337
rect -146 52253 -112 52269
rect -146 51261 -112 51277
rect 112 52253 146 52269
rect 112 51261 146 51277
rect -100 51193 -84 51227
rect 84 51193 100 51227
rect -100 51085 -84 51119
rect 84 51085 100 51119
rect -146 51035 -112 51051
rect -146 50043 -112 50059
rect 112 51035 146 51051
rect 112 50043 146 50059
rect -100 49975 -84 50009
rect 84 49975 100 50009
rect -100 49867 -84 49901
rect 84 49867 100 49901
rect -146 49817 -112 49833
rect -146 48825 -112 48841
rect 112 49817 146 49833
rect 112 48825 146 48841
rect -100 48757 -84 48791
rect 84 48757 100 48791
rect -100 48649 -84 48683
rect 84 48649 100 48683
rect -146 48599 -112 48615
rect -146 47607 -112 47623
rect 112 48599 146 48615
rect 112 47607 146 47623
rect -100 47539 -84 47573
rect 84 47539 100 47573
rect -100 47431 -84 47465
rect 84 47431 100 47465
rect -146 47381 -112 47397
rect -146 46389 -112 46405
rect 112 47381 146 47397
rect 112 46389 146 46405
rect -100 46321 -84 46355
rect 84 46321 100 46355
rect -100 46213 -84 46247
rect 84 46213 100 46247
rect -146 46163 -112 46179
rect -146 45171 -112 45187
rect 112 46163 146 46179
rect 112 45171 146 45187
rect -100 45103 -84 45137
rect 84 45103 100 45137
rect -100 44995 -84 45029
rect 84 44995 100 45029
rect -146 44945 -112 44961
rect -146 43953 -112 43969
rect 112 44945 146 44961
rect 112 43953 146 43969
rect -100 43885 -84 43919
rect 84 43885 100 43919
rect -100 43777 -84 43811
rect 84 43777 100 43811
rect -146 43727 -112 43743
rect -146 42735 -112 42751
rect 112 43727 146 43743
rect 112 42735 146 42751
rect -100 42667 -84 42701
rect 84 42667 100 42701
rect -100 42559 -84 42593
rect 84 42559 100 42593
rect -146 42509 -112 42525
rect -146 41517 -112 41533
rect 112 42509 146 42525
rect 112 41517 146 41533
rect -100 41449 -84 41483
rect 84 41449 100 41483
rect -100 41341 -84 41375
rect 84 41341 100 41375
rect -146 41291 -112 41307
rect -146 40299 -112 40315
rect 112 41291 146 41307
rect 112 40299 146 40315
rect -100 40231 -84 40265
rect 84 40231 100 40265
rect -100 40123 -84 40157
rect 84 40123 100 40157
rect -146 40073 -112 40089
rect -146 39081 -112 39097
rect 112 40073 146 40089
rect 112 39081 146 39097
rect -100 39013 -84 39047
rect 84 39013 100 39047
rect -100 38905 -84 38939
rect 84 38905 100 38939
rect -146 38855 -112 38871
rect -146 37863 -112 37879
rect 112 38855 146 38871
rect 112 37863 146 37879
rect -100 37795 -84 37829
rect 84 37795 100 37829
rect -100 37687 -84 37721
rect 84 37687 100 37721
rect -146 37637 -112 37653
rect -146 36645 -112 36661
rect 112 37637 146 37653
rect 112 36645 146 36661
rect -100 36577 -84 36611
rect 84 36577 100 36611
rect -100 36469 -84 36503
rect 84 36469 100 36503
rect -146 36419 -112 36435
rect -146 35427 -112 35443
rect 112 36419 146 36435
rect 112 35427 146 35443
rect -100 35359 -84 35393
rect 84 35359 100 35393
rect -100 35251 -84 35285
rect 84 35251 100 35285
rect -146 35201 -112 35217
rect -146 34209 -112 34225
rect 112 35201 146 35217
rect 112 34209 146 34225
rect -100 34141 -84 34175
rect 84 34141 100 34175
rect -100 34033 -84 34067
rect 84 34033 100 34067
rect -146 33983 -112 33999
rect -146 32991 -112 33007
rect 112 33983 146 33999
rect 112 32991 146 33007
rect -100 32923 -84 32957
rect 84 32923 100 32957
rect -100 32815 -84 32849
rect 84 32815 100 32849
rect -146 32765 -112 32781
rect -146 31773 -112 31789
rect 112 32765 146 32781
rect 112 31773 146 31789
rect -100 31705 -84 31739
rect 84 31705 100 31739
rect -100 31597 -84 31631
rect 84 31597 100 31631
rect -146 31547 -112 31563
rect -146 30555 -112 30571
rect 112 31547 146 31563
rect 112 30555 146 30571
rect -100 30487 -84 30521
rect 84 30487 100 30521
rect -100 30379 -84 30413
rect 84 30379 100 30413
rect -146 30329 -112 30345
rect -146 29337 -112 29353
rect 112 30329 146 30345
rect 112 29337 146 29353
rect -100 29269 -84 29303
rect 84 29269 100 29303
rect -100 29161 -84 29195
rect 84 29161 100 29195
rect -146 29111 -112 29127
rect -146 28119 -112 28135
rect 112 29111 146 29127
rect 112 28119 146 28135
rect -100 28051 -84 28085
rect 84 28051 100 28085
rect -100 27943 -84 27977
rect 84 27943 100 27977
rect -146 27893 -112 27909
rect -146 26901 -112 26917
rect 112 27893 146 27909
rect 112 26901 146 26917
rect -100 26833 -84 26867
rect 84 26833 100 26867
rect -100 26725 -84 26759
rect 84 26725 100 26759
rect -146 26675 -112 26691
rect -146 25683 -112 25699
rect 112 26675 146 26691
rect 112 25683 146 25699
rect -100 25615 -84 25649
rect 84 25615 100 25649
rect -100 25507 -84 25541
rect 84 25507 100 25541
rect -146 25457 -112 25473
rect -146 24465 -112 24481
rect 112 25457 146 25473
rect 112 24465 146 24481
rect -100 24397 -84 24431
rect 84 24397 100 24431
rect -100 24289 -84 24323
rect 84 24289 100 24323
rect -146 24239 -112 24255
rect -146 23247 -112 23263
rect 112 24239 146 24255
rect 112 23247 146 23263
rect -100 23179 -84 23213
rect 84 23179 100 23213
rect -100 23071 -84 23105
rect 84 23071 100 23105
rect -146 23021 -112 23037
rect -146 22029 -112 22045
rect 112 23021 146 23037
rect 112 22029 146 22045
rect -100 21961 -84 21995
rect 84 21961 100 21995
rect -100 21853 -84 21887
rect 84 21853 100 21887
rect -146 21803 -112 21819
rect -146 20811 -112 20827
rect 112 21803 146 21819
rect 112 20811 146 20827
rect -100 20743 -84 20777
rect 84 20743 100 20777
rect -100 20635 -84 20669
rect 84 20635 100 20669
rect -146 20585 -112 20601
rect -146 19593 -112 19609
rect 112 20585 146 20601
rect 112 19593 146 19609
rect -100 19525 -84 19559
rect 84 19525 100 19559
rect -100 19417 -84 19451
rect 84 19417 100 19451
rect -146 19367 -112 19383
rect -146 18375 -112 18391
rect 112 19367 146 19383
rect 112 18375 146 18391
rect -100 18307 -84 18341
rect 84 18307 100 18341
rect -100 18199 -84 18233
rect 84 18199 100 18233
rect -146 18149 -112 18165
rect -146 17157 -112 17173
rect 112 18149 146 18165
rect 112 17157 146 17173
rect -100 17089 -84 17123
rect 84 17089 100 17123
rect -100 16981 -84 17015
rect 84 16981 100 17015
rect -146 16931 -112 16947
rect -146 15939 -112 15955
rect 112 16931 146 16947
rect 112 15939 146 15955
rect -100 15871 -84 15905
rect 84 15871 100 15905
rect -100 15763 -84 15797
rect 84 15763 100 15797
rect -146 15713 -112 15729
rect -146 14721 -112 14737
rect 112 15713 146 15729
rect 112 14721 146 14737
rect -100 14653 -84 14687
rect 84 14653 100 14687
rect -100 14545 -84 14579
rect 84 14545 100 14579
rect -146 14495 -112 14511
rect -146 13503 -112 13519
rect 112 14495 146 14511
rect 112 13503 146 13519
rect -100 13435 -84 13469
rect 84 13435 100 13469
rect -100 13327 -84 13361
rect 84 13327 100 13361
rect -146 13277 -112 13293
rect -146 12285 -112 12301
rect 112 13277 146 13293
rect 112 12285 146 12301
rect -100 12217 -84 12251
rect 84 12217 100 12251
rect -100 12109 -84 12143
rect 84 12109 100 12143
rect -146 12059 -112 12075
rect -146 11067 -112 11083
rect 112 12059 146 12075
rect 112 11067 146 11083
rect -100 10999 -84 11033
rect 84 10999 100 11033
rect -100 10891 -84 10925
rect 84 10891 100 10925
rect -146 10841 -112 10857
rect -146 9849 -112 9865
rect 112 10841 146 10857
rect 112 9849 146 9865
rect -100 9781 -84 9815
rect 84 9781 100 9815
rect -100 9673 -84 9707
rect 84 9673 100 9707
rect -146 9623 -112 9639
rect -146 8631 -112 8647
rect 112 9623 146 9639
rect 112 8631 146 8647
rect -100 8563 -84 8597
rect 84 8563 100 8597
rect -100 8455 -84 8489
rect 84 8455 100 8489
rect -146 8405 -112 8421
rect -146 7413 -112 7429
rect 112 8405 146 8421
rect 112 7413 146 7429
rect -100 7345 -84 7379
rect 84 7345 100 7379
rect -100 7237 -84 7271
rect 84 7237 100 7271
rect -146 7187 -112 7203
rect -146 6195 -112 6211
rect 112 7187 146 7203
rect 112 6195 146 6211
rect -100 6127 -84 6161
rect 84 6127 100 6161
rect -100 6019 -84 6053
rect 84 6019 100 6053
rect -146 5969 -112 5985
rect -146 4977 -112 4993
rect 112 5969 146 5985
rect 112 4977 146 4993
rect -100 4909 -84 4943
rect 84 4909 100 4943
rect -100 4801 -84 4835
rect 84 4801 100 4835
rect -146 4751 -112 4767
rect -146 3759 -112 3775
rect 112 4751 146 4767
rect 112 3759 146 3775
rect -100 3691 -84 3725
rect 84 3691 100 3725
rect -100 3583 -84 3617
rect 84 3583 100 3617
rect -146 3533 -112 3549
rect -146 2541 -112 2557
rect 112 3533 146 3549
rect 112 2541 146 2557
rect -100 2473 -84 2507
rect 84 2473 100 2507
rect -100 2365 -84 2399
rect 84 2365 100 2399
rect -146 2315 -112 2331
rect -146 1323 -112 1339
rect 112 2315 146 2331
rect 112 1323 146 1339
rect -100 1255 -84 1289
rect 84 1255 100 1289
rect -100 1147 -84 1181
rect 84 1147 100 1181
rect -146 1097 -112 1113
rect -146 105 -112 121
rect 112 1097 146 1113
rect 112 105 146 121
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -121 -112 -105
rect -146 -1113 -112 -1097
rect 112 -121 146 -105
rect 112 -1113 146 -1097
rect -100 -1181 -84 -1147
rect 84 -1181 100 -1147
rect -100 -1289 -84 -1255
rect 84 -1289 100 -1255
rect -146 -1339 -112 -1323
rect -146 -2331 -112 -2315
rect 112 -1339 146 -1323
rect 112 -2331 146 -2315
rect -100 -2399 -84 -2365
rect 84 -2399 100 -2365
rect -100 -2507 -84 -2473
rect 84 -2507 100 -2473
rect -146 -2557 -112 -2541
rect -146 -3549 -112 -3533
rect 112 -2557 146 -2541
rect 112 -3549 146 -3533
rect -100 -3617 -84 -3583
rect 84 -3617 100 -3583
rect -100 -3725 -84 -3691
rect 84 -3725 100 -3691
rect -146 -3775 -112 -3759
rect -146 -4767 -112 -4751
rect 112 -3775 146 -3759
rect 112 -4767 146 -4751
rect -100 -4835 -84 -4801
rect 84 -4835 100 -4801
rect -100 -4943 -84 -4909
rect 84 -4943 100 -4909
rect -146 -4993 -112 -4977
rect -146 -5985 -112 -5969
rect 112 -4993 146 -4977
rect 112 -5985 146 -5969
rect -100 -6053 -84 -6019
rect 84 -6053 100 -6019
rect -100 -6161 -84 -6127
rect 84 -6161 100 -6127
rect -146 -6211 -112 -6195
rect -146 -7203 -112 -7187
rect 112 -6211 146 -6195
rect 112 -7203 146 -7187
rect -100 -7271 -84 -7237
rect 84 -7271 100 -7237
rect -100 -7379 -84 -7345
rect 84 -7379 100 -7345
rect -146 -7429 -112 -7413
rect -146 -8421 -112 -8405
rect 112 -7429 146 -7413
rect 112 -8421 146 -8405
rect -100 -8489 -84 -8455
rect 84 -8489 100 -8455
rect -100 -8597 -84 -8563
rect 84 -8597 100 -8563
rect -146 -8647 -112 -8631
rect -146 -9639 -112 -9623
rect 112 -8647 146 -8631
rect 112 -9639 146 -9623
rect -100 -9707 -84 -9673
rect 84 -9707 100 -9673
rect -100 -9815 -84 -9781
rect 84 -9815 100 -9781
rect -146 -9865 -112 -9849
rect -146 -10857 -112 -10841
rect 112 -9865 146 -9849
rect 112 -10857 146 -10841
rect -100 -10925 -84 -10891
rect 84 -10925 100 -10891
rect -100 -11033 -84 -10999
rect 84 -11033 100 -10999
rect -146 -11083 -112 -11067
rect -146 -12075 -112 -12059
rect 112 -11083 146 -11067
rect 112 -12075 146 -12059
rect -100 -12143 -84 -12109
rect 84 -12143 100 -12109
rect -100 -12251 -84 -12217
rect 84 -12251 100 -12217
rect -146 -12301 -112 -12285
rect -146 -13293 -112 -13277
rect 112 -12301 146 -12285
rect 112 -13293 146 -13277
rect -100 -13361 -84 -13327
rect 84 -13361 100 -13327
rect -100 -13469 -84 -13435
rect 84 -13469 100 -13435
rect -146 -13519 -112 -13503
rect -146 -14511 -112 -14495
rect 112 -13519 146 -13503
rect 112 -14511 146 -14495
rect -100 -14579 -84 -14545
rect 84 -14579 100 -14545
rect -100 -14687 -84 -14653
rect 84 -14687 100 -14653
rect -146 -14737 -112 -14721
rect -146 -15729 -112 -15713
rect 112 -14737 146 -14721
rect 112 -15729 146 -15713
rect -100 -15797 -84 -15763
rect 84 -15797 100 -15763
rect -100 -15905 -84 -15871
rect 84 -15905 100 -15871
rect -146 -15955 -112 -15939
rect -146 -16947 -112 -16931
rect 112 -15955 146 -15939
rect 112 -16947 146 -16931
rect -100 -17015 -84 -16981
rect 84 -17015 100 -16981
rect -100 -17123 -84 -17089
rect 84 -17123 100 -17089
rect -146 -17173 -112 -17157
rect -146 -18165 -112 -18149
rect 112 -17173 146 -17157
rect 112 -18165 146 -18149
rect -100 -18233 -84 -18199
rect 84 -18233 100 -18199
rect -100 -18341 -84 -18307
rect 84 -18341 100 -18307
rect -146 -18391 -112 -18375
rect -146 -19383 -112 -19367
rect 112 -18391 146 -18375
rect 112 -19383 146 -19367
rect -100 -19451 -84 -19417
rect 84 -19451 100 -19417
rect -100 -19559 -84 -19525
rect 84 -19559 100 -19525
rect -146 -19609 -112 -19593
rect -146 -20601 -112 -20585
rect 112 -19609 146 -19593
rect 112 -20601 146 -20585
rect -100 -20669 -84 -20635
rect 84 -20669 100 -20635
rect -100 -20777 -84 -20743
rect 84 -20777 100 -20743
rect -146 -20827 -112 -20811
rect -146 -21819 -112 -21803
rect 112 -20827 146 -20811
rect 112 -21819 146 -21803
rect -100 -21887 -84 -21853
rect 84 -21887 100 -21853
rect -100 -21995 -84 -21961
rect 84 -21995 100 -21961
rect -146 -22045 -112 -22029
rect -146 -23037 -112 -23021
rect 112 -22045 146 -22029
rect 112 -23037 146 -23021
rect -100 -23105 -84 -23071
rect 84 -23105 100 -23071
rect -100 -23213 -84 -23179
rect 84 -23213 100 -23179
rect -146 -23263 -112 -23247
rect -146 -24255 -112 -24239
rect 112 -23263 146 -23247
rect 112 -24255 146 -24239
rect -100 -24323 -84 -24289
rect 84 -24323 100 -24289
rect -100 -24431 -84 -24397
rect 84 -24431 100 -24397
rect -146 -24481 -112 -24465
rect -146 -25473 -112 -25457
rect 112 -24481 146 -24465
rect 112 -25473 146 -25457
rect -100 -25541 -84 -25507
rect 84 -25541 100 -25507
rect -100 -25649 -84 -25615
rect 84 -25649 100 -25615
rect -146 -25699 -112 -25683
rect -146 -26691 -112 -26675
rect 112 -25699 146 -25683
rect 112 -26691 146 -26675
rect -100 -26759 -84 -26725
rect 84 -26759 100 -26725
rect -100 -26867 -84 -26833
rect 84 -26867 100 -26833
rect -146 -26917 -112 -26901
rect -146 -27909 -112 -27893
rect 112 -26917 146 -26901
rect 112 -27909 146 -27893
rect -100 -27977 -84 -27943
rect 84 -27977 100 -27943
rect -100 -28085 -84 -28051
rect 84 -28085 100 -28051
rect -146 -28135 -112 -28119
rect -146 -29127 -112 -29111
rect 112 -28135 146 -28119
rect 112 -29127 146 -29111
rect -100 -29195 -84 -29161
rect 84 -29195 100 -29161
rect -100 -29303 -84 -29269
rect 84 -29303 100 -29269
rect -146 -29353 -112 -29337
rect -146 -30345 -112 -30329
rect 112 -29353 146 -29337
rect 112 -30345 146 -30329
rect -100 -30413 -84 -30379
rect 84 -30413 100 -30379
rect -100 -30521 -84 -30487
rect 84 -30521 100 -30487
rect -146 -30571 -112 -30555
rect -146 -31563 -112 -31547
rect 112 -30571 146 -30555
rect 112 -31563 146 -31547
rect -100 -31631 -84 -31597
rect 84 -31631 100 -31597
rect -100 -31739 -84 -31705
rect 84 -31739 100 -31705
rect -146 -31789 -112 -31773
rect -146 -32781 -112 -32765
rect 112 -31789 146 -31773
rect 112 -32781 146 -32765
rect -100 -32849 -84 -32815
rect 84 -32849 100 -32815
rect -100 -32957 -84 -32923
rect 84 -32957 100 -32923
rect -146 -33007 -112 -32991
rect -146 -33999 -112 -33983
rect 112 -33007 146 -32991
rect 112 -33999 146 -33983
rect -100 -34067 -84 -34033
rect 84 -34067 100 -34033
rect -100 -34175 -84 -34141
rect 84 -34175 100 -34141
rect -146 -34225 -112 -34209
rect -146 -35217 -112 -35201
rect 112 -34225 146 -34209
rect 112 -35217 146 -35201
rect -100 -35285 -84 -35251
rect 84 -35285 100 -35251
rect -100 -35393 -84 -35359
rect 84 -35393 100 -35359
rect -146 -35443 -112 -35427
rect -146 -36435 -112 -36419
rect 112 -35443 146 -35427
rect 112 -36435 146 -36419
rect -100 -36503 -84 -36469
rect 84 -36503 100 -36469
rect -100 -36611 -84 -36577
rect 84 -36611 100 -36577
rect -146 -36661 -112 -36645
rect -146 -37653 -112 -37637
rect 112 -36661 146 -36645
rect 112 -37653 146 -37637
rect -100 -37721 -84 -37687
rect 84 -37721 100 -37687
rect -100 -37829 -84 -37795
rect 84 -37829 100 -37795
rect -146 -37879 -112 -37863
rect -146 -38871 -112 -38855
rect 112 -37879 146 -37863
rect 112 -38871 146 -38855
rect -100 -38939 -84 -38905
rect 84 -38939 100 -38905
rect -100 -39047 -84 -39013
rect 84 -39047 100 -39013
rect -146 -39097 -112 -39081
rect -146 -40089 -112 -40073
rect 112 -39097 146 -39081
rect 112 -40089 146 -40073
rect -100 -40157 -84 -40123
rect 84 -40157 100 -40123
rect -100 -40265 -84 -40231
rect 84 -40265 100 -40231
rect -146 -40315 -112 -40299
rect -146 -41307 -112 -41291
rect 112 -40315 146 -40299
rect 112 -41307 146 -41291
rect -100 -41375 -84 -41341
rect 84 -41375 100 -41341
rect -100 -41483 -84 -41449
rect 84 -41483 100 -41449
rect -146 -41533 -112 -41517
rect -146 -42525 -112 -42509
rect 112 -41533 146 -41517
rect 112 -42525 146 -42509
rect -100 -42593 -84 -42559
rect 84 -42593 100 -42559
rect -100 -42701 -84 -42667
rect 84 -42701 100 -42667
rect -146 -42751 -112 -42735
rect -146 -43743 -112 -43727
rect 112 -42751 146 -42735
rect 112 -43743 146 -43727
rect -100 -43811 -84 -43777
rect 84 -43811 100 -43777
rect -100 -43919 -84 -43885
rect 84 -43919 100 -43885
rect -146 -43969 -112 -43953
rect -146 -44961 -112 -44945
rect 112 -43969 146 -43953
rect 112 -44961 146 -44945
rect -100 -45029 -84 -44995
rect 84 -45029 100 -44995
rect -100 -45137 -84 -45103
rect 84 -45137 100 -45103
rect -146 -45187 -112 -45171
rect -146 -46179 -112 -46163
rect 112 -45187 146 -45171
rect 112 -46179 146 -46163
rect -100 -46247 -84 -46213
rect 84 -46247 100 -46213
rect -100 -46355 -84 -46321
rect 84 -46355 100 -46321
rect -146 -46405 -112 -46389
rect -146 -47397 -112 -47381
rect 112 -46405 146 -46389
rect 112 -47397 146 -47381
rect -100 -47465 -84 -47431
rect 84 -47465 100 -47431
rect -100 -47573 -84 -47539
rect 84 -47573 100 -47539
rect -146 -47623 -112 -47607
rect -146 -48615 -112 -48599
rect 112 -47623 146 -47607
rect 112 -48615 146 -48599
rect -100 -48683 -84 -48649
rect 84 -48683 100 -48649
rect -100 -48791 -84 -48757
rect 84 -48791 100 -48757
rect -146 -48841 -112 -48825
rect -146 -49833 -112 -49817
rect 112 -48841 146 -48825
rect 112 -49833 146 -49817
rect -100 -49901 -84 -49867
rect 84 -49901 100 -49867
rect -100 -50009 -84 -49975
rect 84 -50009 100 -49975
rect -146 -50059 -112 -50043
rect -146 -51051 -112 -51035
rect 112 -50059 146 -50043
rect 112 -51051 146 -51035
rect -100 -51119 -84 -51085
rect 84 -51119 100 -51085
rect -100 -51227 -84 -51193
rect 84 -51227 100 -51193
rect -146 -51277 -112 -51261
rect -146 -52269 -112 -52253
rect 112 -51277 146 -51261
rect 112 -52269 146 -52253
rect -100 -52337 -84 -52303
rect 84 -52337 100 -52303
rect -100 -52445 -84 -52411
rect 84 -52445 100 -52411
rect -146 -52495 -112 -52479
rect -146 -53487 -112 -53471
rect 112 -52495 146 -52479
rect 112 -53487 146 -53471
rect -100 -53555 -84 -53521
rect 84 -53555 100 -53521
rect -100 -53663 -84 -53629
rect 84 -53663 100 -53629
rect -146 -53713 -112 -53697
rect -146 -54705 -112 -54689
rect 112 -53713 146 -53697
rect 112 -54705 146 -54689
rect -100 -54773 -84 -54739
rect 84 -54773 100 -54739
rect -100 -54881 -84 -54847
rect 84 -54881 100 -54847
rect -146 -54931 -112 -54915
rect -146 -55923 -112 -55907
rect 112 -54931 146 -54915
rect 112 -55923 146 -55907
rect -100 -55991 -84 -55957
rect 84 -55991 100 -55957
rect -100 -56099 -84 -56065
rect 84 -56099 100 -56065
rect -146 -56149 -112 -56133
rect -146 -57141 -112 -57125
rect 112 -56149 146 -56133
rect 112 -57141 146 -57125
rect -100 -57209 -84 -57175
rect 84 -57209 100 -57175
rect -100 -57317 -84 -57283
rect 84 -57317 100 -57283
rect -146 -57367 -112 -57351
rect -146 -58359 -112 -58343
rect 112 -57367 146 -57351
rect 112 -58359 146 -58343
rect -100 -58427 -84 -58393
rect 84 -58427 100 -58393
rect -100 -58535 -84 -58501
rect 84 -58535 100 -58501
rect -146 -58585 -112 -58569
rect -146 -59577 -112 -59561
rect 112 -58585 146 -58569
rect 112 -59577 146 -59561
rect -100 -59645 -84 -59611
rect 84 -59645 100 -59611
rect -100 -59753 -84 -59719
rect 84 -59753 100 -59719
rect -146 -59803 -112 -59787
rect -146 -60795 -112 -60779
rect 112 -59803 146 -59787
rect 112 -60795 146 -60779
rect -100 -60863 -84 -60829
rect 84 -60863 100 -60829
rect -100 -60971 -84 -60937
rect 84 -60971 100 -60937
rect -146 -61021 -112 -61005
rect -146 -62013 -112 -61997
rect 112 -61021 146 -61005
rect 112 -62013 146 -61997
rect -100 -62081 -84 -62047
rect 84 -62081 100 -62047
rect -100 -62189 -84 -62155
rect 84 -62189 100 -62155
rect -146 -62239 -112 -62223
rect -146 -63231 -112 -63215
rect 112 -62239 146 -62223
rect 112 -63231 146 -63215
rect -100 -63299 -84 -63265
rect 84 -63299 100 -63265
rect -100 -63407 -84 -63373
rect 84 -63407 100 -63373
rect -146 -63457 -112 -63441
rect -146 -64449 -112 -64433
rect 112 -63457 146 -63441
rect 112 -64449 146 -64433
rect -100 -64517 -84 -64483
rect 84 -64517 100 -64483
rect -100 -64625 -84 -64591
rect 84 -64625 100 -64591
rect -146 -64675 -112 -64659
rect -146 -65667 -112 -65651
rect 112 -64675 146 -64659
rect 112 -65667 146 -65651
rect -100 -65735 -84 -65701
rect 84 -65735 100 -65701
rect -100 -65843 -84 -65809
rect 84 -65843 100 -65809
rect -146 -65893 -112 -65877
rect -146 -66885 -112 -66869
rect 112 -65893 146 -65877
rect 112 -66885 146 -66869
rect -100 -66953 -84 -66919
rect 84 -66953 100 -66919
rect -100 -67061 -84 -67027
rect 84 -67061 100 -67027
rect -146 -67111 -112 -67095
rect -146 -68103 -112 -68087
rect 112 -67111 146 -67095
rect 112 -68103 146 -68087
rect -100 -68171 -84 -68137
rect 84 -68171 100 -68137
rect -100 -68279 -84 -68245
rect 84 -68279 100 -68245
rect -146 -68329 -112 -68313
rect -146 -69321 -112 -69305
rect 112 -68329 146 -68313
rect 112 -69321 146 -69305
rect -100 -69389 -84 -69355
rect 84 -69389 100 -69355
rect -100 -69497 -84 -69463
rect 84 -69497 100 -69463
rect -146 -69547 -112 -69531
rect -146 -70539 -112 -70523
rect 112 -69547 146 -69531
rect 112 -70539 146 -70523
rect -100 -70607 -84 -70573
rect 84 -70607 100 -70573
rect -100 -70715 -84 -70681
rect 84 -70715 100 -70681
rect -146 -70765 -112 -70749
rect -146 -71757 -112 -71741
rect 112 -70765 146 -70749
rect 112 -71757 146 -71741
rect -100 -71825 -84 -71791
rect 84 -71825 100 -71791
rect -100 -71933 -84 -71899
rect 84 -71933 100 -71899
rect -146 -71983 -112 -71967
rect -146 -72975 -112 -72959
rect 112 -71983 146 -71967
rect 112 -72975 146 -72959
rect -100 -73043 -84 -73009
rect 84 -73043 100 -73009
rect -100 -73151 -84 -73117
rect 84 -73151 100 -73117
rect -146 -73201 -112 -73185
rect -146 -74193 -112 -74177
rect 112 -73201 146 -73185
rect 112 -74193 146 -74177
rect -100 -74261 -84 -74227
rect 84 -74261 100 -74227
rect -100 -74369 -84 -74335
rect 84 -74369 100 -74335
rect -146 -74419 -112 -74403
rect -146 -75411 -112 -75395
rect 112 -74419 146 -74403
rect 112 -75411 146 -75395
rect -100 -75479 -84 -75445
rect 84 -75479 100 -75445
rect -100 -75587 -84 -75553
rect 84 -75587 100 -75553
rect -146 -75637 -112 -75621
rect -146 -76629 -112 -76613
rect 112 -75637 146 -75621
rect 112 -76629 146 -76613
rect -100 -76697 -84 -76663
rect 84 -76697 100 -76663
rect -100 -76805 -84 -76771
rect 84 -76805 100 -76771
rect -146 -76855 -112 -76839
rect -146 -77847 -112 -77831
rect 112 -76855 146 -76839
rect 112 -77847 146 -77831
rect -100 -77915 -84 -77881
rect 84 -77915 100 -77881
rect -100 -78023 -84 -77989
rect 84 -78023 100 -77989
rect -146 -78073 -112 -78057
rect -146 -79065 -112 -79049
rect 112 -78073 146 -78057
rect 112 -79065 146 -79049
rect -100 -79133 -84 -79099
rect 84 -79133 100 -79099
rect -100 -79241 -84 -79207
rect 84 -79241 100 -79207
rect -146 -79291 -112 -79275
rect -146 -80283 -112 -80267
rect 112 -79291 146 -79275
rect 112 -80283 146 -80267
rect -100 -80351 -84 -80317
rect 84 -80351 100 -80317
rect -100 -80459 -84 -80425
rect 84 -80459 100 -80425
rect -146 -80509 -112 -80493
rect -146 -81501 -112 -81485
rect 112 -80509 146 -80493
rect 112 -81501 146 -81485
rect -100 -81569 -84 -81535
rect 84 -81569 100 -81535
rect -100 -81677 -84 -81643
rect 84 -81677 100 -81643
rect -146 -81727 -112 -81711
rect -146 -82719 -112 -82703
rect 112 -81727 146 -81711
rect 112 -82719 146 -82703
rect -100 -82787 -84 -82753
rect 84 -82787 100 -82753
rect -100 -82895 -84 -82861
rect 84 -82895 100 -82861
rect -146 -82945 -112 -82929
rect -146 -83937 -112 -83921
rect 112 -82945 146 -82929
rect 112 -83937 146 -83921
rect -100 -84005 -84 -83971
rect 84 -84005 100 -83971
rect -100 -84113 -84 -84079
rect 84 -84113 100 -84079
rect -146 -84163 -112 -84147
rect -146 -85155 -112 -85139
rect 112 -84163 146 -84147
rect 112 -85155 146 -85139
rect -100 -85223 -84 -85189
rect 84 -85223 100 -85189
rect -100 -85331 -84 -85297
rect 84 -85331 100 -85297
rect -146 -85381 -112 -85365
rect -146 -86373 -112 -86357
rect 112 -85381 146 -85365
rect 112 -86373 146 -86357
rect -100 -86441 -84 -86407
rect 84 -86441 100 -86407
rect -100 -86549 -84 -86515
rect 84 -86549 100 -86515
rect -146 -86599 -112 -86583
rect -146 -87591 -112 -87575
rect 112 -86599 146 -86583
rect 112 -87591 146 -87575
rect -100 -87659 -84 -87625
rect 84 -87659 100 -87625
rect -100 -87767 -84 -87733
rect 84 -87767 100 -87733
rect -146 -87817 -112 -87801
rect -146 -88809 -112 -88793
rect 112 -87817 146 -87801
rect 112 -88809 146 -88793
rect -100 -88877 -84 -88843
rect 84 -88877 100 -88843
rect -100 -88985 -84 -88951
rect 84 -88985 100 -88951
rect -146 -89035 -112 -89019
rect -146 -90027 -112 -90011
rect 112 -89035 146 -89019
rect 112 -90027 146 -90011
rect -100 -90095 -84 -90061
rect 84 -90095 100 -90061
rect -100 -90203 -84 -90169
rect 84 -90203 100 -90169
rect -146 -90253 -112 -90237
rect -146 -91245 -112 -91229
rect 112 -90253 146 -90237
rect 112 -91245 146 -91229
rect -100 -91313 -84 -91279
rect 84 -91313 100 -91279
rect -100 -91421 -84 -91387
rect 84 -91421 100 -91387
rect -146 -91471 -112 -91455
rect -146 -92463 -112 -92447
rect 112 -91471 146 -91455
rect 112 -92463 146 -92447
rect -100 -92531 -84 -92497
rect 84 -92531 100 -92497
rect -100 -92639 -84 -92605
rect 84 -92639 100 -92605
rect -146 -92689 -112 -92673
rect -146 -93681 -112 -93665
rect 112 -92689 146 -92673
rect 112 -93681 146 -93665
rect -100 -93749 -84 -93715
rect 84 -93749 100 -93715
rect -100 -93857 -84 -93823
rect 84 -93857 100 -93823
rect -146 -93907 -112 -93891
rect -146 -94899 -112 -94883
rect 112 -93907 146 -93891
rect 112 -94899 146 -94883
rect -100 -94967 -84 -94933
rect 84 -94967 100 -94933
rect -100 -95075 -84 -95041
rect 84 -95075 100 -95041
rect -146 -95125 -112 -95109
rect -146 -96117 -112 -96101
rect 112 -95125 146 -95109
rect 112 -96117 146 -96101
rect -100 -96185 -84 -96151
rect 84 -96185 100 -96151
rect -100 -96293 -84 -96259
rect 84 -96293 100 -96259
rect -146 -96343 -112 -96327
rect -146 -97335 -112 -97319
rect 112 -96343 146 -96327
rect 112 -97335 146 -97319
rect -100 -97403 -84 -97369
rect 84 -97403 100 -97369
rect -100 -97511 -84 -97477
rect 84 -97511 100 -97477
rect -146 -97561 -112 -97545
rect -146 -98553 -112 -98537
rect 112 -97561 146 -97545
rect 112 -98553 146 -98537
rect -100 -98621 -84 -98587
rect 84 -98621 100 -98587
rect -100 -98729 -84 -98695
rect 84 -98729 100 -98695
rect -146 -98779 -112 -98763
rect -146 -99771 -112 -99755
rect 112 -98779 146 -98763
rect 112 -99771 146 -99755
rect -100 -99839 -84 -99805
rect 84 -99839 100 -99805
rect -100 -99947 -84 -99913
rect 84 -99947 100 -99913
rect -146 -99997 -112 -99981
rect -146 -100989 -112 -100973
rect 112 -99997 146 -99981
rect 112 -100989 146 -100973
rect -100 -101057 -84 -101023
rect 84 -101057 100 -101023
rect -100 -101165 -84 -101131
rect 84 -101165 100 -101131
rect -146 -101215 -112 -101199
rect -146 -102207 -112 -102191
rect 112 -101215 146 -101199
rect 112 -102207 146 -102191
rect -100 -102275 -84 -102241
rect 84 -102275 100 -102241
rect -100 -102383 -84 -102349
rect 84 -102383 100 -102349
rect -146 -102433 -112 -102417
rect -146 -103425 -112 -103409
rect 112 -102433 146 -102417
rect 112 -103425 146 -103409
rect -100 -103493 -84 -103459
rect 84 -103493 100 -103459
rect -100 -103601 -84 -103567
rect 84 -103601 100 -103567
rect -146 -103651 -112 -103635
rect -146 -104643 -112 -104627
rect 112 -103651 146 -103635
rect 112 -104643 146 -104627
rect -100 -104711 -84 -104677
rect 84 -104711 100 -104677
rect -100 -104819 -84 -104785
rect 84 -104819 100 -104785
rect -146 -104869 -112 -104853
rect -146 -105861 -112 -105845
rect 112 -104869 146 -104853
rect 112 -105861 146 -105845
rect -100 -105929 -84 -105895
rect 84 -105929 100 -105895
rect -100 -106037 -84 -106003
rect 84 -106037 100 -106003
rect -146 -106087 -112 -106071
rect -146 -107079 -112 -107063
rect 112 -106087 146 -106071
rect 112 -107079 146 -107063
rect -100 -107147 -84 -107113
rect 84 -107147 100 -107113
rect -100 -107255 -84 -107221
rect 84 -107255 100 -107221
rect -146 -107305 -112 -107289
rect -146 -108297 -112 -108281
rect 112 -107305 146 -107289
rect 112 -108297 146 -108281
rect -100 -108365 -84 -108331
rect 84 -108365 100 -108331
rect -100 -108473 -84 -108439
rect 84 -108473 100 -108439
rect -146 -108523 -112 -108507
rect -146 -109515 -112 -109499
rect 112 -108523 146 -108507
rect 112 -109515 146 -109499
rect -100 -109583 -84 -109549
rect 84 -109583 100 -109549
rect -100 -109691 -84 -109657
rect 84 -109691 100 -109657
rect -146 -109741 -112 -109725
rect -146 -110733 -112 -110717
rect 112 -109741 146 -109725
rect 112 -110733 146 -110717
rect -100 -110801 -84 -110767
rect 84 -110801 100 -110767
rect -100 -110909 -84 -110875
rect 84 -110909 100 -110875
rect -146 -110959 -112 -110943
rect -146 -111951 -112 -111935
rect 112 -110959 146 -110943
rect 112 -111951 146 -111935
rect -100 -112019 -84 -111985
rect 84 -112019 100 -111985
rect -100 -112127 -84 -112093
rect 84 -112127 100 -112093
rect -146 -112177 -112 -112161
rect -146 -113169 -112 -113153
rect 112 -112177 146 -112161
rect 112 -113169 146 -113153
rect -100 -113237 -84 -113203
rect 84 -113237 100 -113203
rect -100 -113345 -84 -113311
rect 84 -113345 100 -113311
rect -146 -113395 -112 -113379
rect -146 -114387 -112 -114371
rect 112 -113395 146 -113379
rect 112 -114387 146 -114371
rect -100 -114455 -84 -114421
rect 84 -114455 100 -114421
rect -100 -114563 -84 -114529
rect 84 -114563 100 -114529
rect -146 -114613 -112 -114597
rect -146 -115605 -112 -115589
rect 112 -114613 146 -114597
rect 112 -115605 146 -115589
rect -100 -115673 -84 -115639
rect 84 -115673 100 -115639
rect -100 -115781 -84 -115747
rect 84 -115781 100 -115747
rect -146 -115831 -112 -115815
rect -146 -116823 -112 -116807
rect 112 -115831 146 -115815
rect 112 -116823 146 -116807
rect -100 -116891 -84 -116857
rect 84 -116891 100 -116857
rect -100 -116999 -84 -116965
rect 84 -116999 100 -116965
rect -146 -117049 -112 -117033
rect -146 -118041 -112 -118025
rect 112 -117049 146 -117033
rect 112 -118041 146 -118025
rect -100 -118109 -84 -118075
rect 84 -118109 100 -118075
rect -100 -118217 -84 -118183
rect 84 -118217 100 -118183
rect -146 -118267 -112 -118251
rect -146 -119259 -112 -119243
rect 112 -118267 146 -118251
rect 112 -119259 146 -119243
rect -100 -119327 -84 -119293
rect 84 -119327 100 -119293
rect -100 -119435 -84 -119401
rect 84 -119435 100 -119401
rect -146 -119485 -112 -119469
rect -146 -120477 -112 -120461
rect 112 -119485 146 -119469
rect 112 -120477 146 -120461
rect -100 -120545 -84 -120511
rect 84 -120545 100 -120511
rect -100 -120653 -84 -120619
rect 84 -120653 100 -120619
rect -146 -120703 -112 -120687
rect -146 -121695 -112 -121679
rect 112 -120703 146 -120687
rect 112 -121695 146 -121679
rect -100 -121763 -84 -121729
rect 84 -121763 100 -121729
rect -280 -121867 -246 -121805
rect 246 -121867 280 -121805
rect -280 -121901 -184 -121867
rect 184 -121901 280 -121867
<< viali >>
rect -84 121729 84 121763
rect -146 120703 -112 121679
rect 112 120703 146 121679
rect -84 120619 84 120653
rect -84 120511 84 120545
rect -146 119485 -112 120461
rect 112 119485 146 120461
rect -84 119401 84 119435
rect -84 119293 84 119327
rect -146 118267 -112 119243
rect 112 118267 146 119243
rect -84 118183 84 118217
rect -84 118075 84 118109
rect -146 117049 -112 118025
rect 112 117049 146 118025
rect -84 116965 84 116999
rect -84 116857 84 116891
rect -146 115831 -112 116807
rect 112 115831 146 116807
rect -84 115747 84 115781
rect -84 115639 84 115673
rect -146 114613 -112 115589
rect 112 114613 146 115589
rect -84 114529 84 114563
rect -84 114421 84 114455
rect -146 113395 -112 114371
rect 112 113395 146 114371
rect -84 113311 84 113345
rect -84 113203 84 113237
rect -146 112177 -112 113153
rect 112 112177 146 113153
rect -84 112093 84 112127
rect -84 111985 84 112019
rect -146 110959 -112 111935
rect 112 110959 146 111935
rect -84 110875 84 110909
rect -84 110767 84 110801
rect -146 109741 -112 110717
rect 112 109741 146 110717
rect -84 109657 84 109691
rect -84 109549 84 109583
rect -146 108523 -112 109499
rect 112 108523 146 109499
rect -84 108439 84 108473
rect -84 108331 84 108365
rect -146 107305 -112 108281
rect 112 107305 146 108281
rect -84 107221 84 107255
rect -84 107113 84 107147
rect -146 106087 -112 107063
rect 112 106087 146 107063
rect -84 106003 84 106037
rect -84 105895 84 105929
rect -146 104869 -112 105845
rect 112 104869 146 105845
rect -84 104785 84 104819
rect -84 104677 84 104711
rect -146 103651 -112 104627
rect 112 103651 146 104627
rect -84 103567 84 103601
rect -84 103459 84 103493
rect -146 102433 -112 103409
rect 112 102433 146 103409
rect -84 102349 84 102383
rect -84 102241 84 102275
rect -146 101215 -112 102191
rect 112 101215 146 102191
rect -84 101131 84 101165
rect -84 101023 84 101057
rect -146 99997 -112 100973
rect 112 99997 146 100973
rect -84 99913 84 99947
rect -84 99805 84 99839
rect -146 98779 -112 99755
rect 112 98779 146 99755
rect -84 98695 84 98729
rect -84 98587 84 98621
rect -146 97561 -112 98537
rect 112 97561 146 98537
rect -84 97477 84 97511
rect -84 97369 84 97403
rect -146 96343 -112 97319
rect 112 96343 146 97319
rect -84 96259 84 96293
rect -84 96151 84 96185
rect -146 95125 -112 96101
rect 112 95125 146 96101
rect -84 95041 84 95075
rect -84 94933 84 94967
rect -146 93907 -112 94883
rect 112 93907 146 94883
rect -84 93823 84 93857
rect -84 93715 84 93749
rect -146 92689 -112 93665
rect 112 92689 146 93665
rect -84 92605 84 92639
rect -84 92497 84 92531
rect -146 91471 -112 92447
rect 112 91471 146 92447
rect -84 91387 84 91421
rect -84 91279 84 91313
rect -146 90253 -112 91229
rect 112 90253 146 91229
rect -84 90169 84 90203
rect -84 90061 84 90095
rect -146 89035 -112 90011
rect 112 89035 146 90011
rect -84 88951 84 88985
rect -84 88843 84 88877
rect -146 87817 -112 88793
rect 112 87817 146 88793
rect -84 87733 84 87767
rect -84 87625 84 87659
rect -146 86599 -112 87575
rect 112 86599 146 87575
rect -84 86515 84 86549
rect -84 86407 84 86441
rect -146 85381 -112 86357
rect 112 85381 146 86357
rect -84 85297 84 85331
rect -84 85189 84 85223
rect -146 84163 -112 85139
rect 112 84163 146 85139
rect -84 84079 84 84113
rect -84 83971 84 84005
rect -146 82945 -112 83921
rect 112 82945 146 83921
rect -84 82861 84 82895
rect -84 82753 84 82787
rect -146 81727 -112 82703
rect 112 81727 146 82703
rect -84 81643 84 81677
rect -84 81535 84 81569
rect -146 80509 -112 81485
rect 112 80509 146 81485
rect -84 80425 84 80459
rect -84 80317 84 80351
rect -146 79291 -112 80267
rect 112 79291 146 80267
rect -84 79207 84 79241
rect -84 79099 84 79133
rect -146 78073 -112 79049
rect 112 78073 146 79049
rect -84 77989 84 78023
rect -84 77881 84 77915
rect -146 76855 -112 77831
rect 112 76855 146 77831
rect -84 76771 84 76805
rect -84 76663 84 76697
rect -146 75637 -112 76613
rect 112 75637 146 76613
rect -84 75553 84 75587
rect -84 75445 84 75479
rect -146 74419 -112 75395
rect 112 74419 146 75395
rect -84 74335 84 74369
rect -84 74227 84 74261
rect -146 73201 -112 74177
rect 112 73201 146 74177
rect -84 73117 84 73151
rect -84 73009 84 73043
rect -146 71983 -112 72959
rect 112 71983 146 72959
rect -84 71899 84 71933
rect -84 71791 84 71825
rect -146 70765 -112 71741
rect 112 70765 146 71741
rect -84 70681 84 70715
rect -84 70573 84 70607
rect -146 69547 -112 70523
rect 112 69547 146 70523
rect -84 69463 84 69497
rect -84 69355 84 69389
rect -146 68329 -112 69305
rect 112 68329 146 69305
rect -84 68245 84 68279
rect -84 68137 84 68171
rect -146 67111 -112 68087
rect 112 67111 146 68087
rect -84 67027 84 67061
rect -84 66919 84 66953
rect -146 65893 -112 66869
rect 112 65893 146 66869
rect -84 65809 84 65843
rect -84 65701 84 65735
rect -146 64675 -112 65651
rect 112 64675 146 65651
rect -84 64591 84 64625
rect -84 64483 84 64517
rect -146 63457 -112 64433
rect 112 63457 146 64433
rect -84 63373 84 63407
rect -84 63265 84 63299
rect -146 62239 -112 63215
rect 112 62239 146 63215
rect -84 62155 84 62189
rect -84 62047 84 62081
rect -146 61021 -112 61997
rect 112 61021 146 61997
rect -84 60937 84 60971
rect -84 60829 84 60863
rect -146 59803 -112 60779
rect 112 59803 146 60779
rect -84 59719 84 59753
rect -84 59611 84 59645
rect -146 58585 -112 59561
rect 112 58585 146 59561
rect -84 58501 84 58535
rect -84 58393 84 58427
rect -146 57367 -112 58343
rect 112 57367 146 58343
rect -84 57283 84 57317
rect -84 57175 84 57209
rect -146 56149 -112 57125
rect 112 56149 146 57125
rect -84 56065 84 56099
rect -84 55957 84 55991
rect -146 54931 -112 55907
rect 112 54931 146 55907
rect -84 54847 84 54881
rect -84 54739 84 54773
rect -146 53713 -112 54689
rect 112 53713 146 54689
rect -84 53629 84 53663
rect -84 53521 84 53555
rect -146 52495 -112 53471
rect 112 52495 146 53471
rect -84 52411 84 52445
rect -84 52303 84 52337
rect -146 51277 -112 52253
rect 112 51277 146 52253
rect -84 51193 84 51227
rect -84 51085 84 51119
rect -146 50059 -112 51035
rect 112 50059 146 51035
rect -84 49975 84 50009
rect -84 49867 84 49901
rect -146 48841 -112 49817
rect 112 48841 146 49817
rect -84 48757 84 48791
rect -84 48649 84 48683
rect -146 47623 -112 48599
rect 112 47623 146 48599
rect -84 47539 84 47573
rect -84 47431 84 47465
rect -146 46405 -112 47381
rect 112 46405 146 47381
rect -84 46321 84 46355
rect -84 46213 84 46247
rect -146 45187 -112 46163
rect 112 45187 146 46163
rect -84 45103 84 45137
rect -84 44995 84 45029
rect -146 43969 -112 44945
rect 112 43969 146 44945
rect -84 43885 84 43919
rect -84 43777 84 43811
rect -146 42751 -112 43727
rect 112 42751 146 43727
rect -84 42667 84 42701
rect -84 42559 84 42593
rect -146 41533 -112 42509
rect 112 41533 146 42509
rect -84 41449 84 41483
rect -84 41341 84 41375
rect -146 40315 -112 41291
rect 112 40315 146 41291
rect -84 40231 84 40265
rect -84 40123 84 40157
rect -146 39097 -112 40073
rect 112 39097 146 40073
rect -84 39013 84 39047
rect -84 38905 84 38939
rect -146 37879 -112 38855
rect 112 37879 146 38855
rect -84 37795 84 37829
rect -84 37687 84 37721
rect -146 36661 -112 37637
rect 112 36661 146 37637
rect -84 36577 84 36611
rect -84 36469 84 36503
rect -146 35443 -112 36419
rect 112 35443 146 36419
rect -84 35359 84 35393
rect -84 35251 84 35285
rect -146 34225 -112 35201
rect 112 34225 146 35201
rect -84 34141 84 34175
rect -84 34033 84 34067
rect -146 33007 -112 33983
rect 112 33007 146 33983
rect -84 32923 84 32957
rect -84 32815 84 32849
rect -146 31789 -112 32765
rect 112 31789 146 32765
rect -84 31705 84 31739
rect -84 31597 84 31631
rect -146 30571 -112 31547
rect 112 30571 146 31547
rect -84 30487 84 30521
rect -84 30379 84 30413
rect -146 29353 -112 30329
rect 112 29353 146 30329
rect -84 29269 84 29303
rect -84 29161 84 29195
rect -146 28135 -112 29111
rect 112 28135 146 29111
rect -84 28051 84 28085
rect -84 27943 84 27977
rect -146 26917 -112 27893
rect 112 26917 146 27893
rect -84 26833 84 26867
rect -84 26725 84 26759
rect -146 25699 -112 26675
rect 112 25699 146 26675
rect -84 25615 84 25649
rect -84 25507 84 25541
rect -146 24481 -112 25457
rect 112 24481 146 25457
rect -84 24397 84 24431
rect -84 24289 84 24323
rect -146 23263 -112 24239
rect 112 23263 146 24239
rect -84 23179 84 23213
rect -84 23071 84 23105
rect -146 22045 -112 23021
rect 112 22045 146 23021
rect -84 21961 84 21995
rect -84 21853 84 21887
rect -146 20827 -112 21803
rect 112 20827 146 21803
rect -84 20743 84 20777
rect -84 20635 84 20669
rect -146 19609 -112 20585
rect 112 19609 146 20585
rect -84 19525 84 19559
rect -84 19417 84 19451
rect -146 18391 -112 19367
rect 112 18391 146 19367
rect -84 18307 84 18341
rect -84 18199 84 18233
rect -146 17173 -112 18149
rect 112 17173 146 18149
rect -84 17089 84 17123
rect -84 16981 84 17015
rect -146 15955 -112 16931
rect 112 15955 146 16931
rect -84 15871 84 15905
rect -84 15763 84 15797
rect -146 14737 -112 15713
rect 112 14737 146 15713
rect -84 14653 84 14687
rect -84 14545 84 14579
rect -146 13519 -112 14495
rect 112 13519 146 14495
rect -84 13435 84 13469
rect -84 13327 84 13361
rect -146 12301 -112 13277
rect 112 12301 146 13277
rect -84 12217 84 12251
rect -84 12109 84 12143
rect -146 11083 -112 12059
rect 112 11083 146 12059
rect -84 10999 84 11033
rect -84 10891 84 10925
rect -146 9865 -112 10841
rect 112 9865 146 10841
rect -84 9781 84 9815
rect -84 9673 84 9707
rect -146 8647 -112 9623
rect 112 8647 146 9623
rect -84 8563 84 8597
rect -84 8455 84 8489
rect -146 7429 -112 8405
rect 112 7429 146 8405
rect -84 7345 84 7379
rect -84 7237 84 7271
rect -146 6211 -112 7187
rect 112 6211 146 7187
rect -84 6127 84 6161
rect -84 6019 84 6053
rect -146 4993 -112 5969
rect 112 4993 146 5969
rect -84 4909 84 4943
rect -84 4801 84 4835
rect -146 3775 -112 4751
rect 112 3775 146 4751
rect -84 3691 84 3725
rect -84 3583 84 3617
rect -146 2557 -112 3533
rect 112 2557 146 3533
rect -84 2473 84 2507
rect -84 2365 84 2399
rect -146 1339 -112 2315
rect 112 1339 146 2315
rect -84 1255 84 1289
rect -84 1147 84 1181
rect -146 121 -112 1097
rect 112 121 146 1097
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -1097 -112 -121
rect 112 -1097 146 -121
rect -84 -1181 84 -1147
rect -84 -1289 84 -1255
rect -146 -2315 -112 -1339
rect 112 -2315 146 -1339
rect -84 -2399 84 -2365
rect -84 -2507 84 -2473
rect -146 -3533 -112 -2557
rect 112 -3533 146 -2557
rect -84 -3617 84 -3583
rect -84 -3725 84 -3691
rect -146 -4751 -112 -3775
rect 112 -4751 146 -3775
rect -84 -4835 84 -4801
rect -84 -4943 84 -4909
rect -146 -5969 -112 -4993
rect 112 -5969 146 -4993
rect -84 -6053 84 -6019
rect -84 -6161 84 -6127
rect -146 -7187 -112 -6211
rect 112 -7187 146 -6211
rect -84 -7271 84 -7237
rect -84 -7379 84 -7345
rect -146 -8405 -112 -7429
rect 112 -8405 146 -7429
rect -84 -8489 84 -8455
rect -84 -8597 84 -8563
rect -146 -9623 -112 -8647
rect 112 -9623 146 -8647
rect -84 -9707 84 -9673
rect -84 -9815 84 -9781
rect -146 -10841 -112 -9865
rect 112 -10841 146 -9865
rect -84 -10925 84 -10891
rect -84 -11033 84 -10999
rect -146 -12059 -112 -11083
rect 112 -12059 146 -11083
rect -84 -12143 84 -12109
rect -84 -12251 84 -12217
rect -146 -13277 -112 -12301
rect 112 -13277 146 -12301
rect -84 -13361 84 -13327
rect -84 -13469 84 -13435
rect -146 -14495 -112 -13519
rect 112 -14495 146 -13519
rect -84 -14579 84 -14545
rect -84 -14687 84 -14653
rect -146 -15713 -112 -14737
rect 112 -15713 146 -14737
rect -84 -15797 84 -15763
rect -84 -15905 84 -15871
rect -146 -16931 -112 -15955
rect 112 -16931 146 -15955
rect -84 -17015 84 -16981
rect -84 -17123 84 -17089
rect -146 -18149 -112 -17173
rect 112 -18149 146 -17173
rect -84 -18233 84 -18199
rect -84 -18341 84 -18307
rect -146 -19367 -112 -18391
rect 112 -19367 146 -18391
rect -84 -19451 84 -19417
rect -84 -19559 84 -19525
rect -146 -20585 -112 -19609
rect 112 -20585 146 -19609
rect -84 -20669 84 -20635
rect -84 -20777 84 -20743
rect -146 -21803 -112 -20827
rect 112 -21803 146 -20827
rect -84 -21887 84 -21853
rect -84 -21995 84 -21961
rect -146 -23021 -112 -22045
rect 112 -23021 146 -22045
rect -84 -23105 84 -23071
rect -84 -23213 84 -23179
rect -146 -24239 -112 -23263
rect 112 -24239 146 -23263
rect -84 -24323 84 -24289
rect -84 -24431 84 -24397
rect -146 -25457 -112 -24481
rect 112 -25457 146 -24481
rect -84 -25541 84 -25507
rect -84 -25649 84 -25615
rect -146 -26675 -112 -25699
rect 112 -26675 146 -25699
rect -84 -26759 84 -26725
rect -84 -26867 84 -26833
rect -146 -27893 -112 -26917
rect 112 -27893 146 -26917
rect -84 -27977 84 -27943
rect -84 -28085 84 -28051
rect -146 -29111 -112 -28135
rect 112 -29111 146 -28135
rect -84 -29195 84 -29161
rect -84 -29303 84 -29269
rect -146 -30329 -112 -29353
rect 112 -30329 146 -29353
rect -84 -30413 84 -30379
rect -84 -30521 84 -30487
rect -146 -31547 -112 -30571
rect 112 -31547 146 -30571
rect -84 -31631 84 -31597
rect -84 -31739 84 -31705
rect -146 -32765 -112 -31789
rect 112 -32765 146 -31789
rect -84 -32849 84 -32815
rect -84 -32957 84 -32923
rect -146 -33983 -112 -33007
rect 112 -33983 146 -33007
rect -84 -34067 84 -34033
rect -84 -34175 84 -34141
rect -146 -35201 -112 -34225
rect 112 -35201 146 -34225
rect -84 -35285 84 -35251
rect -84 -35393 84 -35359
rect -146 -36419 -112 -35443
rect 112 -36419 146 -35443
rect -84 -36503 84 -36469
rect -84 -36611 84 -36577
rect -146 -37637 -112 -36661
rect 112 -37637 146 -36661
rect -84 -37721 84 -37687
rect -84 -37829 84 -37795
rect -146 -38855 -112 -37879
rect 112 -38855 146 -37879
rect -84 -38939 84 -38905
rect -84 -39047 84 -39013
rect -146 -40073 -112 -39097
rect 112 -40073 146 -39097
rect -84 -40157 84 -40123
rect -84 -40265 84 -40231
rect -146 -41291 -112 -40315
rect 112 -41291 146 -40315
rect -84 -41375 84 -41341
rect -84 -41483 84 -41449
rect -146 -42509 -112 -41533
rect 112 -42509 146 -41533
rect -84 -42593 84 -42559
rect -84 -42701 84 -42667
rect -146 -43727 -112 -42751
rect 112 -43727 146 -42751
rect -84 -43811 84 -43777
rect -84 -43919 84 -43885
rect -146 -44945 -112 -43969
rect 112 -44945 146 -43969
rect -84 -45029 84 -44995
rect -84 -45137 84 -45103
rect -146 -46163 -112 -45187
rect 112 -46163 146 -45187
rect -84 -46247 84 -46213
rect -84 -46355 84 -46321
rect -146 -47381 -112 -46405
rect 112 -47381 146 -46405
rect -84 -47465 84 -47431
rect -84 -47573 84 -47539
rect -146 -48599 -112 -47623
rect 112 -48599 146 -47623
rect -84 -48683 84 -48649
rect -84 -48791 84 -48757
rect -146 -49817 -112 -48841
rect 112 -49817 146 -48841
rect -84 -49901 84 -49867
rect -84 -50009 84 -49975
rect -146 -51035 -112 -50059
rect 112 -51035 146 -50059
rect -84 -51119 84 -51085
rect -84 -51227 84 -51193
rect -146 -52253 -112 -51277
rect 112 -52253 146 -51277
rect -84 -52337 84 -52303
rect -84 -52445 84 -52411
rect -146 -53471 -112 -52495
rect 112 -53471 146 -52495
rect -84 -53555 84 -53521
rect -84 -53663 84 -53629
rect -146 -54689 -112 -53713
rect 112 -54689 146 -53713
rect -84 -54773 84 -54739
rect -84 -54881 84 -54847
rect -146 -55907 -112 -54931
rect 112 -55907 146 -54931
rect -84 -55991 84 -55957
rect -84 -56099 84 -56065
rect -146 -57125 -112 -56149
rect 112 -57125 146 -56149
rect -84 -57209 84 -57175
rect -84 -57317 84 -57283
rect -146 -58343 -112 -57367
rect 112 -58343 146 -57367
rect -84 -58427 84 -58393
rect -84 -58535 84 -58501
rect -146 -59561 -112 -58585
rect 112 -59561 146 -58585
rect -84 -59645 84 -59611
rect -84 -59753 84 -59719
rect -146 -60779 -112 -59803
rect 112 -60779 146 -59803
rect -84 -60863 84 -60829
rect -84 -60971 84 -60937
rect -146 -61997 -112 -61021
rect 112 -61997 146 -61021
rect -84 -62081 84 -62047
rect -84 -62189 84 -62155
rect -146 -63215 -112 -62239
rect 112 -63215 146 -62239
rect -84 -63299 84 -63265
rect -84 -63407 84 -63373
rect -146 -64433 -112 -63457
rect 112 -64433 146 -63457
rect -84 -64517 84 -64483
rect -84 -64625 84 -64591
rect -146 -65651 -112 -64675
rect 112 -65651 146 -64675
rect -84 -65735 84 -65701
rect -84 -65843 84 -65809
rect -146 -66869 -112 -65893
rect 112 -66869 146 -65893
rect -84 -66953 84 -66919
rect -84 -67061 84 -67027
rect -146 -68087 -112 -67111
rect 112 -68087 146 -67111
rect -84 -68171 84 -68137
rect -84 -68279 84 -68245
rect -146 -69305 -112 -68329
rect 112 -69305 146 -68329
rect -84 -69389 84 -69355
rect -84 -69497 84 -69463
rect -146 -70523 -112 -69547
rect 112 -70523 146 -69547
rect -84 -70607 84 -70573
rect -84 -70715 84 -70681
rect -146 -71741 -112 -70765
rect 112 -71741 146 -70765
rect -84 -71825 84 -71791
rect -84 -71933 84 -71899
rect -146 -72959 -112 -71983
rect 112 -72959 146 -71983
rect -84 -73043 84 -73009
rect -84 -73151 84 -73117
rect -146 -74177 -112 -73201
rect 112 -74177 146 -73201
rect -84 -74261 84 -74227
rect -84 -74369 84 -74335
rect -146 -75395 -112 -74419
rect 112 -75395 146 -74419
rect -84 -75479 84 -75445
rect -84 -75587 84 -75553
rect -146 -76613 -112 -75637
rect 112 -76613 146 -75637
rect -84 -76697 84 -76663
rect -84 -76805 84 -76771
rect -146 -77831 -112 -76855
rect 112 -77831 146 -76855
rect -84 -77915 84 -77881
rect -84 -78023 84 -77989
rect -146 -79049 -112 -78073
rect 112 -79049 146 -78073
rect -84 -79133 84 -79099
rect -84 -79241 84 -79207
rect -146 -80267 -112 -79291
rect 112 -80267 146 -79291
rect -84 -80351 84 -80317
rect -84 -80459 84 -80425
rect -146 -81485 -112 -80509
rect 112 -81485 146 -80509
rect -84 -81569 84 -81535
rect -84 -81677 84 -81643
rect -146 -82703 -112 -81727
rect 112 -82703 146 -81727
rect -84 -82787 84 -82753
rect -84 -82895 84 -82861
rect -146 -83921 -112 -82945
rect 112 -83921 146 -82945
rect -84 -84005 84 -83971
rect -84 -84113 84 -84079
rect -146 -85139 -112 -84163
rect 112 -85139 146 -84163
rect -84 -85223 84 -85189
rect -84 -85331 84 -85297
rect -146 -86357 -112 -85381
rect 112 -86357 146 -85381
rect -84 -86441 84 -86407
rect -84 -86549 84 -86515
rect -146 -87575 -112 -86599
rect 112 -87575 146 -86599
rect -84 -87659 84 -87625
rect -84 -87767 84 -87733
rect -146 -88793 -112 -87817
rect 112 -88793 146 -87817
rect -84 -88877 84 -88843
rect -84 -88985 84 -88951
rect -146 -90011 -112 -89035
rect 112 -90011 146 -89035
rect -84 -90095 84 -90061
rect -84 -90203 84 -90169
rect -146 -91229 -112 -90253
rect 112 -91229 146 -90253
rect -84 -91313 84 -91279
rect -84 -91421 84 -91387
rect -146 -92447 -112 -91471
rect 112 -92447 146 -91471
rect -84 -92531 84 -92497
rect -84 -92639 84 -92605
rect -146 -93665 -112 -92689
rect 112 -93665 146 -92689
rect -84 -93749 84 -93715
rect -84 -93857 84 -93823
rect -146 -94883 -112 -93907
rect 112 -94883 146 -93907
rect -84 -94967 84 -94933
rect -84 -95075 84 -95041
rect -146 -96101 -112 -95125
rect 112 -96101 146 -95125
rect -84 -96185 84 -96151
rect -84 -96293 84 -96259
rect -146 -97319 -112 -96343
rect 112 -97319 146 -96343
rect -84 -97403 84 -97369
rect -84 -97511 84 -97477
rect -146 -98537 -112 -97561
rect 112 -98537 146 -97561
rect -84 -98621 84 -98587
rect -84 -98729 84 -98695
rect -146 -99755 -112 -98779
rect 112 -99755 146 -98779
rect -84 -99839 84 -99805
rect -84 -99947 84 -99913
rect -146 -100973 -112 -99997
rect 112 -100973 146 -99997
rect -84 -101057 84 -101023
rect -84 -101165 84 -101131
rect -146 -102191 -112 -101215
rect 112 -102191 146 -101215
rect -84 -102275 84 -102241
rect -84 -102383 84 -102349
rect -146 -103409 -112 -102433
rect 112 -103409 146 -102433
rect -84 -103493 84 -103459
rect -84 -103601 84 -103567
rect -146 -104627 -112 -103651
rect 112 -104627 146 -103651
rect -84 -104711 84 -104677
rect -84 -104819 84 -104785
rect -146 -105845 -112 -104869
rect 112 -105845 146 -104869
rect -84 -105929 84 -105895
rect -84 -106037 84 -106003
rect -146 -107063 -112 -106087
rect 112 -107063 146 -106087
rect -84 -107147 84 -107113
rect -84 -107255 84 -107221
rect -146 -108281 -112 -107305
rect 112 -108281 146 -107305
rect -84 -108365 84 -108331
rect -84 -108473 84 -108439
rect -146 -109499 -112 -108523
rect 112 -109499 146 -108523
rect -84 -109583 84 -109549
rect -84 -109691 84 -109657
rect -146 -110717 -112 -109741
rect 112 -110717 146 -109741
rect -84 -110801 84 -110767
rect -84 -110909 84 -110875
rect -146 -111935 -112 -110959
rect 112 -111935 146 -110959
rect -84 -112019 84 -111985
rect -84 -112127 84 -112093
rect -146 -113153 -112 -112177
rect 112 -113153 146 -112177
rect -84 -113237 84 -113203
rect -84 -113345 84 -113311
rect -146 -114371 -112 -113395
rect 112 -114371 146 -113395
rect -84 -114455 84 -114421
rect -84 -114563 84 -114529
rect -146 -115589 -112 -114613
rect 112 -115589 146 -114613
rect -84 -115673 84 -115639
rect -84 -115781 84 -115747
rect -146 -116807 -112 -115831
rect 112 -116807 146 -115831
rect -84 -116891 84 -116857
rect -84 -116999 84 -116965
rect -146 -118025 -112 -117049
rect 112 -118025 146 -117049
rect -84 -118109 84 -118075
rect -84 -118217 84 -118183
rect -146 -119243 -112 -118267
rect 112 -119243 146 -118267
rect -84 -119327 84 -119293
rect -84 -119435 84 -119401
rect -146 -120461 -112 -119485
rect 112 -120461 146 -119485
rect -84 -120545 84 -120511
rect -84 -120653 84 -120619
rect -146 -121679 -112 -120703
rect 112 -121679 146 -120703
rect -84 -121763 84 -121729
<< metal1 >>
rect -96 121763 96 121769
rect -96 121729 -84 121763
rect 84 121729 96 121763
rect -96 121723 96 121729
rect -152 121679 -106 121691
rect -152 120703 -146 121679
rect -112 120703 -106 121679
rect -152 120691 -106 120703
rect 106 121679 152 121691
rect 106 120703 112 121679
rect 146 120703 152 121679
rect 106 120691 152 120703
rect -96 120653 96 120659
rect -96 120619 -84 120653
rect 84 120619 96 120653
rect -96 120613 96 120619
rect -96 120545 96 120551
rect -96 120511 -84 120545
rect 84 120511 96 120545
rect -96 120505 96 120511
rect -152 120461 -106 120473
rect -152 119485 -146 120461
rect -112 119485 -106 120461
rect -152 119473 -106 119485
rect 106 120461 152 120473
rect 106 119485 112 120461
rect 146 119485 152 120461
rect 106 119473 152 119485
rect -96 119435 96 119441
rect -96 119401 -84 119435
rect 84 119401 96 119435
rect -96 119395 96 119401
rect -96 119327 96 119333
rect -96 119293 -84 119327
rect 84 119293 96 119327
rect -96 119287 96 119293
rect -152 119243 -106 119255
rect -152 118267 -146 119243
rect -112 118267 -106 119243
rect -152 118255 -106 118267
rect 106 119243 152 119255
rect 106 118267 112 119243
rect 146 118267 152 119243
rect 106 118255 152 118267
rect -96 118217 96 118223
rect -96 118183 -84 118217
rect 84 118183 96 118217
rect -96 118177 96 118183
rect -96 118109 96 118115
rect -96 118075 -84 118109
rect 84 118075 96 118109
rect -96 118069 96 118075
rect -152 118025 -106 118037
rect -152 117049 -146 118025
rect -112 117049 -106 118025
rect -152 117037 -106 117049
rect 106 118025 152 118037
rect 106 117049 112 118025
rect 146 117049 152 118025
rect 106 117037 152 117049
rect -96 116999 96 117005
rect -96 116965 -84 116999
rect 84 116965 96 116999
rect -96 116959 96 116965
rect -96 116891 96 116897
rect -96 116857 -84 116891
rect 84 116857 96 116891
rect -96 116851 96 116857
rect -152 116807 -106 116819
rect -152 115831 -146 116807
rect -112 115831 -106 116807
rect -152 115819 -106 115831
rect 106 116807 152 116819
rect 106 115831 112 116807
rect 146 115831 152 116807
rect 106 115819 152 115831
rect -96 115781 96 115787
rect -96 115747 -84 115781
rect 84 115747 96 115781
rect -96 115741 96 115747
rect -96 115673 96 115679
rect -96 115639 -84 115673
rect 84 115639 96 115673
rect -96 115633 96 115639
rect -152 115589 -106 115601
rect -152 114613 -146 115589
rect -112 114613 -106 115589
rect -152 114601 -106 114613
rect 106 115589 152 115601
rect 106 114613 112 115589
rect 146 114613 152 115589
rect 106 114601 152 114613
rect -96 114563 96 114569
rect -96 114529 -84 114563
rect 84 114529 96 114563
rect -96 114523 96 114529
rect -96 114455 96 114461
rect -96 114421 -84 114455
rect 84 114421 96 114455
rect -96 114415 96 114421
rect -152 114371 -106 114383
rect -152 113395 -146 114371
rect -112 113395 -106 114371
rect -152 113383 -106 113395
rect 106 114371 152 114383
rect 106 113395 112 114371
rect 146 113395 152 114371
rect 106 113383 152 113395
rect -96 113345 96 113351
rect -96 113311 -84 113345
rect 84 113311 96 113345
rect -96 113305 96 113311
rect -96 113237 96 113243
rect -96 113203 -84 113237
rect 84 113203 96 113237
rect -96 113197 96 113203
rect -152 113153 -106 113165
rect -152 112177 -146 113153
rect -112 112177 -106 113153
rect -152 112165 -106 112177
rect 106 113153 152 113165
rect 106 112177 112 113153
rect 146 112177 152 113153
rect 106 112165 152 112177
rect -96 112127 96 112133
rect -96 112093 -84 112127
rect 84 112093 96 112127
rect -96 112087 96 112093
rect -96 112019 96 112025
rect -96 111985 -84 112019
rect 84 111985 96 112019
rect -96 111979 96 111985
rect -152 111935 -106 111947
rect -152 110959 -146 111935
rect -112 110959 -106 111935
rect -152 110947 -106 110959
rect 106 111935 152 111947
rect 106 110959 112 111935
rect 146 110959 152 111935
rect 106 110947 152 110959
rect -96 110909 96 110915
rect -96 110875 -84 110909
rect 84 110875 96 110909
rect -96 110869 96 110875
rect -96 110801 96 110807
rect -96 110767 -84 110801
rect 84 110767 96 110801
rect -96 110761 96 110767
rect -152 110717 -106 110729
rect -152 109741 -146 110717
rect -112 109741 -106 110717
rect -152 109729 -106 109741
rect 106 110717 152 110729
rect 106 109741 112 110717
rect 146 109741 152 110717
rect 106 109729 152 109741
rect -96 109691 96 109697
rect -96 109657 -84 109691
rect 84 109657 96 109691
rect -96 109651 96 109657
rect -96 109583 96 109589
rect -96 109549 -84 109583
rect 84 109549 96 109583
rect -96 109543 96 109549
rect -152 109499 -106 109511
rect -152 108523 -146 109499
rect -112 108523 -106 109499
rect -152 108511 -106 108523
rect 106 109499 152 109511
rect 106 108523 112 109499
rect 146 108523 152 109499
rect 106 108511 152 108523
rect -96 108473 96 108479
rect -96 108439 -84 108473
rect 84 108439 96 108473
rect -96 108433 96 108439
rect -96 108365 96 108371
rect -96 108331 -84 108365
rect 84 108331 96 108365
rect -96 108325 96 108331
rect -152 108281 -106 108293
rect -152 107305 -146 108281
rect -112 107305 -106 108281
rect -152 107293 -106 107305
rect 106 108281 152 108293
rect 106 107305 112 108281
rect 146 107305 152 108281
rect 106 107293 152 107305
rect -96 107255 96 107261
rect -96 107221 -84 107255
rect 84 107221 96 107255
rect -96 107215 96 107221
rect -96 107147 96 107153
rect -96 107113 -84 107147
rect 84 107113 96 107147
rect -96 107107 96 107113
rect -152 107063 -106 107075
rect -152 106087 -146 107063
rect -112 106087 -106 107063
rect -152 106075 -106 106087
rect 106 107063 152 107075
rect 106 106087 112 107063
rect 146 106087 152 107063
rect 106 106075 152 106087
rect -96 106037 96 106043
rect -96 106003 -84 106037
rect 84 106003 96 106037
rect -96 105997 96 106003
rect -96 105929 96 105935
rect -96 105895 -84 105929
rect 84 105895 96 105929
rect -96 105889 96 105895
rect -152 105845 -106 105857
rect -152 104869 -146 105845
rect -112 104869 -106 105845
rect -152 104857 -106 104869
rect 106 105845 152 105857
rect 106 104869 112 105845
rect 146 104869 152 105845
rect 106 104857 152 104869
rect -96 104819 96 104825
rect -96 104785 -84 104819
rect 84 104785 96 104819
rect -96 104779 96 104785
rect -96 104711 96 104717
rect -96 104677 -84 104711
rect 84 104677 96 104711
rect -96 104671 96 104677
rect -152 104627 -106 104639
rect -152 103651 -146 104627
rect -112 103651 -106 104627
rect -152 103639 -106 103651
rect 106 104627 152 104639
rect 106 103651 112 104627
rect 146 103651 152 104627
rect 106 103639 152 103651
rect -96 103601 96 103607
rect -96 103567 -84 103601
rect 84 103567 96 103601
rect -96 103561 96 103567
rect -96 103493 96 103499
rect -96 103459 -84 103493
rect 84 103459 96 103493
rect -96 103453 96 103459
rect -152 103409 -106 103421
rect -152 102433 -146 103409
rect -112 102433 -106 103409
rect -152 102421 -106 102433
rect 106 103409 152 103421
rect 106 102433 112 103409
rect 146 102433 152 103409
rect 106 102421 152 102433
rect -96 102383 96 102389
rect -96 102349 -84 102383
rect 84 102349 96 102383
rect -96 102343 96 102349
rect -96 102275 96 102281
rect -96 102241 -84 102275
rect 84 102241 96 102275
rect -96 102235 96 102241
rect -152 102191 -106 102203
rect -152 101215 -146 102191
rect -112 101215 -106 102191
rect -152 101203 -106 101215
rect 106 102191 152 102203
rect 106 101215 112 102191
rect 146 101215 152 102191
rect 106 101203 152 101215
rect -96 101165 96 101171
rect -96 101131 -84 101165
rect 84 101131 96 101165
rect -96 101125 96 101131
rect -96 101057 96 101063
rect -96 101023 -84 101057
rect 84 101023 96 101057
rect -96 101017 96 101023
rect -152 100973 -106 100985
rect -152 99997 -146 100973
rect -112 99997 -106 100973
rect -152 99985 -106 99997
rect 106 100973 152 100985
rect 106 99997 112 100973
rect 146 99997 152 100973
rect 106 99985 152 99997
rect -96 99947 96 99953
rect -96 99913 -84 99947
rect 84 99913 96 99947
rect -96 99907 96 99913
rect -96 99839 96 99845
rect -96 99805 -84 99839
rect 84 99805 96 99839
rect -96 99799 96 99805
rect -152 99755 -106 99767
rect -152 98779 -146 99755
rect -112 98779 -106 99755
rect -152 98767 -106 98779
rect 106 99755 152 99767
rect 106 98779 112 99755
rect 146 98779 152 99755
rect 106 98767 152 98779
rect -96 98729 96 98735
rect -96 98695 -84 98729
rect 84 98695 96 98729
rect -96 98689 96 98695
rect -96 98621 96 98627
rect -96 98587 -84 98621
rect 84 98587 96 98621
rect -96 98581 96 98587
rect -152 98537 -106 98549
rect -152 97561 -146 98537
rect -112 97561 -106 98537
rect -152 97549 -106 97561
rect 106 98537 152 98549
rect 106 97561 112 98537
rect 146 97561 152 98537
rect 106 97549 152 97561
rect -96 97511 96 97517
rect -96 97477 -84 97511
rect 84 97477 96 97511
rect -96 97471 96 97477
rect -96 97403 96 97409
rect -96 97369 -84 97403
rect 84 97369 96 97403
rect -96 97363 96 97369
rect -152 97319 -106 97331
rect -152 96343 -146 97319
rect -112 96343 -106 97319
rect -152 96331 -106 96343
rect 106 97319 152 97331
rect 106 96343 112 97319
rect 146 96343 152 97319
rect 106 96331 152 96343
rect -96 96293 96 96299
rect -96 96259 -84 96293
rect 84 96259 96 96293
rect -96 96253 96 96259
rect -96 96185 96 96191
rect -96 96151 -84 96185
rect 84 96151 96 96185
rect -96 96145 96 96151
rect -152 96101 -106 96113
rect -152 95125 -146 96101
rect -112 95125 -106 96101
rect -152 95113 -106 95125
rect 106 96101 152 96113
rect 106 95125 112 96101
rect 146 95125 152 96101
rect 106 95113 152 95125
rect -96 95075 96 95081
rect -96 95041 -84 95075
rect 84 95041 96 95075
rect -96 95035 96 95041
rect -96 94967 96 94973
rect -96 94933 -84 94967
rect 84 94933 96 94967
rect -96 94927 96 94933
rect -152 94883 -106 94895
rect -152 93907 -146 94883
rect -112 93907 -106 94883
rect -152 93895 -106 93907
rect 106 94883 152 94895
rect 106 93907 112 94883
rect 146 93907 152 94883
rect 106 93895 152 93907
rect -96 93857 96 93863
rect -96 93823 -84 93857
rect 84 93823 96 93857
rect -96 93817 96 93823
rect -96 93749 96 93755
rect -96 93715 -84 93749
rect 84 93715 96 93749
rect -96 93709 96 93715
rect -152 93665 -106 93677
rect -152 92689 -146 93665
rect -112 92689 -106 93665
rect -152 92677 -106 92689
rect 106 93665 152 93677
rect 106 92689 112 93665
rect 146 92689 152 93665
rect 106 92677 152 92689
rect -96 92639 96 92645
rect -96 92605 -84 92639
rect 84 92605 96 92639
rect -96 92599 96 92605
rect -96 92531 96 92537
rect -96 92497 -84 92531
rect 84 92497 96 92531
rect -96 92491 96 92497
rect -152 92447 -106 92459
rect -152 91471 -146 92447
rect -112 91471 -106 92447
rect -152 91459 -106 91471
rect 106 92447 152 92459
rect 106 91471 112 92447
rect 146 91471 152 92447
rect 106 91459 152 91471
rect -96 91421 96 91427
rect -96 91387 -84 91421
rect 84 91387 96 91421
rect -96 91381 96 91387
rect -96 91313 96 91319
rect -96 91279 -84 91313
rect 84 91279 96 91313
rect -96 91273 96 91279
rect -152 91229 -106 91241
rect -152 90253 -146 91229
rect -112 90253 -106 91229
rect -152 90241 -106 90253
rect 106 91229 152 91241
rect 106 90253 112 91229
rect 146 90253 152 91229
rect 106 90241 152 90253
rect -96 90203 96 90209
rect -96 90169 -84 90203
rect 84 90169 96 90203
rect -96 90163 96 90169
rect -96 90095 96 90101
rect -96 90061 -84 90095
rect 84 90061 96 90095
rect -96 90055 96 90061
rect -152 90011 -106 90023
rect -152 89035 -146 90011
rect -112 89035 -106 90011
rect -152 89023 -106 89035
rect 106 90011 152 90023
rect 106 89035 112 90011
rect 146 89035 152 90011
rect 106 89023 152 89035
rect -96 88985 96 88991
rect -96 88951 -84 88985
rect 84 88951 96 88985
rect -96 88945 96 88951
rect -96 88877 96 88883
rect -96 88843 -84 88877
rect 84 88843 96 88877
rect -96 88837 96 88843
rect -152 88793 -106 88805
rect -152 87817 -146 88793
rect -112 87817 -106 88793
rect -152 87805 -106 87817
rect 106 88793 152 88805
rect 106 87817 112 88793
rect 146 87817 152 88793
rect 106 87805 152 87817
rect -96 87767 96 87773
rect -96 87733 -84 87767
rect 84 87733 96 87767
rect -96 87727 96 87733
rect -96 87659 96 87665
rect -96 87625 -84 87659
rect 84 87625 96 87659
rect -96 87619 96 87625
rect -152 87575 -106 87587
rect -152 86599 -146 87575
rect -112 86599 -106 87575
rect -152 86587 -106 86599
rect 106 87575 152 87587
rect 106 86599 112 87575
rect 146 86599 152 87575
rect 106 86587 152 86599
rect -96 86549 96 86555
rect -96 86515 -84 86549
rect 84 86515 96 86549
rect -96 86509 96 86515
rect -96 86441 96 86447
rect -96 86407 -84 86441
rect 84 86407 96 86441
rect -96 86401 96 86407
rect -152 86357 -106 86369
rect -152 85381 -146 86357
rect -112 85381 -106 86357
rect -152 85369 -106 85381
rect 106 86357 152 86369
rect 106 85381 112 86357
rect 146 85381 152 86357
rect 106 85369 152 85381
rect -96 85331 96 85337
rect -96 85297 -84 85331
rect 84 85297 96 85331
rect -96 85291 96 85297
rect -96 85223 96 85229
rect -96 85189 -84 85223
rect 84 85189 96 85223
rect -96 85183 96 85189
rect -152 85139 -106 85151
rect -152 84163 -146 85139
rect -112 84163 -106 85139
rect -152 84151 -106 84163
rect 106 85139 152 85151
rect 106 84163 112 85139
rect 146 84163 152 85139
rect 106 84151 152 84163
rect -96 84113 96 84119
rect -96 84079 -84 84113
rect 84 84079 96 84113
rect -96 84073 96 84079
rect -96 84005 96 84011
rect -96 83971 -84 84005
rect 84 83971 96 84005
rect -96 83965 96 83971
rect -152 83921 -106 83933
rect -152 82945 -146 83921
rect -112 82945 -106 83921
rect -152 82933 -106 82945
rect 106 83921 152 83933
rect 106 82945 112 83921
rect 146 82945 152 83921
rect 106 82933 152 82945
rect -96 82895 96 82901
rect -96 82861 -84 82895
rect 84 82861 96 82895
rect -96 82855 96 82861
rect -96 82787 96 82793
rect -96 82753 -84 82787
rect 84 82753 96 82787
rect -96 82747 96 82753
rect -152 82703 -106 82715
rect -152 81727 -146 82703
rect -112 81727 -106 82703
rect -152 81715 -106 81727
rect 106 82703 152 82715
rect 106 81727 112 82703
rect 146 81727 152 82703
rect 106 81715 152 81727
rect -96 81677 96 81683
rect -96 81643 -84 81677
rect 84 81643 96 81677
rect -96 81637 96 81643
rect -96 81569 96 81575
rect -96 81535 -84 81569
rect 84 81535 96 81569
rect -96 81529 96 81535
rect -152 81485 -106 81497
rect -152 80509 -146 81485
rect -112 80509 -106 81485
rect -152 80497 -106 80509
rect 106 81485 152 81497
rect 106 80509 112 81485
rect 146 80509 152 81485
rect 106 80497 152 80509
rect -96 80459 96 80465
rect -96 80425 -84 80459
rect 84 80425 96 80459
rect -96 80419 96 80425
rect -96 80351 96 80357
rect -96 80317 -84 80351
rect 84 80317 96 80351
rect -96 80311 96 80317
rect -152 80267 -106 80279
rect -152 79291 -146 80267
rect -112 79291 -106 80267
rect -152 79279 -106 79291
rect 106 80267 152 80279
rect 106 79291 112 80267
rect 146 79291 152 80267
rect 106 79279 152 79291
rect -96 79241 96 79247
rect -96 79207 -84 79241
rect 84 79207 96 79241
rect -96 79201 96 79207
rect -96 79133 96 79139
rect -96 79099 -84 79133
rect 84 79099 96 79133
rect -96 79093 96 79099
rect -152 79049 -106 79061
rect -152 78073 -146 79049
rect -112 78073 -106 79049
rect -152 78061 -106 78073
rect 106 79049 152 79061
rect 106 78073 112 79049
rect 146 78073 152 79049
rect 106 78061 152 78073
rect -96 78023 96 78029
rect -96 77989 -84 78023
rect 84 77989 96 78023
rect -96 77983 96 77989
rect -96 77915 96 77921
rect -96 77881 -84 77915
rect 84 77881 96 77915
rect -96 77875 96 77881
rect -152 77831 -106 77843
rect -152 76855 -146 77831
rect -112 76855 -106 77831
rect -152 76843 -106 76855
rect 106 77831 152 77843
rect 106 76855 112 77831
rect 146 76855 152 77831
rect 106 76843 152 76855
rect -96 76805 96 76811
rect -96 76771 -84 76805
rect 84 76771 96 76805
rect -96 76765 96 76771
rect -96 76697 96 76703
rect -96 76663 -84 76697
rect 84 76663 96 76697
rect -96 76657 96 76663
rect -152 76613 -106 76625
rect -152 75637 -146 76613
rect -112 75637 -106 76613
rect -152 75625 -106 75637
rect 106 76613 152 76625
rect 106 75637 112 76613
rect 146 75637 152 76613
rect 106 75625 152 75637
rect -96 75587 96 75593
rect -96 75553 -84 75587
rect 84 75553 96 75587
rect -96 75547 96 75553
rect -96 75479 96 75485
rect -96 75445 -84 75479
rect 84 75445 96 75479
rect -96 75439 96 75445
rect -152 75395 -106 75407
rect -152 74419 -146 75395
rect -112 74419 -106 75395
rect -152 74407 -106 74419
rect 106 75395 152 75407
rect 106 74419 112 75395
rect 146 74419 152 75395
rect 106 74407 152 74419
rect -96 74369 96 74375
rect -96 74335 -84 74369
rect 84 74335 96 74369
rect -96 74329 96 74335
rect -96 74261 96 74267
rect -96 74227 -84 74261
rect 84 74227 96 74261
rect -96 74221 96 74227
rect -152 74177 -106 74189
rect -152 73201 -146 74177
rect -112 73201 -106 74177
rect -152 73189 -106 73201
rect 106 74177 152 74189
rect 106 73201 112 74177
rect 146 73201 152 74177
rect 106 73189 152 73201
rect -96 73151 96 73157
rect -96 73117 -84 73151
rect 84 73117 96 73151
rect -96 73111 96 73117
rect -96 73043 96 73049
rect -96 73009 -84 73043
rect 84 73009 96 73043
rect -96 73003 96 73009
rect -152 72959 -106 72971
rect -152 71983 -146 72959
rect -112 71983 -106 72959
rect -152 71971 -106 71983
rect 106 72959 152 72971
rect 106 71983 112 72959
rect 146 71983 152 72959
rect 106 71971 152 71983
rect -96 71933 96 71939
rect -96 71899 -84 71933
rect 84 71899 96 71933
rect -96 71893 96 71899
rect -96 71825 96 71831
rect -96 71791 -84 71825
rect 84 71791 96 71825
rect -96 71785 96 71791
rect -152 71741 -106 71753
rect -152 70765 -146 71741
rect -112 70765 -106 71741
rect -152 70753 -106 70765
rect 106 71741 152 71753
rect 106 70765 112 71741
rect 146 70765 152 71741
rect 106 70753 152 70765
rect -96 70715 96 70721
rect -96 70681 -84 70715
rect 84 70681 96 70715
rect -96 70675 96 70681
rect -96 70607 96 70613
rect -96 70573 -84 70607
rect 84 70573 96 70607
rect -96 70567 96 70573
rect -152 70523 -106 70535
rect -152 69547 -146 70523
rect -112 69547 -106 70523
rect -152 69535 -106 69547
rect 106 70523 152 70535
rect 106 69547 112 70523
rect 146 69547 152 70523
rect 106 69535 152 69547
rect -96 69497 96 69503
rect -96 69463 -84 69497
rect 84 69463 96 69497
rect -96 69457 96 69463
rect -96 69389 96 69395
rect -96 69355 -84 69389
rect 84 69355 96 69389
rect -96 69349 96 69355
rect -152 69305 -106 69317
rect -152 68329 -146 69305
rect -112 68329 -106 69305
rect -152 68317 -106 68329
rect 106 69305 152 69317
rect 106 68329 112 69305
rect 146 68329 152 69305
rect 106 68317 152 68329
rect -96 68279 96 68285
rect -96 68245 -84 68279
rect 84 68245 96 68279
rect -96 68239 96 68245
rect -96 68171 96 68177
rect -96 68137 -84 68171
rect 84 68137 96 68171
rect -96 68131 96 68137
rect -152 68087 -106 68099
rect -152 67111 -146 68087
rect -112 67111 -106 68087
rect -152 67099 -106 67111
rect 106 68087 152 68099
rect 106 67111 112 68087
rect 146 67111 152 68087
rect 106 67099 152 67111
rect -96 67061 96 67067
rect -96 67027 -84 67061
rect 84 67027 96 67061
rect -96 67021 96 67027
rect -96 66953 96 66959
rect -96 66919 -84 66953
rect 84 66919 96 66953
rect -96 66913 96 66919
rect -152 66869 -106 66881
rect -152 65893 -146 66869
rect -112 65893 -106 66869
rect -152 65881 -106 65893
rect 106 66869 152 66881
rect 106 65893 112 66869
rect 146 65893 152 66869
rect 106 65881 152 65893
rect -96 65843 96 65849
rect -96 65809 -84 65843
rect 84 65809 96 65843
rect -96 65803 96 65809
rect -96 65735 96 65741
rect -96 65701 -84 65735
rect 84 65701 96 65735
rect -96 65695 96 65701
rect -152 65651 -106 65663
rect -152 64675 -146 65651
rect -112 64675 -106 65651
rect -152 64663 -106 64675
rect 106 65651 152 65663
rect 106 64675 112 65651
rect 146 64675 152 65651
rect 106 64663 152 64675
rect -96 64625 96 64631
rect -96 64591 -84 64625
rect 84 64591 96 64625
rect -96 64585 96 64591
rect -96 64517 96 64523
rect -96 64483 -84 64517
rect 84 64483 96 64517
rect -96 64477 96 64483
rect -152 64433 -106 64445
rect -152 63457 -146 64433
rect -112 63457 -106 64433
rect -152 63445 -106 63457
rect 106 64433 152 64445
rect 106 63457 112 64433
rect 146 63457 152 64433
rect 106 63445 152 63457
rect -96 63407 96 63413
rect -96 63373 -84 63407
rect 84 63373 96 63407
rect -96 63367 96 63373
rect -96 63299 96 63305
rect -96 63265 -84 63299
rect 84 63265 96 63299
rect -96 63259 96 63265
rect -152 63215 -106 63227
rect -152 62239 -146 63215
rect -112 62239 -106 63215
rect -152 62227 -106 62239
rect 106 63215 152 63227
rect 106 62239 112 63215
rect 146 62239 152 63215
rect 106 62227 152 62239
rect -96 62189 96 62195
rect -96 62155 -84 62189
rect 84 62155 96 62189
rect -96 62149 96 62155
rect -96 62081 96 62087
rect -96 62047 -84 62081
rect 84 62047 96 62081
rect -96 62041 96 62047
rect -152 61997 -106 62009
rect -152 61021 -146 61997
rect -112 61021 -106 61997
rect -152 61009 -106 61021
rect 106 61997 152 62009
rect 106 61021 112 61997
rect 146 61021 152 61997
rect 106 61009 152 61021
rect -96 60971 96 60977
rect -96 60937 -84 60971
rect 84 60937 96 60971
rect -96 60931 96 60937
rect -96 60863 96 60869
rect -96 60829 -84 60863
rect 84 60829 96 60863
rect -96 60823 96 60829
rect -152 60779 -106 60791
rect -152 59803 -146 60779
rect -112 59803 -106 60779
rect -152 59791 -106 59803
rect 106 60779 152 60791
rect 106 59803 112 60779
rect 146 59803 152 60779
rect 106 59791 152 59803
rect -96 59753 96 59759
rect -96 59719 -84 59753
rect 84 59719 96 59753
rect -96 59713 96 59719
rect -96 59645 96 59651
rect -96 59611 -84 59645
rect 84 59611 96 59645
rect -96 59605 96 59611
rect -152 59561 -106 59573
rect -152 58585 -146 59561
rect -112 58585 -106 59561
rect -152 58573 -106 58585
rect 106 59561 152 59573
rect 106 58585 112 59561
rect 146 58585 152 59561
rect 106 58573 152 58585
rect -96 58535 96 58541
rect -96 58501 -84 58535
rect 84 58501 96 58535
rect -96 58495 96 58501
rect -96 58427 96 58433
rect -96 58393 -84 58427
rect 84 58393 96 58427
rect -96 58387 96 58393
rect -152 58343 -106 58355
rect -152 57367 -146 58343
rect -112 57367 -106 58343
rect -152 57355 -106 57367
rect 106 58343 152 58355
rect 106 57367 112 58343
rect 146 57367 152 58343
rect 106 57355 152 57367
rect -96 57317 96 57323
rect -96 57283 -84 57317
rect 84 57283 96 57317
rect -96 57277 96 57283
rect -96 57209 96 57215
rect -96 57175 -84 57209
rect 84 57175 96 57209
rect -96 57169 96 57175
rect -152 57125 -106 57137
rect -152 56149 -146 57125
rect -112 56149 -106 57125
rect -152 56137 -106 56149
rect 106 57125 152 57137
rect 106 56149 112 57125
rect 146 56149 152 57125
rect 106 56137 152 56149
rect -96 56099 96 56105
rect -96 56065 -84 56099
rect 84 56065 96 56099
rect -96 56059 96 56065
rect -96 55991 96 55997
rect -96 55957 -84 55991
rect 84 55957 96 55991
rect -96 55951 96 55957
rect -152 55907 -106 55919
rect -152 54931 -146 55907
rect -112 54931 -106 55907
rect -152 54919 -106 54931
rect 106 55907 152 55919
rect 106 54931 112 55907
rect 146 54931 152 55907
rect 106 54919 152 54931
rect -96 54881 96 54887
rect -96 54847 -84 54881
rect 84 54847 96 54881
rect -96 54841 96 54847
rect -96 54773 96 54779
rect -96 54739 -84 54773
rect 84 54739 96 54773
rect -96 54733 96 54739
rect -152 54689 -106 54701
rect -152 53713 -146 54689
rect -112 53713 -106 54689
rect -152 53701 -106 53713
rect 106 54689 152 54701
rect 106 53713 112 54689
rect 146 53713 152 54689
rect 106 53701 152 53713
rect -96 53663 96 53669
rect -96 53629 -84 53663
rect 84 53629 96 53663
rect -96 53623 96 53629
rect -96 53555 96 53561
rect -96 53521 -84 53555
rect 84 53521 96 53555
rect -96 53515 96 53521
rect -152 53471 -106 53483
rect -152 52495 -146 53471
rect -112 52495 -106 53471
rect -152 52483 -106 52495
rect 106 53471 152 53483
rect 106 52495 112 53471
rect 146 52495 152 53471
rect 106 52483 152 52495
rect -96 52445 96 52451
rect -96 52411 -84 52445
rect 84 52411 96 52445
rect -96 52405 96 52411
rect -96 52337 96 52343
rect -96 52303 -84 52337
rect 84 52303 96 52337
rect -96 52297 96 52303
rect -152 52253 -106 52265
rect -152 51277 -146 52253
rect -112 51277 -106 52253
rect -152 51265 -106 51277
rect 106 52253 152 52265
rect 106 51277 112 52253
rect 146 51277 152 52253
rect 106 51265 152 51277
rect -96 51227 96 51233
rect -96 51193 -84 51227
rect 84 51193 96 51227
rect -96 51187 96 51193
rect -96 51119 96 51125
rect -96 51085 -84 51119
rect 84 51085 96 51119
rect -96 51079 96 51085
rect -152 51035 -106 51047
rect -152 50059 -146 51035
rect -112 50059 -106 51035
rect -152 50047 -106 50059
rect 106 51035 152 51047
rect 106 50059 112 51035
rect 146 50059 152 51035
rect 106 50047 152 50059
rect -96 50009 96 50015
rect -96 49975 -84 50009
rect 84 49975 96 50009
rect -96 49969 96 49975
rect -96 49901 96 49907
rect -96 49867 -84 49901
rect 84 49867 96 49901
rect -96 49861 96 49867
rect -152 49817 -106 49829
rect -152 48841 -146 49817
rect -112 48841 -106 49817
rect -152 48829 -106 48841
rect 106 49817 152 49829
rect 106 48841 112 49817
rect 146 48841 152 49817
rect 106 48829 152 48841
rect -96 48791 96 48797
rect -96 48757 -84 48791
rect 84 48757 96 48791
rect -96 48751 96 48757
rect -96 48683 96 48689
rect -96 48649 -84 48683
rect 84 48649 96 48683
rect -96 48643 96 48649
rect -152 48599 -106 48611
rect -152 47623 -146 48599
rect -112 47623 -106 48599
rect -152 47611 -106 47623
rect 106 48599 152 48611
rect 106 47623 112 48599
rect 146 47623 152 48599
rect 106 47611 152 47623
rect -96 47573 96 47579
rect -96 47539 -84 47573
rect 84 47539 96 47573
rect -96 47533 96 47539
rect -96 47465 96 47471
rect -96 47431 -84 47465
rect 84 47431 96 47465
rect -96 47425 96 47431
rect -152 47381 -106 47393
rect -152 46405 -146 47381
rect -112 46405 -106 47381
rect -152 46393 -106 46405
rect 106 47381 152 47393
rect 106 46405 112 47381
rect 146 46405 152 47381
rect 106 46393 152 46405
rect -96 46355 96 46361
rect -96 46321 -84 46355
rect 84 46321 96 46355
rect -96 46315 96 46321
rect -96 46247 96 46253
rect -96 46213 -84 46247
rect 84 46213 96 46247
rect -96 46207 96 46213
rect -152 46163 -106 46175
rect -152 45187 -146 46163
rect -112 45187 -106 46163
rect -152 45175 -106 45187
rect 106 46163 152 46175
rect 106 45187 112 46163
rect 146 45187 152 46163
rect 106 45175 152 45187
rect -96 45137 96 45143
rect -96 45103 -84 45137
rect 84 45103 96 45137
rect -96 45097 96 45103
rect -96 45029 96 45035
rect -96 44995 -84 45029
rect 84 44995 96 45029
rect -96 44989 96 44995
rect -152 44945 -106 44957
rect -152 43969 -146 44945
rect -112 43969 -106 44945
rect -152 43957 -106 43969
rect 106 44945 152 44957
rect 106 43969 112 44945
rect 146 43969 152 44945
rect 106 43957 152 43969
rect -96 43919 96 43925
rect -96 43885 -84 43919
rect 84 43885 96 43919
rect -96 43879 96 43885
rect -96 43811 96 43817
rect -96 43777 -84 43811
rect 84 43777 96 43811
rect -96 43771 96 43777
rect -152 43727 -106 43739
rect -152 42751 -146 43727
rect -112 42751 -106 43727
rect -152 42739 -106 42751
rect 106 43727 152 43739
rect 106 42751 112 43727
rect 146 42751 152 43727
rect 106 42739 152 42751
rect -96 42701 96 42707
rect -96 42667 -84 42701
rect 84 42667 96 42701
rect -96 42661 96 42667
rect -96 42593 96 42599
rect -96 42559 -84 42593
rect 84 42559 96 42593
rect -96 42553 96 42559
rect -152 42509 -106 42521
rect -152 41533 -146 42509
rect -112 41533 -106 42509
rect -152 41521 -106 41533
rect 106 42509 152 42521
rect 106 41533 112 42509
rect 146 41533 152 42509
rect 106 41521 152 41533
rect -96 41483 96 41489
rect -96 41449 -84 41483
rect 84 41449 96 41483
rect -96 41443 96 41449
rect -96 41375 96 41381
rect -96 41341 -84 41375
rect 84 41341 96 41375
rect -96 41335 96 41341
rect -152 41291 -106 41303
rect -152 40315 -146 41291
rect -112 40315 -106 41291
rect -152 40303 -106 40315
rect 106 41291 152 41303
rect 106 40315 112 41291
rect 146 40315 152 41291
rect 106 40303 152 40315
rect -96 40265 96 40271
rect -96 40231 -84 40265
rect 84 40231 96 40265
rect -96 40225 96 40231
rect -96 40157 96 40163
rect -96 40123 -84 40157
rect 84 40123 96 40157
rect -96 40117 96 40123
rect -152 40073 -106 40085
rect -152 39097 -146 40073
rect -112 39097 -106 40073
rect -152 39085 -106 39097
rect 106 40073 152 40085
rect 106 39097 112 40073
rect 146 39097 152 40073
rect 106 39085 152 39097
rect -96 39047 96 39053
rect -96 39013 -84 39047
rect 84 39013 96 39047
rect -96 39007 96 39013
rect -96 38939 96 38945
rect -96 38905 -84 38939
rect 84 38905 96 38939
rect -96 38899 96 38905
rect -152 38855 -106 38867
rect -152 37879 -146 38855
rect -112 37879 -106 38855
rect -152 37867 -106 37879
rect 106 38855 152 38867
rect 106 37879 112 38855
rect 146 37879 152 38855
rect 106 37867 152 37879
rect -96 37829 96 37835
rect -96 37795 -84 37829
rect 84 37795 96 37829
rect -96 37789 96 37795
rect -96 37721 96 37727
rect -96 37687 -84 37721
rect 84 37687 96 37721
rect -96 37681 96 37687
rect -152 37637 -106 37649
rect -152 36661 -146 37637
rect -112 36661 -106 37637
rect -152 36649 -106 36661
rect 106 37637 152 37649
rect 106 36661 112 37637
rect 146 36661 152 37637
rect 106 36649 152 36661
rect -96 36611 96 36617
rect -96 36577 -84 36611
rect 84 36577 96 36611
rect -96 36571 96 36577
rect -96 36503 96 36509
rect -96 36469 -84 36503
rect 84 36469 96 36503
rect -96 36463 96 36469
rect -152 36419 -106 36431
rect -152 35443 -146 36419
rect -112 35443 -106 36419
rect -152 35431 -106 35443
rect 106 36419 152 36431
rect 106 35443 112 36419
rect 146 35443 152 36419
rect 106 35431 152 35443
rect -96 35393 96 35399
rect -96 35359 -84 35393
rect 84 35359 96 35393
rect -96 35353 96 35359
rect -96 35285 96 35291
rect -96 35251 -84 35285
rect 84 35251 96 35285
rect -96 35245 96 35251
rect -152 35201 -106 35213
rect -152 34225 -146 35201
rect -112 34225 -106 35201
rect -152 34213 -106 34225
rect 106 35201 152 35213
rect 106 34225 112 35201
rect 146 34225 152 35201
rect 106 34213 152 34225
rect -96 34175 96 34181
rect -96 34141 -84 34175
rect 84 34141 96 34175
rect -96 34135 96 34141
rect -96 34067 96 34073
rect -96 34033 -84 34067
rect 84 34033 96 34067
rect -96 34027 96 34033
rect -152 33983 -106 33995
rect -152 33007 -146 33983
rect -112 33007 -106 33983
rect -152 32995 -106 33007
rect 106 33983 152 33995
rect 106 33007 112 33983
rect 146 33007 152 33983
rect 106 32995 152 33007
rect -96 32957 96 32963
rect -96 32923 -84 32957
rect 84 32923 96 32957
rect -96 32917 96 32923
rect -96 32849 96 32855
rect -96 32815 -84 32849
rect 84 32815 96 32849
rect -96 32809 96 32815
rect -152 32765 -106 32777
rect -152 31789 -146 32765
rect -112 31789 -106 32765
rect -152 31777 -106 31789
rect 106 32765 152 32777
rect 106 31789 112 32765
rect 146 31789 152 32765
rect 106 31777 152 31789
rect -96 31739 96 31745
rect -96 31705 -84 31739
rect 84 31705 96 31739
rect -96 31699 96 31705
rect -96 31631 96 31637
rect -96 31597 -84 31631
rect 84 31597 96 31631
rect -96 31591 96 31597
rect -152 31547 -106 31559
rect -152 30571 -146 31547
rect -112 30571 -106 31547
rect -152 30559 -106 30571
rect 106 31547 152 31559
rect 106 30571 112 31547
rect 146 30571 152 31547
rect 106 30559 152 30571
rect -96 30521 96 30527
rect -96 30487 -84 30521
rect 84 30487 96 30521
rect -96 30481 96 30487
rect -96 30413 96 30419
rect -96 30379 -84 30413
rect 84 30379 96 30413
rect -96 30373 96 30379
rect -152 30329 -106 30341
rect -152 29353 -146 30329
rect -112 29353 -106 30329
rect -152 29341 -106 29353
rect 106 30329 152 30341
rect 106 29353 112 30329
rect 146 29353 152 30329
rect 106 29341 152 29353
rect -96 29303 96 29309
rect -96 29269 -84 29303
rect 84 29269 96 29303
rect -96 29263 96 29269
rect -96 29195 96 29201
rect -96 29161 -84 29195
rect 84 29161 96 29195
rect -96 29155 96 29161
rect -152 29111 -106 29123
rect -152 28135 -146 29111
rect -112 28135 -106 29111
rect -152 28123 -106 28135
rect 106 29111 152 29123
rect 106 28135 112 29111
rect 146 28135 152 29111
rect 106 28123 152 28135
rect -96 28085 96 28091
rect -96 28051 -84 28085
rect 84 28051 96 28085
rect -96 28045 96 28051
rect -96 27977 96 27983
rect -96 27943 -84 27977
rect 84 27943 96 27977
rect -96 27937 96 27943
rect -152 27893 -106 27905
rect -152 26917 -146 27893
rect -112 26917 -106 27893
rect -152 26905 -106 26917
rect 106 27893 152 27905
rect 106 26917 112 27893
rect 146 26917 152 27893
rect 106 26905 152 26917
rect -96 26867 96 26873
rect -96 26833 -84 26867
rect 84 26833 96 26867
rect -96 26827 96 26833
rect -96 26759 96 26765
rect -96 26725 -84 26759
rect 84 26725 96 26759
rect -96 26719 96 26725
rect -152 26675 -106 26687
rect -152 25699 -146 26675
rect -112 25699 -106 26675
rect -152 25687 -106 25699
rect 106 26675 152 26687
rect 106 25699 112 26675
rect 146 25699 152 26675
rect 106 25687 152 25699
rect -96 25649 96 25655
rect -96 25615 -84 25649
rect 84 25615 96 25649
rect -96 25609 96 25615
rect -96 25541 96 25547
rect -96 25507 -84 25541
rect 84 25507 96 25541
rect -96 25501 96 25507
rect -152 25457 -106 25469
rect -152 24481 -146 25457
rect -112 24481 -106 25457
rect -152 24469 -106 24481
rect 106 25457 152 25469
rect 106 24481 112 25457
rect 146 24481 152 25457
rect 106 24469 152 24481
rect -96 24431 96 24437
rect -96 24397 -84 24431
rect 84 24397 96 24431
rect -96 24391 96 24397
rect -96 24323 96 24329
rect -96 24289 -84 24323
rect 84 24289 96 24323
rect -96 24283 96 24289
rect -152 24239 -106 24251
rect -152 23263 -146 24239
rect -112 23263 -106 24239
rect -152 23251 -106 23263
rect 106 24239 152 24251
rect 106 23263 112 24239
rect 146 23263 152 24239
rect 106 23251 152 23263
rect -96 23213 96 23219
rect -96 23179 -84 23213
rect 84 23179 96 23213
rect -96 23173 96 23179
rect -96 23105 96 23111
rect -96 23071 -84 23105
rect 84 23071 96 23105
rect -96 23065 96 23071
rect -152 23021 -106 23033
rect -152 22045 -146 23021
rect -112 22045 -106 23021
rect -152 22033 -106 22045
rect 106 23021 152 23033
rect 106 22045 112 23021
rect 146 22045 152 23021
rect 106 22033 152 22045
rect -96 21995 96 22001
rect -96 21961 -84 21995
rect 84 21961 96 21995
rect -96 21955 96 21961
rect -96 21887 96 21893
rect -96 21853 -84 21887
rect 84 21853 96 21887
rect -96 21847 96 21853
rect -152 21803 -106 21815
rect -152 20827 -146 21803
rect -112 20827 -106 21803
rect -152 20815 -106 20827
rect 106 21803 152 21815
rect 106 20827 112 21803
rect 146 20827 152 21803
rect 106 20815 152 20827
rect -96 20777 96 20783
rect -96 20743 -84 20777
rect 84 20743 96 20777
rect -96 20737 96 20743
rect -96 20669 96 20675
rect -96 20635 -84 20669
rect 84 20635 96 20669
rect -96 20629 96 20635
rect -152 20585 -106 20597
rect -152 19609 -146 20585
rect -112 19609 -106 20585
rect -152 19597 -106 19609
rect 106 20585 152 20597
rect 106 19609 112 20585
rect 146 19609 152 20585
rect 106 19597 152 19609
rect -96 19559 96 19565
rect -96 19525 -84 19559
rect 84 19525 96 19559
rect -96 19519 96 19525
rect -96 19451 96 19457
rect -96 19417 -84 19451
rect 84 19417 96 19451
rect -96 19411 96 19417
rect -152 19367 -106 19379
rect -152 18391 -146 19367
rect -112 18391 -106 19367
rect -152 18379 -106 18391
rect 106 19367 152 19379
rect 106 18391 112 19367
rect 146 18391 152 19367
rect 106 18379 152 18391
rect -96 18341 96 18347
rect -96 18307 -84 18341
rect 84 18307 96 18341
rect -96 18301 96 18307
rect -96 18233 96 18239
rect -96 18199 -84 18233
rect 84 18199 96 18233
rect -96 18193 96 18199
rect -152 18149 -106 18161
rect -152 17173 -146 18149
rect -112 17173 -106 18149
rect -152 17161 -106 17173
rect 106 18149 152 18161
rect 106 17173 112 18149
rect 146 17173 152 18149
rect 106 17161 152 17173
rect -96 17123 96 17129
rect -96 17089 -84 17123
rect 84 17089 96 17123
rect -96 17083 96 17089
rect -96 17015 96 17021
rect -96 16981 -84 17015
rect 84 16981 96 17015
rect -96 16975 96 16981
rect -152 16931 -106 16943
rect -152 15955 -146 16931
rect -112 15955 -106 16931
rect -152 15943 -106 15955
rect 106 16931 152 16943
rect 106 15955 112 16931
rect 146 15955 152 16931
rect 106 15943 152 15955
rect -96 15905 96 15911
rect -96 15871 -84 15905
rect 84 15871 96 15905
rect -96 15865 96 15871
rect -96 15797 96 15803
rect -96 15763 -84 15797
rect 84 15763 96 15797
rect -96 15757 96 15763
rect -152 15713 -106 15725
rect -152 14737 -146 15713
rect -112 14737 -106 15713
rect -152 14725 -106 14737
rect 106 15713 152 15725
rect 106 14737 112 15713
rect 146 14737 152 15713
rect 106 14725 152 14737
rect -96 14687 96 14693
rect -96 14653 -84 14687
rect 84 14653 96 14687
rect -96 14647 96 14653
rect -96 14579 96 14585
rect -96 14545 -84 14579
rect 84 14545 96 14579
rect -96 14539 96 14545
rect -152 14495 -106 14507
rect -152 13519 -146 14495
rect -112 13519 -106 14495
rect -152 13507 -106 13519
rect 106 14495 152 14507
rect 106 13519 112 14495
rect 146 13519 152 14495
rect 106 13507 152 13519
rect -96 13469 96 13475
rect -96 13435 -84 13469
rect 84 13435 96 13469
rect -96 13429 96 13435
rect -96 13361 96 13367
rect -96 13327 -84 13361
rect 84 13327 96 13361
rect -96 13321 96 13327
rect -152 13277 -106 13289
rect -152 12301 -146 13277
rect -112 12301 -106 13277
rect -152 12289 -106 12301
rect 106 13277 152 13289
rect 106 12301 112 13277
rect 146 12301 152 13277
rect 106 12289 152 12301
rect -96 12251 96 12257
rect -96 12217 -84 12251
rect 84 12217 96 12251
rect -96 12211 96 12217
rect -96 12143 96 12149
rect -96 12109 -84 12143
rect 84 12109 96 12143
rect -96 12103 96 12109
rect -152 12059 -106 12071
rect -152 11083 -146 12059
rect -112 11083 -106 12059
rect -152 11071 -106 11083
rect 106 12059 152 12071
rect 106 11083 112 12059
rect 146 11083 152 12059
rect 106 11071 152 11083
rect -96 11033 96 11039
rect -96 10999 -84 11033
rect 84 10999 96 11033
rect -96 10993 96 10999
rect -96 10925 96 10931
rect -96 10891 -84 10925
rect 84 10891 96 10925
rect -96 10885 96 10891
rect -152 10841 -106 10853
rect -152 9865 -146 10841
rect -112 9865 -106 10841
rect -152 9853 -106 9865
rect 106 10841 152 10853
rect 106 9865 112 10841
rect 146 9865 152 10841
rect 106 9853 152 9865
rect -96 9815 96 9821
rect -96 9781 -84 9815
rect 84 9781 96 9815
rect -96 9775 96 9781
rect -96 9707 96 9713
rect -96 9673 -84 9707
rect 84 9673 96 9707
rect -96 9667 96 9673
rect -152 9623 -106 9635
rect -152 8647 -146 9623
rect -112 8647 -106 9623
rect -152 8635 -106 8647
rect 106 9623 152 9635
rect 106 8647 112 9623
rect 146 8647 152 9623
rect 106 8635 152 8647
rect -96 8597 96 8603
rect -96 8563 -84 8597
rect 84 8563 96 8597
rect -96 8557 96 8563
rect -96 8489 96 8495
rect -96 8455 -84 8489
rect 84 8455 96 8489
rect -96 8449 96 8455
rect -152 8405 -106 8417
rect -152 7429 -146 8405
rect -112 7429 -106 8405
rect -152 7417 -106 7429
rect 106 8405 152 8417
rect 106 7429 112 8405
rect 146 7429 152 8405
rect 106 7417 152 7429
rect -96 7379 96 7385
rect -96 7345 -84 7379
rect 84 7345 96 7379
rect -96 7339 96 7345
rect -96 7271 96 7277
rect -96 7237 -84 7271
rect 84 7237 96 7271
rect -96 7231 96 7237
rect -152 7187 -106 7199
rect -152 6211 -146 7187
rect -112 6211 -106 7187
rect -152 6199 -106 6211
rect 106 7187 152 7199
rect 106 6211 112 7187
rect 146 6211 152 7187
rect 106 6199 152 6211
rect -96 6161 96 6167
rect -96 6127 -84 6161
rect 84 6127 96 6161
rect -96 6121 96 6127
rect -96 6053 96 6059
rect -96 6019 -84 6053
rect 84 6019 96 6053
rect -96 6013 96 6019
rect -152 5969 -106 5981
rect -152 4993 -146 5969
rect -112 4993 -106 5969
rect -152 4981 -106 4993
rect 106 5969 152 5981
rect 106 4993 112 5969
rect 146 4993 152 5969
rect 106 4981 152 4993
rect -96 4943 96 4949
rect -96 4909 -84 4943
rect 84 4909 96 4943
rect -96 4903 96 4909
rect -96 4835 96 4841
rect -96 4801 -84 4835
rect 84 4801 96 4835
rect -96 4795 96 4801
rect -152 4751 -106 4763
rect -152 3775 -146 4751
rect -112 3775 -106 4751
rect -152 3763 -106 3775
rect 106 4751 152 4763
rect 106 3775 112 4751
rect 146 3775 152 4751
rect 106 3763 152 3775
rect -96 3725 96 3731
rect -96 3691 -84 3725
rect 84 3691 96 3725
rect -96 3685 96 3691
rect -96 3617 96 3623
rect -96 3583 -84 3617
rect 84 3583 96 3617
rect -96 3577 96 3583
rect -152 3533 -106 3545
rect -152 2557 -146 3533
rect -112 2557 -106 3533
rect -152 2545 -106 2557
rect 106 3533 152 3545
rect 106 2557 112 3533
rect 146 2557 152 3533
rect 106 2545 152 2557
rect -96 2507 96 2513
rect -96 2473 -84 2507
rect 84 2473 96 2507
rect -96 2467 96 2473
rect -96 2399 96 2405
rect -96 2365 -84 2399
rect 84 2365 96 2399
rect -96 2359 96 2365
rect -152 2315 -106 2327
rect -152 1339 -146 2315
rect -112 1339 -106 2315
rect -152 1327 -106 1339
rect 106 2315 152 2327
rect 106 1339 112 2315
rect 146 1339 152 2315
rect 106 1327 152 1339
rect -96 1289 96 1295
rect -96 1255 -84 1289
rect 84 1255 96 1289
rect -96 1249 96 1255
rect -96 1181 96 1187
rect -96 1147 -84 1181
rect 84 1147 96 1181
rect -96 1141 96 1147
rect -152 1097 -106 1109
rect -152 121 -146 1097
rect -112 121 -106 1097
rect -152 109 -106 121
rect 106 1097 152 1109
rect 106 121 112 1097
rect 146 121 152 1097
rect 106 109 152 121
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -121 -106 -109
rect -152 -1097 -146 -121
rect -112 -1097 -106 -121
rect -152 -1109 -106 -1097
rect 106 -121 152 -109
rect 106 -1097 112 -121
rect 146 -1097 152 -121
rect 106 -1109 152 -1097
rect -96 -1147 96 -1141
rect -96 -1181 -84 -1147
rect 84 -1181 96 -1147
rect -96 -1187 96 -1181
rect -96 -1255 96 -1249
rect -96 -1289 -84 -1255
rect 84 -1289 96 -1255
rect -96 -1295 96 -1289
rect -152 -1339 -106 -1327
rect -152 -2315 -146 -1339
rect -112 -2315 -106 -1339
rect -152 -2327 -106 -2315
rect 106 -1339 152 -1327
rect 106 -2315 112 -1339
rect 146 -2315 152 -1339
rect 106 -2327 152 -2315
rect -96 -2365 96 -2359
rect -96 -2399 -84 -2365
rect 84 -2399 96 -2365
rect -96 -2405 96 -2399
rect -96 -2473 96 -2467
rect -96 -2507 -84 -2473
rect 84 -2507 96 -2473
rect -96 -2513 96 -2507
rect -152 -2557 -106 -2545
rect -152 -3533 -146 -2557
rect -112 -3533 -106 -2557
rect -152 -3545 -106 -3533
rect 106 -2557 152 -2545
rect 106 -3533 112 -2557
rect 146 -3533 152 -2557
rect 106 -3545 152 -3533
rect -96 -3583 96 -3577
rect -96 -3617 -84 -3583
rect 84 -3617 96 -3583
rect -96 -3623 96 -3617
rect -96 -3691 96 -3685
rect -96 -3725 -84 -3691
rect 84 -3725 96 -3691
rect -96 -3731 96 -3725
rect -152 -3775 -106 -3763
rect -152 -4751 -146 -3775
rect -112 -4751 -106 -3775
rect -152 -4763 -106 -4751
rect 106 -3775 152 -3763
rect 106 -4751 112 -3775
rect 146 -4751 152 -3775
rect 106 -4763 152 -4751
rect -96 -4801 96 -4795
rect -96 -4835 -84 -4801
rect 84 -4835 96 -4801
rect -96 -4841 96 -4835
rect -96 -4909 96 -4903
rect -96 -4943 -84 -4909
rect 84 -4943 96 -4909
rect -96 -4949 96 -4943
rect -152 -4993 -106 -4981
rect -152 -5969 -146 -4993
rect -112 -5969 -106 -4993
rect -152 -5981 -106 -5969
rect 106 -4993 152 -4981
rect 106 -5969 112 -4993
rect 146 -5969 152 -4993
rect 106 -5981 152 -5969
rect -96 -6019 96 -6013
rect -96 -6053 -84 -6019
rect 84 -6053 96 -6019
rect -96 -6059 96 -6053
rect -96 -6127 96 -6121
rect -96 -6161 -84 -6127
rect 84 -6161 96 -6127
rect -96 -6167 96 -6161
rect -152 -6211 -106 -6199
rect -152 -7187 -146 -6211
rect -112 -7187 -106 -6211
rect -152 -7199 -106 -7187
rect 106 -6211 152 -6199
rect 106 -7187 112 -6211
rect 146 -7187 152 -6211
rect 106 -7199 152 -7187
rect -96 -7237 96 -7231
rect -96 -7271 -84 -7237
rect 84 -7271 96 -7237
rect -96 -7277 96 -7271
rect -96 -7345 96 -7339
rect -96 -7379 -84 -7345
rect 84 -7379 96 -7345
rect -96 -7385 96 -7379
rect -152 -7429 -106 -7417
rect -152 -8405 -146 -7429
rect -112 -8405 -106 -7429
rect -152 -8417 -106 -8405
rect 106 -7429 152 -7417
rect 106 -8405 112 -7429
rect 146 -8405 152 -7429
rect 106 -8417 152 -8405
rect -96 -8455 96 -8449
rect -96 -8489 -84 -8455
rect 84 -8489 96 -8455
rect -96 -8495 96 -8489
rect -96 -8563 96 -8557
rect -96 -8597 -84 -8563
rect 84 -8597 96 -8563
rect -96 -8603 96 -8597
rect -152 -8647 -106 -8635
rect -152 -9623 -146 -8647
rect -112 -9623 -106 -8647
rect -152 -9635 -106 -9623
rect 106 -8647 152 -8635
rect 106 -9623 112 -8647
rect 146 -9623 152 -8647
rect 106 -9635 152 -9623
rect -96 -9673 96 -9667
rect -96 -9707 -84 -9673
rect 84 -9707 96 -9673
rect -96 -9713 96 -9707
rect -96 -9781 96 -9775
rect -96 -9815 -84 -9781
rect 84 -9815 96 -9781
rect -96 -9821 96 -9815
rect -152 -9865 -106 -9853
rect -152 -10841 -146 -9865
rect -112 -10841 -106 -9865
rect -152 -10853 -106 -10841
rect 106 -9865 152 -9853
rect 106 -10841 112 -9865
rect 146 -10841 152 -9865
rect 106 -10853 152 -10841
rect -96 -10891 96 -10885
rect -96 -10925 -84 -10891
rect 84 -10925 96 -10891
rect -96 -10931 96 -10925
rect -96 -10999 96 -10993
rect -96 -11033 -84 -10999
rect 84 -11033 96 -10999
rect -96 -11039 96 -11033
rect -152 -11083 -106 -11071
rect -152 -12059 -146 -11083
rect -112 -12059 -106 -11083
rect -152 -12071 -106 -12059
rect 106 -11083 152 -11071
rect 106 -12059 112 -11083
rect 146 -12059 152 -11083
rect 106 -12071 152 -12059
rect -96 -12109 96 -12103
rect -96 -12143 -84 -12109
rect 84 -12143 96 -12109
rect -96 -12149 96 -12143
rect -96 -12217 96 -12211
rect -96 -12251 -84 -12217
rect 84 -12251 96 -12217
rect -96 -12257 96 -12251
rect -152 -12301 -106 -12289
rect -152 -13277 -146 -12301
rect -112 -13277 -106 -12301
rect -152 -13289 -106 -13277
rect 106 -12301 152 -12289
rect 106 -13277 112 -12301
rect 146 -13277 152 -12301
rect 106 -13289 152 -13277
rect -96 -13327 96 -13321
rect -96 -13361 -84 -13327
rect 84 -13361 96 -13327
rect -96 -13367 96 -13361
rect -96 -13435 96 -13429
rect -96 -13469 -84 -13435
rect 84 -13469 96 -13435
rect -96 -13475 96 -13469
rect -152 -13519 -106 -13507
rect -152 -14495 -146 -13519
rect -112 -14495 -106 -13519
rect -152 -14507 -106 -14495
rect 106 -13519 152 -13507
rect 106 -14495 112 -13519
rect 146 -14495 152 -13519
rect 106 -14507 152 -14495
rect -96 -14545 96 -14539
rect -96 -14579 -84 -14545
rect 84 -14579 96 -14545
rect -96 -14585 96 -14579
rect -96 -14653 96 -14647
rect -96 -14687 -84 -14653
rect 84 -14687 96 -14653
rect -96 -14693 96 -14687
rect -152 -14737 -106 -14725
rect -152 -15713 -146 -14737
rect -112 -15713 -106 -14737
rect -152 -15725 -106 -15713
rect 106 -14737 152 -14725
rect 106 -15713 112 -14737
rect 146 -15713 152 -14737
rect 106 -15725 152 -15713
rect -96 -15763 96 -15757
rect -96 -15797 -84 -15763
rect 84 -15797 96 -15763
rect -96 -15803 96 -15797
rect -96 -15871 96 -15865
rect -96 -15905 -84 -15871
rect 84 -15905 96 -15871
rect -96 -15911 96 -15905
rect -152 -15955 -106 -15943
rect -152 -16931 -146 -15955
rect -112 -16931 -106 -15955
rect -152 -16943 -106 -16931
rect 106 -15955 152 -15943
rect 106 -16931 112 -15955
rect 146 -16931 152 -15955
rect 106 -16943 152 -16931
rect -96 -16981 96 -16975
rect -96 -17015 -84 -16981
rect 84 -17015 96 -16981
rect -96 -17021 96 -17015
rect -96 -17089 96 -17083
rect -96 -17123 -84 -17089
rect 84 -17123 96 -17089
rect -96 -17129 96 -17123
rect -152 -17173 -106 -17161
rect -152 -18149 -146 -17173
rect -112 -18149 -106 -17173
rect -152 -18161 -106 -18149
rect 106 -17173 152 -17161
rect 106 -18149 112 -17173
rect 146 -18149 152 -17173
rect 106 -18161 152 -18149
rect -96 -18199 96 -18193
rect -96 -18233 -84 -18199
rect 84 -18233 96 -18199
rect -96 -18239 96 -18233
rect -96 -18307 96 -18301
rect -96 -18341 -84 -18307
rect 84 -18341 96 -18307
rect -96 -18347 96 -18341
rect -152 -18391 -106 -18379
rect -152 -19367 -146 -18391
rect -112 -19367 -106 -18391
rect -152 -19379 -106 -19367
rect 106 -18391 152 -18379
rect 106 -19367 112 -18391
rect 146 -19367 152 -18391
rect 106 -19379 152 -19367
rect -96 -19417 96 -19411
rect -96 -19451 -84 -19417
rect 84 -19451 96 -19417
rect -96 -19457 96 -19451
rect -96 -19525 96 -19519
rect -96 -19559 -84 -19525
rect 84 -19559 96 -19525
rect -96 -19565 96 -19559
rect -152 -19609 -106 -19597
rect -152 -20585 -146 -19609
rect -112 -20585 -106 -19609
rect -152 -20597 -106 -20585
rect 106 -19609 152 -19597
rect 106 -20585 112 -19609
rect 146 -20585 152 -19609
rect 106 -20597 152 -20585
rect -96 -20635 96 -20629
rect -96 -20669 -84 -20635
rect 84 -20669 96 -20635
rect -96 -20675 96 -20669
rect -96 -20743 96 -20737
rect -96 -20777 -84 -20743
rect 84 -20777 96 -20743
rect -96 -20783 96 -20777
rect -152 -20827 -106 -20815
rect -152 -21803 -146 -20827
rect -112 -21803 -106 -20827
rect -152 -21815 -106 -21803
rect 106 -20827 152 -20815
rect 106 -21803 112 -20827
rect 146 -21803 152 -20827
rect 106 -21815 152 -21803
rect -96 -21853 96 -21847
rect -96 -21887 -84 -21853
rect 84 -21887 96 -21853
rect -96 -21893 96 -21887
rect -96 -21961 96 -21955
rect -96 -21995 -84 -21961
rect 84 -21995 96 -21961
rect -96 -22001 96 -21995
rect -152 -22045 -106 -22033
rect -152 -23021 -146 -22045
rect -112 -23021 -106 -22045
rect -152 -23033 -106 -23021
rect 106 -22045 152 -22033
rect 106 -23021 112 -22045
rect 146 -23021 152 -22045
rect 106 -23033 152 -23021
rect -96 -23071 96 -23065
rect -96 -23105 -84 -23071
rect 84 -23105 96 -23071
rect -96 -23111 96 -23105
rect -96 -23179 96 -23173
rect -96 -23213 -84 -23179
rect 84 -23213 96 -23179
rect -96 -23219 96 -23213
rect -152 -23263 -106 -23251
rect -152 -24239 -146 -23263
rect -112 -24239 -106 -23263
rect -152 -24251 -106 -24239
rect 106 -23263 152 -23251
rect 106 -24239 112 -23263
rect 146 -24239 152 -23263
rect 106 -24251 152 -24239
rect -96 -24289 96 -24283
rect -96 -24323 -84 -24289
rect 84 -24323 96 -24289
rect -96 -24329 96 -24323
rect -96 -24397 96 -24391
rect -96 -24431 -84 -24397
rect 84 -24431 96 -24397
rect -96 -24437 96 -24431
rect -152 -24481 -106 -24469
rect -152 -25457 -146 -24481
rect -112 -25457 -106 -24481
rect -152 -25469 -106 -25457
rect 106 -24481 152 -24469
rect 106 -25457 112 -24481
rect 146 -25457 152 -24481
rect 106 -25469 152 -25457
rect -96 -25507 96 -25501
rect -96 -25541 -84 -25507
rect 84 -25541 96 -25507
rect -96 -25547 96 -25541
rect -96 -25615 96 -25609
rect -96 -25649 -84 -25615
rect 84 -25649 96 -25615
rect -96 -25655 96 -25649
rect -152 -25699 -106 -25687
rect -152 -26675 -146 -25699
rect -112 -26675 -106 -25699
rect -152 -26687 -106 -26675
rect 106 -25699 152 -25687
rect 106 -26675 112 -25699
rect 146 -26675 152 -25699
rect 106 -26687 152 -26675
rect -96 -26725 96 -26719
rect -96 -26759 -84 -26725
rect 84 -26759 96 -26725
rect -96 -26765 96 -26759
rect -96 -26833 96 -26827
rect -96 -26867 -84 -26833
rect 84 -26867 96 -26833
rect -96 -26873 96 -26867
rect -152 -26917 -106 -26905
rect -152 -27893 -146 -26917
rect -112 -27893 -106 -26917
rect -152 -27905 -106 -27893
rect 106 -26917 152 -26905
rect 106 -27893 112 -26917
rect 146 -27893 152 -26917
rect 106 -27905 152 -27893
rect -96 -27943 96 -27937
rect -96 -27977 -84 -27943
rect 84 -27977 96 -27943
rect -96 -27983 96 -27977
rect -96 -28051 96 -28045
rect -96 -28085 -84 -28051
rect 84 -28085 96 -28051
rect -96 -28091 96 -28085
rect -152 -28135 -106 -28123
rect -152 -29111 -146 -28135
rect -112 -29111 -106 -28135
rect -152 -29123 -106 -29111
rect 106 -28135 152 -28123
rect 106 -29111 112 -28135
rect 146 -29111 152 -28135
rect 106 -29123 152 -29111
rect -96 -29161 96 -29155
rect -96 -29195 -84 -29161
rect 84 -29195 96 -29161
rect -96 -29201 96 -29195
rect -96 -29269 96 -29263
rect -96 -29303 -84 -29269
rect 84 -29303 96 -29269
rect -96 -29309 96 -29303
rect -152 -29353 -106 -29341
rect -152 -30329 -146 -29353
rect -112 -30329 -106 -29353
rect -152 -30341 -106 -30329
rect 106 -29353 152 -29341
rect 106 -30329 112 -29353
rect 146 -30329 152 -29353
rect 106 -30341 152 -30329
rect -96 -30379 96 -30373
rect -96 -30413 -84 -30379
rect 84 -30413 96 -30379
rect -96 -30419 96 -30413
rect -96 -30487 96 -30481
rect -96 -30521 -84 -30487
rect 84 -30521 96 -30487
rect -96 -30527 96 -30521
rect -152 -30571 -106 -30559
rect -152 -31547 -146 -30571
rect -112 -31547 -106 -30571
rect -152 -31559 -106 -31547
rect 106 -30571 152 -30559
rect 106 -31547 112 -30571
rect 146 -31547 152 -30571
rect 106 -31559 152 -31547
rect -96 -31597 96 -31591
rect -96 -31631 -84 -31597
rect 84 -31631 96 -31597
rect -96 -31637 96 -31631
rect -96 -31705 96 -31699
rect -96 -31739 -84 -31705
rect 84 -31739 96 -31705
rect -96 -31745 96 -31739
rect -152 -31789 -106 -31777
rect -152 -32765 -146 -31789
rect -112 -32765 -106 -31789
rect -152 -32777 -106 -32765
rect 106 -31789 152 -31777
rect 106 -32765 112 -31789
rect 146 -32765 152 -31789
rect 106 -32777 152 -32765
rect -96 -32815 96 -32809
rect -96 -32849 -84 -32815
rect 84 -32849 96 -32815
rect -96 -32855 96 -32849
rect -96 -32923 96 -32917
rect -96 -32957 -84 -32923
rect 84 -32957 96 -32923
rect -96 -32963 96 -32957
rect -152 -33007 -106 -32995
rect -152 -33983 -146 -33007
rect -112 -33983 -106 -33007
rect -152 -33995 -106 -33983
rect 106 -33007 152 -32995
rect 106 -33983 112 -33007
rect 146 -33983 152 -33007
rect 106 -33995 152 -33983
rect -96 -34033 96 -34027
rect -96 -34067 -84 -34033
rect 84 -34067 96 -34033
rect -96 -34073 96 -34067
rect -96 -34141 96 -34135
rect -96 -34175 -84 -34141
rect 84 -34175 96 -34141
rect -96 -34181 96 -34175
rect -152 -34225 -106 -34213
rect -152 -35201 -146 -34225
rect -112 -35201 -106 -34225
rect -152 -35213 -106 -35201
rect 106 -34225 152 -34213
rect 106 -35201 112 -34225
rect 146 -35201 152 -34225
rect 106 -35213 152 -35201
rect -96 -35251 96 -35245
rect -96 -35285 -84 -35251
rect 84 -35285 96 -35251
rect -96 -35291 96 -35285
rect -96 -35359 96 -35353
rect -96 -35393 -84 -35359
rect 84 -35393 96 -35359
rect -96 -35399 96 -35393
rect -152 -35443 -106 -35431
rect -152 -36419 -146 -35443
rect -112 -36419 -106 -35443
rect -152 -36431 -106 -36419
rect 106 -35443 152 -35431
rect 106 -36419 112 -35443
rect 146 -36419 152 -35443
rect 106 -36431 152 -36419
rect -96 -36469 96 -36463
rect -96 -36503 -84 -36469
rect 84 -36503 96 -36469
rect -96 -36509 96 -36503
rect -96 -36577 96 -36571
rect -96 -36611 -84 -36577
rect 84 -36611 96 -36577
rect -96 -36617 96 -36611
rect -152 -36661 -106 -36649
rect -152 -37637 -146 -36661
rect -112 -37637 -106 -36661
rect -152 -37649 -106 -37637
rect 106 -36661 152 -36649
rect 106 -37637 112 -36661
rect 146 -37637 152 -36661
rect 106 -37649 152 -37637
rect -96 -37687 96 -37681
rect -96 -37721 -84 -37687
rect 84 -37721 96 -37687
rect -96 -37727 96 -37721
rect -96 -37795 96 -37789
rect -96 -37829 -84 -37795
rect 84 -37829 96 -37795
rect -96 -37835 96 -37829
rect -152 -37879 -106 -37867
rect -152 -38855 -146 -37879
rect -112 -38855 -106 -37879
rect -152 -38867 -106 -38855
rect 106 -37879 152 -37867
rect 106 -38855 112 -37879
rect 146 -38855 152 -37879
rect 106 -38867 152 -38855
rect -96 -38905 96 -38899
rect -96 -38939 -84 -38905
rect 84 -38939 96 -38905
rect -96 -38945 96 -38939
rect -96 -39013 96 -39007
rect -96 -39047 -84 -39013
rect 84 -39047 96 -39013
rect -96 -39053 96 -39047
rect -152 -39097 -106 -39085
rect -152 -40073 -146 -39097
rect -112 -40073 -106 -39097
rect -152 -40085 -106 -40073
rect 106 -39097 152 -39085
rect 106 -40073 112 -39097
rect 146 -40073 152 -39097
rect 106 -40085 152 -40073
rect -96 -40123 96 -40117
rect -96 -40157 -84 -40123
rect 84 -40157 96 -40123
rect -96 -40163 96 -40157
rect -96 -40231 96 -40225
rect -96 -40265 -84 -40231
rect 84 -40265 96 -40231
rect -96 -40271 96 -40265
rect -152 -40315 -106 -40303
rect -152 -41291 -146 -40315
rect -112 -41291 -106 -40315
rect -152 -41303 -106 -41291
rect 106 -40315 152 -40303
rect 106 -41291 112 -40315
rect 146 -41291 152 -40315
rect 106 -41303 152 -41291
rect -96 -41341 96 -41335
rect -96 -41375 -84 -41341
rect 84 -41375 96 -41341
rect -96 -41381 96 -41375
rect -96 -41449 96 -41443
rect -96 -41483 -84 -41449
rect 84 -41483 96 -41449
rect -96 -41489 96 -41483
rect -152 -41533 -106 -41521
rect -152 -42509 -146 -41533
rect -112 -42509 -106 -41533
rect -152 -42521 -106 -42509
rect 106 -41533 152 -41521
rect 106 -42509 112 -41533
rect 146 -42509 152 -41533
rect 106 -42521 152 -42509
rect -96 -42559 96 -42553
rect -96 -42593 -84 -42559
rect 84 -42593 96 -42559
rect -96 -42599 96 -42593
rect -96 -42667 96 -42661
rect -96 -42701 -84 -42667
rect 84 -42701 96 -42667
rect -96 -42707 96 -42701
rect -152 -42751 -106 -42739
rect -152 -43727 -146 -42751
rect -112 -43727 -106 -42751
rect -152 -43739 -106 -43727
rect 106 -42751 152 -42739
rect 106 -43727 112 -42751
rect 146 -43727 152 -42751
rect 106 -43739 152 -43727
rect -96 -43777 96 -43771
rect -96 -43811 -84 -43777
rect 84 -43811 96 -43777
rect -96 -43817 96 -43811
rect -96 -43885 96 -43879
rect -96 -43919 -84 -43885
rect 84 -43919 96 -43885
rect -96 -43925 96 -43919
rect -152 -43969 -106 -43957
rect -152 -44945 -146 -43969
rect -112 -44945 -106 -43969
rect -152 -44957 -106 -44945
rect 106 -43969 152 -43957
rect 106 -44945 112 -43969
rect 146 -44945 152 -43969
rect 106 -44957 152 -44945
rect -96 -44995 96 -44989
rect -96 -45029 -84 -44995
rect 84 -45029 96 -44995
rect -96 -45035 96 -45029
rect -96 -45103 96 -45097
rect -96 -45137 -84 -45103
rect 84 -45137 96 -45103
rect -96 -45143 96 -45137
rect -152 -45187 -106 -45175
rect -152 -46163 -146 -45187
rect -112 -46163 -106 -45187
rect -152 -46175 -106 -46163
rect 106 -45187 152 -45175
rect 106 -46163 112 -45187
rect 146 -46163 152 -45187
rect 106 -46175 152 -46163
rect -96 -46213 96 -46207
rect -96 -46247 -84 -46213
rect 84 -46247 96 -46213
rect -96 -46253 96 -46247
rect -96 -46321 96 -46315
rect -96 -46355 -84 -46321
rect 84 -46355 96 -46321
rect -96 -46361 96 -46355
rect -152 -46405 -106 -46393
rect -152 -47381 -146 -46405
rect -112 -47381 -106 -46405
rect -152 -47393 -106 -47381
rect 106 -46405 152 -46393
rect 106 -47381 112 -46405
rect 146 -47381 152 -46405
rect 106 -47393 152 -47381
rect -96 -47431 96 -47425
rect -96 -47465 -84 -47431
rect 84 -47465 96 -47431
rect -96 -47471 96 -47465
rect -96 -47539 96 -47533
rect -96 -47573 -84 -47539
rect 84 -47573 96 -47539
rect -96 -47579 96 -47573
rect -152 -47623 -106 -47611
rect -152 -48599 -146 -47623
rect -112 -48599 -106 -47623
rect -152 -48611 -106 -48599
rect 106 -47623 152 -47611
rect 106 -48599 112 -47623
rect 146 -48599 152 -47623
rect 106 -48611 152 -48599
rect -96 -48649 96 -48643
rect -96 -48683 -84 -48649
rect 84 -48683 96 -48649
rect -96 -48689 96 -48683
rect -96 -48757 96 -48751
rect -96 -48791 -84 -48757
rect 84 -48791 96 -48757
rect -96 -48797 96 -48791
rect -152 -48841 -106 -48829
rect -152 -49817 -146 -48841
rect -112 -49817 -106 -48841
rect -152 -49829 -106 -49817
rect 106 -48841 152 -48829
rect 106 -49817 112 -48841
rect 146 -49817 152 -48841
rect 106 -49829 152 -49817
rect -96 -49867 96 -49861
rect -96 -49901 -84 -49867
rect 84 -49901 96 -49867
rect -96 -49907 96 -49901
rect -96 -49975 96 -49969
rect -96 -50009 -84 -49975
rect 84 -50009 96 -49975
rect -96 -50015 96 -50009
rect -152 -50059 -106 -50047
rect -152 -51035 -146 -50059
rect -112 -51035 -106 -50059
rect -152 -51047 -106 -51035
rect 106 -50059 152 -50047
rect 106 -51035 112 -50059
rect 146 -51035 152 -50059
rect 106 -51047 152 -51035
rect -96 -51085 96 -51079
rect -96 -51119 -84 -51085
rect 84 -51119 96 -51085
rect -96 -51125 96 -51119
rect -96 -51193 96 -51187
rect -96 -51227 -84 -51193
rect 84 -51227 96 -51193
rect -96 -51233 96 -51227
rect -152 -51277 -106 -51265
rect -152 -52253 -146 -51277
rect -112 -52253 -106 -51277
rect -152 -52265 -106 -52253
rect 106 -51277 152 -51265
rect 106 -52253 112 -51277
rect 146 -52253 152 -51277
rect 106 -52265 152 -52253
rect -96 -52303 96 -52297
rect -96 -52337 -84 -52303
rect 84 -52337 96 -52303
rect -96 -52343 96 -52337
rect -96 -52411 96 -52405
rect -96 -52445 -84 -52411
rect 84 -52445 96 -52411
rect -96 -52451 96 -52445
rect -152 -52495 -106 -52483
rect -152 -53471 -146 -52495
rect -112 -53471 -106 -52495
rect -152 -53483 -106 -53471
rect 106 -52495 152 -52483
rect 106 -53471 112 -52495
rect 146 -53471 152 -52495
rect 106 -53483 152 -53471
rect -96 -53521 96 -53515
rect -96 -53555 -84 -53521
rect 84 -53555 96 -53521
rect -96 -53561 96 -53555
rect -96 -53629 96 -53623
rect -96 -53663 -84 -53629
rect 84 -53663 96 -53629
rect -96 -53669 96 -53663
rect -152 -53713 -106 -53701
rect -152 -54689 -146 -53713
rect -112 -54689 -106 -53713
rect -152 -54701 -106 -54689
rect 106 -53713 152 -53701
rect 106 -54689 112 -53713
rect 146 -54689 152 -53713
rect 106 -54701 152 -54689
rect -96 -54739 96 -54733
rect -96 -54773 -84 -54739
rect 84 -54773 96 -54739
rect -96 -54779 96 -54773
rect -96 -54847 96 -54841
rect -96 -54881 -84 -54847
rect 84 -54881 96 -54847
rect -96 -54887 96 -54881
rect -152 -54931 -106 -54919
rect -152 -55907 -146 -54931
rect -112 -55907 -106 -54931
rect -152 -55919 -106 -55907
rect 106 -54931 152 -54919
rect 106 -55907 112 -54931
rect 146 -55907 152 -54931
rect 106 -55919 152 -55907
rect -96 -55957 96 -55951
rect -96 -55991 -84 -55957
rect 84 -55991 96 -55957
rect -96 -55997 96 -55991
rect -96 -56065 96 -56059
rect -96 -56099 -84 -56065
rect 84 -56099 96 -56065
rect -96 -56105 96 -56099
rect -152 -56149 -106 -56137
rect -152 -57125 -146 -56149
rect -112 -57125 -106 -56149
rect -152 -57137 -106 -57125
rect 106 -56149 152 -56137
rect 106 -57125 112 -56149
rect 146 -57125 152 -56149
rect 106 -57137 152 -57125
rect -96 -57175 96 -57169
rect -96 -57209 -84 -57175
rect 84 -57209 96 -57175
rect -96 -57215 96 -57209
rect -96 -57283 96 -57277
rect -96 -57317 -84 -57283
rect 84 -57317 96 -57283
rect -96 -57323 96 -57317
rect -152 -57367 -106 -57355
rect -152 -58343 -146 -57367
rect -112 -58343 -106 -57367
rect -152 -58355 -106 -58343
rect 106 -57367 152 -57355
rect 106 -58343 112 -57367
rect 146 -58343 152 -57367
rect 106 -58355 152 -58343
rect -96 -58393 96 -58387
rect -96 -58427 -84 -58393
rect 84 -58427 96 -58393
rect -96 -58433 96 -58427
rect -96 -58501 96 -58495
rect -96 -58535 -84 -58501
rect 84 -58535 96 -58501
rect -96 -58541 96 -58535
rect -152 -58585 -106 -58573
rect -152 -59561 -146 -58585
rect -112 -59561 -106 -58585
rect -152 -59573 -106 -59561
rect 106 -58585 152 -58573
rect 106 -59561 112 -58585
rect 146 -59561 152 -58585
rect 106 -59573 152 -59561
rect -96 -59611 96 -59605
rect -96 -59645 -84 -59611
rect 84 -59645 96 -59611
rect -96 -59651 96 -59645
rect -96 -59719 96 -59713
rect -96 -59753 -84 -59719
rect 84 -59753 96 -59719
rect -96 -59759 96 -59753
rect -152 -59803 -106 -59791
rect -152 -60779 -146 -59803
rect -112 -60779 -106 -59803
rect -152 -60791 -106 -60779
rect 106 -59803 152 -59791
rect 106 -60779 112 -59803
rect 146 -60779 152 -59803
rect 106 -60791 152 -60779
rect -96 -60829 96 -60823
rect -96 -60863 -84 -60829
rect 84 -60863 96 -60829
rect -96 -60869 96 -60863
rect -96 -60937 96 -60931
rect -96 -60971 -84 -60937
rect 84 -60971 96 -60937
rect -96 -60977 96 -60971
rect -152 -61021 -106 -61009
rect -152 -61997 -146 -61021
rect -112 -61997 -106 -61021
rect -152 -62009 -106 -61997
rect 106 -61021 152 -61009
rect 106 -61997 112 -61021
rect 146 -61997 152 -61021
rect 106 -62009 152 -61997
rect -96 -62047 96 -62041
rect -96 -62081 -84 -62047
rect 84 -62081 96 -62047
rect -96 -62087 96 -62081
rect -96 -62155 96 -62149
rect -96 -62189 -84 -62155
rect 84 -62189 96 -62155
rect -96 -62195 96 -62189
rect -152 -62239 -106 -62227
rect -152 -63215 -146 -62239
rect -112 -63215 -106 -62239
rect -152 -63227 -106 -63215
rect 106 -62239 152 -62227
rect 106 -63215 112 -62239
rect 146 -63215 152 -62239
rect 106 -63227 152 -63215
rect -96 -63265 96 -63259
rect -96 -63299 -84 -63265
rect 84 -63299 96 -63265
rect -96 -63305 96 -63299
rect -96 -63373 96 -63367
rect -96 -63407 -84 -63373
rect 84 -63407 96 -63373
rect -96 -63413 96 -63407
rect -152 -63457 -106 -63445
rect -152 -64433 -146 -63457
rect -112 -64433 -106 -63457
rect -152 -64445 -106 -64433
rect 106 -63457 152 -63445
rect 106 -64433 112 -63457
rect 146 -64433 152 -63457
rect 106 -64445 152 -64433
rect -96 -64483 96 -64477
rect -96 -64517 -84 -64483
rect 84 -64517 96 -64483
rect -96 -64523 96 -64517
rect -96 -64591 96 -64585
rect -96 -64625 -84 -64591
rect 84 -64625 96 -64591
rect -96 -64631 96 -64625
rect -152 -64675 -106 -64663
rect -152 -65651 -146 -64675
rect -112 -65651 -106 -64675
rect -152 -65663 -106 -65651
rect 106 -64675 152 -64663
rect 106 -65651 112 -64675
rect 146 -65651 152 -64675
rect 106 -65663 152 -65651
rect -96 -65701 96 -65695
rect -96 -65735 -84 -65701
rect 84 -65735 96 -65701
rect -96 -65741 96 -65735
rect -96 -65809 96 -65803
rect -96 -65843 -84 -65809
rect 84 -65843 96 -65809
rect -96 -65849 96 -65843
rect -152 -65893 -106 -65881
rect -152 -66869 -146 -65893
rect -112 -66869 -106 -65893
rect -152 -66881 -106 -66869
rect 106 -65893 152 -65881
rect 106 -66869 112 -65893
rect 146 -66869 152 -65893
rect 106 -66881 152 -66869
rect -96 -66919 96 -66913
rect -96 -66953 -84 -66919
rect 84 -66953 96 -66919
rect -96 -66959 96 -66953
rect -96 -67027 96 -67021
rect -96 -67061 -84 -67027
rect 84 -67061 96 -67027
rect -96 -67067 96 -67061
rect -152 -67111 -106 -67099
rect -152 -68087 -146 -67111
rect -112 -68087 -106 -67111
rect -152 -68099 -106 -68087
rect 106 -67111 152 -67099
rect 106 -68087 112 -67111
rect 146 -68087 152 -67111
rect 106 -68099 152 -68087
rect -96 -68137 96 -68131
rect -96 -68171 -84 -68137
rect 84 -68171 96 -68137
rect -96 -68177 96 -68171
rect -96 -68245 96 -68239
rect -96 -68279 -84 -68245
rect 84 -68279 96 -68245
rect -96 -68285 96 -68279
rect -152 -68329 -106 -68317
rect -152 -69305 -146 -68329
rect -112 -69305 -106 -68329
rect -152 -69317 -106 -69305
rect 106 -68329 152 -68317
rect 106 -69305 112 -68329
rect 146 -69305 152 -68329
rect 106 -69317 152 -69305
rect -96 -69355 96 -69349
rect -96 -69389 -84 -69355
rect 84 -69389 96 -69355
rect -96 -69395 96 -69389
rect -96 -69463 96 -69457
rect -96 -69497 -84 -69463
rect 84 -69497 96 -69463
rect -96 -69503 96 -69497
rect -152 -69547 -106 -69535
rect -152 -70523 -146 -69547
rect -112 -70523 -106 -69547
rect -152 -70535 -106 -70523
rect 106 -69547 152 -69535
rect 106 -70523 112 -69547
rect 146 -70523 152 -69547
rect 106 -70535 152 -70523
rect -96 -70573 96 -70567
rect -96 -70607 -84 -70573
rect 84 -70607 96 -70573
rect -96 -70613 96 -70607
rect -96 -70681 96 -70675
rect -96 -70715 -84 -70681
rect 84 -70715 96 -70681
rect -96 -70721 96 -70715
rect -152 -70765 -106 -70753
rect -152 -71741 -146 -70765
rect -112 -71741 -106 -70765
rect -152 -71753 -106 -71741
rect 106 -70765 152 -70753
rect 106 -71741 112 -70765
rect 146 -71741 152 -70765
rect 106 -71753 152 -71741
rect -96 -71791 96 -71785
rect -96 -71825 -84 -71791
rect 84 -71825 96 -71791
rect -96 -71831 96 -71825
rect -96 -71899 96 -71893
rect -96 -71933 -84 -71899
rect 84 -71933 96 -71899
rect -96 -71939 96 -71933
rect -152 -71983 -106 -71971
rect -152 -72959 -146 -71983
rect -112 -72959 -106 -71983
rect -152 -72971 -106 -72959
rect 106 -71983 152 -71971
rect 106 -72959 112 -71983
rect 146 -72959 152 -71983
rect 106 -72971 152 -72959
rect -96 -73009 96 -73003
rect -96 -73043 -84 -73009
rect 84 -73043 96 -73009
rect -96 -73049 96 -73043
rect -96 -73117 96 -73111
rect -96 -73151 -84 -73117
rect 84 -73151 96 -73117
rect -96 -73157 96 -73151
rect -152 -73201 -106 -73189
rect -152 -74177 -146 -73201
rect -112 -74177 -106 -73201
rect -152 -74189 -106 -74177
rect 106 -73201 152 -73189
rect 106 -74177 112 -73201
rect 146 -74177 152 -73201
rect 106 -74189 152 -74177
rect -96 -74227 96 -74221
rect -96 -74261 -84 -74227
rect 84 -74261 96 -74227
rect -96 -74267 96 -74261
rect -96 -74335 96 -74329
rect -96 -74369 -84 -74335
rect 84 -74369 96 -74335
rect -96 -74375 96 -74369
rect -152 -74419 -106 -74407
rect -152 -75395 -146 -74419
rect -112 -75395 -106 -74419
rect -152 -75407 -106 -75395
rect 106 -74419 152 -74407
rect 106 -75395 112 -74419
rect 146 -75395 152 -74419
rect 106 -75407 152 -75395
rect -96 -75445 96 -75439
rect -96 -75479 -84 -75445
rect 84 -75479 96 -75445
rect -96 -75485 96 -75479
rect -96 -75553 96 -75547
rect -96 -75587 -84 -75553
rect 84 -75587 96 -75553
rect -96 -75593 96 -75587
rect -152 -75637 -106 -75625
rect -152 -76613 -146 -75637
rect -112 -76613 -106 -75637
rect -152 -76625 -106 -76613
rect 106 -75637 152 -75625
rect 106 -76613 112 -75637
rect 146 -76613 152 -75637
rect 106 -76625 152 -76613
rect -96 -76663 96 -76657
rect -96 -76697 -84 -76663
rect 84 -76697 96 -76663
rect -96 -76703 96 -76697
rect -96 -76771 96 -76765
rect -96 -76805 -84 -76771
rect 84 -76805 96 -76771
rect -96 -76811 96 -76805
rect -152 -76855 -106 -76843
rect -152 -77831 -146 -76855
rect -112 -77831 -106 -76855
rect -152 -77843 -106 -77831
rect 106 -76855 152 -76843
rect 106 -77831 112 -76855
rect 146 -77831 152 -76855
rect 106 -77843 152 -77831
rect -96 -77881 96 -77875
rect -96 -77915 -84 -77881
rect 84 -77915 96 -77881
rect -96 -77921 96 -77915
rect -96 -77989 96 -77983
rect -96 -78023 -84 -77989
rect 84 -78023 96 -77989
rect -96 -78029 96 -78023
rect -152 -78073 -106 -78061
rect -152 -79049 -146 -78073
rect -112 -79049 -106 -78073
rect -152 -79061 -106 -79049
rect 106 -78073 152 -78061
rect 106 -79049 112 -78073
rect 146 -79049 152 -78073
rect 106 -79061 152 -79049
rect -96 -79099 96 -79093
rect -96 -79133 -84 -79099
rect 84 -79133 96 -79099
rect -96 -79139 96 -79133
rect -96 -79207 96 -79201
rect -96 -79241 -84 -79207
rect 84 -79241 96 -79207
rect -96 -79247 96 -79241
rect -152 -79291 -106 -79279
rect -152 -80267 -146 -79291
rect -112 -80267 -106 -79291
rect -152 -80279 -106 -80267
rect 106 -79291 152 -79279
rect 106 -80267 112 -79291
rect 146 -80267 152 -79291
rect 106 -80279 152 -80267
rect -96 -80317 96 -80311
rect -96 -80351 -84 -80317
rect 84 -80351 96 -80317
rect -96 -80357 96 -80351
rect -96 -80425 96 -80419
rect -96 -80459 -84 -80425
rect 84 -80459 96 -80425
rect -96 -80465 96 -80459
rect -152 -80509 -106 -80497
rect -152 -81485 -146 -80509
rect -112 -81485 -106 -80509
rect -152 -81497 -106 -81485
rect 106 -80509 152 -80497
rect 106 -81485 112 -80509
rect 146 -81485 152 -80509
rect 106 -81497 152 -81485
rect -96 -81535 96 -81529
rect -96 -81569 -84 -81535
rect 84 -81569 96 -81535
rect -96 -81575 96 -81569
rect -96 -81643 96 -81637
rect -96 -81677 -84 -81643
rect 84 -81677 96 -81643
rect -96 -81683 96 -81677
rect -152 -81727 -106 -81715
rect -152 -82703 -146 -81727
rect -112 -82703 -106 -81727
rect -152 -82715 -106 -82703
rect 106 -81727 152 -81715
rect 106 -82703 112 -81727
rect 146 -82703 152 -81727
rect 106 -82715 152 -82703
rect -96 -82753 96 -82747
rect -96 -82787 -84 -82753
rect 84 -82787 96 -82753
rect -96 -82793 96 -82787
rect -96 -82861 96 -82855
rect -96 -82895 -84 -82861
rect 84 -82895 96 -82861
rect -96 -82901 96 -82895
rect -152 -82945 -106 -82933
rect -152 -83921 -146 -82945
rect -112 -83921 -106 -82945
rect -152 -83933 -106 -83921
rect 106 -82945 152 -82933
rect 106 -83921 112 -82945
rect 146 -83921 152 -82945
rect 106 -83933 152 -83921
rect -96 -83971 96 -83965
rect -96 -84005 -84 -83971
rect 84 -84005 96 -83971
rect -96 -84011 96 -84005
rect -96 -84079 96 -84073
rect -96 -84113 -84 -84079
rect 84 -84113 96 -84079
rect -96 -84119 96 -84113
rect -152 -84163 -106 -84151
rect -152 -85139 -146 -84163
rect -112 -85139 -106 -84163
rect -152 -85151 -106 -85139
rect 106 -84163 152 -84151
rect 106 -85139 112 -84163
rect 146 -85139 152 -84163
rect 106 -85151 152 -85139
rect -96 -85189 96 -85183
rect -96 -85223 -84 -85189
rect 84 -85223 96 -85189
rect -96 -85229 96 -85223
rect -96 -85297 96 -85291
rect -96 -85331 -84 -85297
rect 84 -85331 96 -85297
rect -96 -85337 96 -85331
rect -152 -85381 -106 -85369
rect -152 -86357 -146 -85381
rect -112 -86357 -106 -85381
rect -152 -86369 -106 -86357
rect 106 -85381 152 -85369
rect 106 -86357 112 -85381
rect 146 -86357 152 -85381
rect 106 -86369 152 -86357
rect -96 -86407 96 -86401
rect -96 -86441 -84 -86407
rect 84 -86441 96 -86407
rect -96 -86447 96 -86441
rect -96 -86515 96 -86509
rect -96 -86549 -84 -86515
rect 84 -86549 96 -86515
rect -96 -86555 96 -86549
rect -152 -86599 -106 -86587
rect -152 -87575 -146 -86599
rect -112 -87575 -106 -86599
rect -152 -87587 -106 -87575
rect 106 -86599 152 -86587
rect 106 -87575 112 -86599
rect 146 -87575 152 -86599
rect 106 -87587 152 -87575
rect -96 -87625 96 -87619
rect -96 -87659 -84 -87625
rect 84 -87659 96 -87625
rect -96 -87665 96 -87659
rect -96 -87733 96 -87727
rect -96 -87767 -84 -87733
rect 84 -87767 96 -87733
rect -96 -87773 96 -87767
rect -152 -87817 -106 -87805
rect -152 -88793 -146 -87817
rect -112 -88793 -106 -87817
rect -152 -88805 -106 -88793
rect 106 -87817 152 -87805
rect 106 -88793 112 -87817
rect 146 -88793 152 -87817
rect 106 -88805 152 -88793
rect -96 -88843 96 -88837
rect -96 -88877 -84 -88843
rect 84 -88877 96 -88843
rect -96 -88883 96 -88877
rect -96 -88951 96 -88945
rect -96 -88985 -84 -88951
rect 84 -88985 96 -88951
rect -96 -88991 96 -88985
rect -152 -89035 -106 -89023
rect -152 -90011 -146 -89035
rect -112 -90011 -106 -89035
rect -152 -90023 -106 -90011
rect 106 -89035 152 -89023
rect 106 -90011 112 -89035
rect 146 -90011 152 -89035
rect 106 -90023 152 -90011
rect -96 -90061 96 -90055
rect -96 -90095 -84 -90061
rect 84 -90095 96 -90061
rect -96 -90101 96 -90095
rect -96 -90169 96 -90163
rect -96 -90203 -84 -90169
rect 84 -90203 96 -90169
rect -96 -90209 96 -90203
rect -152 -90253 -106 -90241
rect -152 -91229 -146 -90253
rect -112 -91229 -106 -90253
rect -152 -91241 -106 -91229
rect 106 -90253 152 -90241
rect 106 -91229 112 -90253
rect 146 -91229 152 -90253
rect 106 -91241 152 -91229
rect -96 -91279 96 -91273
rect -96 -91313 -84 -91279
rect 84 -91313 96 -91279
rect -96 -91319 96 -91313
rect -96 -91387 96 -91381
rect -96 -91421 -84 -91387
rect 84 -91421 96 -91387
rect -96 -91427 96 -91421
rect -152 -91471 -106 -91459
rect -152 -92447 -146 -91471
rect -112 -92447 -106 -91471
rect -152 -92459 -106 -92447
rect 106 -91471 152 -91459
rect 106 -92447 112 -91471
rect 146 -92447 152 -91471
rect 106 -92459 152 -92447
rect -96 -92497 96 -92491
rect -96 -92531 -84 -92497
rect 84 -92531 96 -92497
rect -96 -92537 96 -92531
rect -96 -92605 96 -92599
rect -96 -92639 -84 -92605
rect 84 -92639 96 -92605
rect -96 -92645 96 -92639
rect -152 -92689 -106 -92677
rect -152 -93665 -146 -92689
rect -112 -93665 -106 -92689
rect -152 -93677 -106 -93665
rect 106 -92689 152 -92677
rect 106 -93665 112 -92689
rect 146 -93665 152 -92689
rect 106 -93677 152 -93665
rect -96 -93715 96 -93709
rect -96 -93749 -84 -93715
rect 84 -93749 96 -93715
rect -96 -93755 96 -93749
rect -96 -93823 96 -93817
rect -96 -93857 -84 -93823
rect 84 -93857 96 -93823
rect -96 -93863 96 -93857
rect -152 -93907 -106 -93895
rect -152 -94883 -146 -93907
rect -112 -94883 -106 -93907
rect -152 -94895 -106 -94883
rect 106 -93907 152 -93895
rect 106 -94883 112 -93907
rect 146 -94883 152 -93907
rect 106 -94895 152 -94883
rect -96 -94933 96 -94927
rect -96 -94967 -84 -94933
rect 84 -94967 96 -94933
rect -96 -94973 96 -94967
rect -96 -95041 96 -95035
rect -96 -95075 -84 -95041
rect 84 -95075 96 -95041
rect -96 -95081 96 -95075
rect -152 -95125 -106 -95113
rect -152 -96101 -146 -95125
rect -112 -96101 -106 -95125
rect -152 -96113 -106 -96101
rect 106 -95125 152 -95113
rect 106 -96101 112 -95125
rect 146 -96101 152 -95125
rect 106 -96113 152 -96101
rect -96 -96151 96 -96145
rect -96 -96185 -84 -96151
rect 84 -96185 96 -96151
rect -96 -96191 96 -96185
rect -96 -96259 96 -96253
rect -96 -96293 -84 -96259
rect 84 -96293 96 -96259
rect -96 -96299 96 -96293
rect -152 -96343 -106 -96331
rect -152 -97319 -146 -96343
rect -112 -97319 -106 -96343
rect -152 -97331 -106 -97319
rect 106 -96343 152 -96331
rect 106 -97319 112 -96343
rect 146 -97319 152 -96343
rect 106 -97331 152 -97319
rect -96 -97369 96 -97363
rect -96 -97403 -84 -97369
rect 84 -97403 96 -97369
rect -96 -97409 96 -97403
rect -96 -97477 96 -97471
rect -96 -97511 -84 -97477
rect 84 -97511 96 -97477
rect -96 -97517 96 -97511
rect -152 -97561 -106 -97549
rect -152 -98537 -146 -97561
rect -112 -98537 -106 -97561
rect -152 -98549 -106 -98537
rect 106 -97561 152 -97549
rect 106 -98537 112 -97561
rect 146 -98537 152 -97561
rect 106 -98549 152 -98537
rect -96 -98587 96 -98581
rect -96 -98621 -84 -98587
rect 84 -98621 96 -98587
rect -96 -98627 96 -98621
rect -96 -98695 96 -98689
rect -96 -98729 -84 -98695
rect 84 -98729 96 -98695
rect -96 -98735 96 -98729
rect -152 -98779 -106 -98767
rect -152 -99755 -146 -98779
rect -112 -99755 -106 -98779
rect -152 -99767 -106 -99755
rect 106 -98779 152 -98767
rect 106 -99755 112 -98779
rect 146 -99755 152 -98779
rect 106 -99767 152 -99755
rect -96 -99805 96 -99799
rect -96 -99839 -84 -99805
rect 84 -99839 96 -99805
rect -96 -99845 96 -99839
rect -96 -99913 96 -99907
rect -96 -99947 -84 -99913
rect 84 -99947 96 -99913
rect -96 -99953 96 -99947
rect -152 -99997 -106 -99985
rect -152 -100973 -146 -99997
rect -112 -100973 -106 -99997
rect -152 -100985 -106 -100973
rect 106 -99997 152 -99985
rect 106 -100973 112 -99997
rect 146 -100973 152 -99997
rect 106 -100985 152 -100973
rect -96 -101023 96 -101017
rect -96 -101057 -84 -101023
rect 84 -101057 96 -101023
rect -96 -101063 96 -101057
rect -96 -101131 96 -101125
rect -96 -101165 -84 -101131
rect 84 -101165 96 -101131
rect -96 -101171 96 -101165
rect -152 -101215 -106 -101203
rect -152 -102191 -146 -101215
rect -112 -102191 -106 -101215
rect -152 -102203 -106 -102191
rect 106 -101215 152 -101203
rect 106 -102191 112 -101215
rect 146 -102191 152 -101215
rect 106 -102203 152 -102191
rect -96 -102241 96 -102235
rect -96 -102275 -84 -102241
rect 84 -102275 96 -102241
rect -96 -102281 96 -102275
rect -96 -102349 96 -102343
rect -96 -102383 -84 -102349
rect 84 -102383 96 -102349
rect -96 -102389 96 -102383
rect -152 -102433 -106 -102421
rect -152 -103409 -146 -102433
rect -112 -103409 -106 -102433
rect -152 -103421 -106 -103409
rect 106 -102433 152 -102421
rect 106 -103409 112 -102433
rect 146 -103409 152 -102433
rect 106 -103421 152 -103409
rect -96 -103459 96 -103453
rect -96 -103493 -84 -103459
rect 84 -103493 96 -103459
rect -96 -103499 96 -103493
rect -96 -103567 96 -103561
rect -96 -103601 -84 -103567
rect 84 -103601 96 -103567
rect -96 -103607 96 -103601
rect -152 -103651 -106 -103639
rect -152 -104627 -146 -103651
rect -112 -104627 -106 -103651
rect -152 -104639 -106 -104627
rect 106 -103651 152 -103639
rect 106 -104627 112 -103651
rect 146 -104627 152 -103651
rect 106 -104639 152 -104627
rect -96 -104677 96 -104671
rect -96 -104711 -84 -104677
rect 84 -104711 96 -104677
rect -96 -104717 96 -104711
rect -96 -104785 96 -104779
rect -96 -104819 -84 -104785
rect 84 -104819 96 -104785
rect -96 -104825 96 -104819
rect -152 -104869 -106 -104857
rect -152 -105845 -146 -104869
rect -112 -105845 -106 -104869
rect -152 -105857 -106 -105845
rect 106 -104869 152 -104857
rect 106 -105845 112 -104869
rect 146 -105845 152 -104869
rect 106 -105857 152 -105845
rect -96 -105895 96 -105889
rect -96 -105929 -84 -105895
rect 84 -105929 96 -105895
rect -96 -105935 96 -105929
rect -96 -106003 96 -105997
rect -96 -106037 -84 -106003
rect 84 -106037 96 -106003
rect -96 -106043 96 -106037
rect -152 -106087 -106 -106075
rect -152 -107063 -146 -106087
rect -112 -107063 -106 -106087
rect -152 -107075 -106 -107063
rect 106 -106087 152 -106075
rect 106 -107063 112 -106087
rect 146 -107063 152 -106087
rect 106 -107075 152 -107063
rect -96 -107113 96 -107107
rect -96 -107147 -84 -107113
rect 84 -107147 96 -107113
rect -96 -107153 96 -107147
rect -96 -107221 96 -107215
rect -96 -107255 -84 -107221
rect 84 -107255 96 -107221
rect -96 -107261 96 -107255
rect -152 -107305 -106 -107293
rect -152 -108281 -146 -107305
rect -112 -108281 -106 -107305
rect -152 -108293 -106 -108281
rect 106 -107305 152 -107293
rect 106 -108281 112 -107305
rect 146 -108281 152 -107305
rect 106 -108293 152 -108281
rect -96 -108331 96 -108325
rect -96 -108365 -84 -108331
rect 84 -108365 96 -108331
rect -96 -108371 96 -108365
rect -96 -108439 96 -108433
rect -96 -108473 -84 -108439
rect 84 -108473 96 -108439
rect -96 -108479 96 -108473
rect -152 -108523 -106 -108511
rect -152 -109499 -146 -108523
rect -112 -109499 -106 -108523
rect -152 -109511 -106 -109499
rect 106 -108523 152 -108511
rect 106 -109499 112 -108523
rect 146 -109499 152 -108523
rect 106 -109511 152 -109499
rect -96 -109549 96 -109543
rect -96 -109583 -84 -109549
rect 84 -109583 96 -109549
rect -96 -109589 96 -109583
rect -96 -109657 96 -109651
rect -96 -109691 -84 -109657
rect 84 -109691 96 -109657
rect -96 -109697 96 -109691
rect -152 -109741 -106 -109729
rect -152 -110717 -146 -109741
rect -112 -110717 -106 -109741
rect -152 -110729 -106 -110717
rect 106 -109741 152 -109729
rect 106 -110717 112 -109741
rect 146 -110717 152 -109741
rect 106 -110729 152 -110717
rect -96 -110767 96 -110761
rect -96 -110801 -84 -110767
rect 84 -110801 96 -110767
rect -96 -110807 96 -110801
rect -96 -110875 96 -110869
rect -96 -110909 -84 -110875
rect 84 -110909 96 -110875
rect -96 -110915 96 -110909
rect -152 -110959 -106 -110947
rect -152 -111935 -146 -110959
rect -112 -111935 -106 -110959
rect -152 -111947 -106 -111935
rect 106 -110959 152 -110947
rect 106 -111935 112 -110959
rect 146 -111935 152 -110959
rect 106 -111947 152 -111935
rect -96 -111985 96 -111979
rect -96 -112019 -84 -111985
rect 84 -112019 96 -111985
rect -96 -112025 96 -112019
rect -96 -112093 96 -112087
rect -96 -112127 -84 -112093
rect 84 -112127 96 -112093
rect -96 -112133 96 -112127
rect -152 -112177 -106 -112165
rect -152 -113153 -146 -112177
rect -112 -113153 -106 -112177
rect -152 -113165 -106 -113153
rect 106 -112177 152 -112165
rect 106 -113153 112 -112177
rect 146 -113153 152 -112177
rect 106 -113165 152 -113153
rect -96 -113203 96 -113197
rect -96 -113237 -84 -113203
rect 84 -113237 96 -113203
rect -96 -113243 96 -113237
rect -96 -113311 96 -113305
rect -96 -113345 -84 -113311
rect 84 -113345 96 -113311
rect -96 -113351 96 -113345
rect -152 -113395 -106 -113383
rect -152 -114371 -146 -113395
rect -112 -114371 -106 -113395
rect -152 -114383 -106 -114371
rect 106 -113395 152 -113383
rect 106 -114371 112 -113395
rect 146 -114371 152 -113395
rect 106 -114383 152 -114371
rect -96 -114421 96 -114415
rect -96 -114455 -84 -114421
rect 84 -114455 96 -114421
rect -96 -114461 96 -114455
rect -96 -114529 96 -114523
rect -96 -114563 -84 -114529
rect 84 -114563 96 -114529
rect -96 -114569 96 -114563
rect -152 -114613 -106 -114601
rect -152 -115589 -146 -114613
rect -112 -115589 -106 -114613
rect -152 -115601 -106 -115589
rect 106 -114613 152 -114601
rect 106 -115589 112 -114613
rect 146 -115589 152 -114613
rect 106 -115601 152 -115589
rect -96 -115639 96 -115633
rect -96 -115673 -84 -115639
rect 84 -115673 96 -115639
rect -96 -115679 96 -115673
rect -96 -115747 96 -115741
rect -96 -115781 -84 -115747
rect 84 -115781 96 -115747
rect -96 -115787 96 -115781
rect -152 -115831 -106 -115819
rect -152 -116807 -146 -115831
rect -112 -116807 -106 -115831
rect -152 -116819 -106 -116807
rect 106 -115831 152 -115819
rect 106 -116807 112 -115831
rect 146 -116807 152 -115831
rect 106 -116819 152 -116807
rect -96 -116857 96 -116851
rect -96 -116891 -84 -116857
rect 84 -116891 96 -116857
rect -96 -116897 96 -116891
rect -96 -116965 96 -116959
rect -96 -116999 -84 -116965
rect 84 -116999 96 -116965
rect -96 -117005 96 -116999
rect -152 -117049 -106 -117037
rect -152 -118025 -146 -117049
rect -112 -118025 -106 -117049
rect -152 -118037 -106 -118025
rect 106 -117049 152 -117037
rect 106 -118025 112 -117049
rect 146 -118025 152 -117049
rect 106 -118037 152 -118025
rect -96 -118075 96 -118069
rect -96 -118109 -84 -118075
rect 84 -118109 96 -118075
rect -96 -118115 96 -118109
rect -96 -118183 96 -118177
rect -96 -118217 -84 -118183
rect 84 -118217 96 -118183
rect -96 -118223 96 -118217
rect -152 -118267 -106 -118255
rect -152 -119243 -146 -118267
rect -112 -119243 -106 -118267
rect -152 -119255 -106 -119243
rect 106 -118267 152 -118255
rect 106 -119243 112 -118267
rect 146 -119243 152 -118267
rect 106 -119255 152 -119243
rect -96 -119293 96 -119287
rect -96 -119327 -84 -119293
rect 84 -119327 96 -119293
rect -96 -119333 96 -119327
rect -96 -119401 96 -119395
rect -96 -119435 -84 -119401
rect 84 -119435 96 -119401
rect -96 -119441 96 -119435
rect -152 -119485 -106 -119473
rect -152 -120461 -146 -119485
rect -112 -120461 -106 -119485
rect -152 -120473 -106 -120461
rect 106 -119485 152 -119473
rect 106 -120461 112 -119485
rect 146 -120461 152 -119485
rect 106 -120473 152 -120461
rect -96 -120511 96 -120505
rect -96 -120545 -84 -120511
rect 84 -120545 96 -120511
rect -96 -120551 96 -120545
rect -96 -120619 96 -120613
rect -96 -120653 -84 -120619
rect 84 -120653 96 -120619
rect -96 -120659 96 -120653
rect -152 -120703 -106 -120691
rect -152 -121679 -146 -120703
rect -112 -121679 -106 -120703
rect -152 -121691 -106 -121679
rect 106 -120703 152 -120691
rect 106 -121679 112 -120703
rect 146 -121679 152 -120703
rect 106 -121691 152 -121679
rect -96 -121729 96 -121723
rect -96 -121763 -84 -121729
rect 84 -121763 96 -121729
rect -96 -121769 96 -121763
<< properties >>
string FIXED_BBOX -263 -121884 263 121884
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 1.0 m 200 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 ad {int((nf+1)/2) * W/nf * 0.29} as {int((nf+2)/2) * W/nf * 0.29} pd {2*int((nf+1)/2) * (W/nf + 0.29)} ps {2*int((nf+2)/2) * (W/nf + 0.29)} nrd {0.29 / W} nrs {0.29 / W} sa 0 sb 0 sd 0 mult 200
<< end >>
