magic
tech sky130A
magscale 1 2
timestamp 1730992408
<< pwell >>
rect -14394 -2070 14394 2070
<< psubdiff >>
rect -14358 2000 -14262 2034
rect 14262 2000 14358 2034
rect -14358 1938 -14324 2000
rect 14324 1938 14358 2000
rect -14358 -2000 -14324 -1938
rect 14324 -2000 14358 -1938
rect -14358 -2034 -14262 -2000
rect 14262 -2034 14358 -2000
<< psubdiffcont >>
rect -14262 2000 14262 2034
rect -14358 -1938 -14324 1938
rect 14324 -1938 14358 1938
rect -14262 -2034 14262 -2000
<< xpolycontact >>
rect -14228 1472 -14158 1904
rect -14228 -1904 -14158 -1472
rect -14062 1472 -13992 1904
rect -14062 -1904 -13992 -1472
rect -13896 1472 -13826 1904
rect -13896 -1904 -13826 -1472
rect -13730 1472 -13660 1904
rect -13730 -1904 -13660 -1472
rect -13564 1472 -13494 1904
rect -13564 -1904 -13494 -1472
rect -13398 1472 -13328 1904
rect -13398 -1904 -13328 -1472
rect -13232 1472 -13162 1904
rect -13232 -1904 -13162 -1472
rect -13066 1472 -12996 1904
rect -13066 -1904 -12996 -1472
rect -12900 1472 -12830 1904
rect -12900 -1904 -12830 -1472
rect -12734 1472 -12664 1904
rect -12734 -1904 -12664 -1472
rect -12568 1472 -12498 1904
rect -12568 -1904 -12498 -1472
rect -12402 1472 -12332 1904
rect -12402 -1904 -12332 -1472
rect -12236 1472 -12166 1904
rect -12236 -1904 -12166 -1472
rect -12070 1472 -12000 1904
rect -12070 -1904 -12000 -1472
rect -11904 1472 -11834 1904
rect -11904 -1904 -11834 -1472
rect -11738 1472 -11668 1904
rect -11738 -1904 -11668 -1472
rect -11572 1472 -11502 1904
rect -11572 -1904 -11502 -1472
rect -11406 1472 -11336 1904
rect -11406 -1904 -11336 -1472
rect -11240 1472 -11170 1904
rect -11240 -1904 -11170 -1472
rect -11074 1472 -11004 1904
rect -11074 -1904 -11004 -1472
rect -10908 1472 -10838 1904
rect -10908 -1904 -10838 -1472
rect -10742 1472 -10672 1904
rect -10742 -1904 -10672 -1472
rect -10576 1472 -10506 1904
rect -10576 -1904 -10506 -1472
rect -10410 1472 -10340 1904
rect -10410 -1904 -10340 -1472
rect -10244 1472 -10174 1904
rect -10244 -1904 -10174 -1472
rect -10078 1472 -10008 1904
rect -10078 -1904 -10008 -1472
rect -9912 1472 -9842 1904
rect -9912 -1904 -9842 -1472
rect -9746 1472 -9676 1904
rect -9746 -1904 -9676 -1472
rect -9580 1472 -9510 1904
rect -9580 -1904 -9510 -1472
rect -9414 1472 -9344 1904
rect -9414 -1904 -9344 -1472
rect -9248 1472 -9178 1904
rect -9248 -1904 -9178 -1472
rect -9082 1472 -9012 1904
rect -9082 -1904 -9012 -1472
rect -8916 1472 -8846 1904
rect -8916 -1904 -8846 -1472
rect -8750 1472 -8680 1904
rect -8750 -1904 -8680 -1472
rect -8584 1472 -8514 1904
rect -8584 -1904 -8514 -1472
rect -8418 1472 -8348 1904
rect -8418 -1904 -8348 -1472
rect -8252 1472 -8182 1904
rect -8252 -1904 -8182 -1472
rect -8086 1472 -8016 1904
rect -8086 -1904 -8016 -1472
rect -7920 1472 -7850 1904
rect -7920 -1904 -7850 -1472
rect -7754 1472 -7684 1904
rect -7754 -1904 -7684 -1472
rect -7588 1472 -7518 1904
rect -7588 -1904 -7518 -1472
rect -7422 1472 -7352 1904
rect -7422 -1904 -7352 -1472
rect -7256 1472 -7186 1904
rect -7256 -1904 -7186 -1472
rect -7090 1472 -7020 1904
rect -7090 -1904 -7020 -1472
rect -6924 1472 -6854 1904
rect -6924 -1904 -6854 -1472
rect -6758 1472 -6688 1904
rect -6758 -1904 -6688 -1472
rect -6592 1472 -6522 1904
rect -6592 -1904 -6522 -1472
rect -6426 1472 -6356 1904
rect -6426 -1904 -6356 -1472
rect -6260 1472 -6190 1904
rect -6260 -1904 -6190 -1472
rect -6094 1472 -6024 1904
rect -6094 -1904 -6024 -1472
rect -5928 1472 -5858 1904
rect -5928 -1904 -5858 -1472
rect -5762 1472 -5692 1904
rect -5762 -1904 -5692 -1472
rect -5596 1472 -5526 1904
rect -5596 -1904 -5526 -1472
rect -5430 1472 -5360 1904
rect -5430 -1904 -5360 -1472
rect -5264 1472 -5194 1904
rect -5264 -1904 -5194 -1472
rect -5098 1472 -5028 1904
rect -5098 -1904 -5028 -1472
rect -4932 1472 -4862 1904
rect -4932 -1904 -4862 -1472
rect -4766 1472 -4696 1904
rect -4766 -1904 -4696 -1472
rect -4600 1472 -4530 1904
rect -4600 -1904 -4530 -1472
rect -4434 1472 -4364 1904
rect -4434 -1904 -4364 -1472
rect -4268 1472 -4198 1904
rect -4268 -1904 -4198 -1472
rect -4102 1472 -4032 1904
rect -4102 -1904 -4032 -1472
rect -3936 1472 -3866 1904
rect -3936 -1904 -3866 -1472
rect -3770 1472 -3700 1904
rect -3770 -1904 -3700 -1472
rect -3604 1472 -3534 1904
rect -3604 -1904 -3534 -1472
rect -3438 1472 -3368 1904
rect -3438 -1904 -3368 -1472
rect -3272 1472 -3202 1904
rect -3272 -1904 -3202 -1472
rect -3106 1472 -3036 1904
rect -3106 -1904 -3036 -1472
rect -2940 1472 -2870 1904
rect -2940 -1904 -2870 -1472
rect -2774 1472 -2704 1904
rect -2774 -1904 -2704 -1472
rect -2608 1472 -2538 1904
rect -2608 -1904 -2538 -1472
rect -2442 1472 -2372 1904
rect -2442 -1904 -2372 -1472
rect -2276 1472 -2206 1904
rect -2276 -1904 -2206 -1472
rect -2110 1472 -2040 1904
rect -2110 -1904 -2040 -1472
rect -1944 1472 -1874 1904
rect -1944 -1904 -1874 -1472
rect -1778 1472 -1708 1904
rect -1778 -1904 -1708 -1472
rect -1612 1472 -1542 1904
rect -1612 -1904 -1542 -1472
rect -1446 1472 -1376 1904
rect -1446 -1904 -1376 -1472
rect -1280 1472 -1210 1904
rect -1280 -1904 -1210 -1472
rect -1114 1472 -1044 1904
rect -1114 -1904 -1044 -1472
rect -948 1472 -878 1904
rect -948 -1904 -878 -1472
rect -782 1472 -712 1904
rect -782 -1904 -712 -1472
rect -616 1472 -546 1904
rect -616 -1904 -546 -1472
rect -450 1472 -380 1904
rect -450 -1904 -380 -1472
rect -284 1472 -214 1904
rect -284 -1904 -214 -1472
rect -118 1472 -48 1904
rect -118 -1904 -48 -1472
rect 48 1472 118 1904
rect 48 -1904 118 -1472
rect 214 1472 284 1904
rect 214 -1904 284 -1472
rect 380 1472 450 1904
rect 380 -1904 450 -1472
rect 546 1472 616 1904
rect 546 -1904 616 -1472
rect 712 1472 782 1904
rect 712 -1904 782 -1472
rect 878 1472 948 1904
rect 878 -1904 948 -1472
rect 1044 1472 1114 1904
rect 1044 -1904 1114 -1472
rect 1210 1472 1280 1904
rect 1210 -1904 1280 -1472
rect 1376 1472 1446 1904
rect 1376 -1904 1446 -1472
rect 1542 1472 1612 1904
rect 1542 -1904 1612 -1472
rect 1708 1472 1778 1904
rect 1708 -1904 1778 -1472
rect 1874 1472 1944 1904
rect 1874 -1904 1944 -1472
rect 2040 1472 2110 1904
rect 2040 -1904 2110 -1472
rect 2206 1472 2276 1904
rect 2206 -1904 2276 -1472
rect 2372 1472 2442 1904
rect 2372 -1904 2442 -1472
rect 2538 1472 2608 1904
rect 2538 -1904 2608 -1472
rect 2704 1472 2774 1904
rect 2704 -1904 2774 -1472
rect 2870 1472 2940 1904
rect 2870 -1904 2940 -1472
rect 3036 1472 3106 1904
rect 3036 -1904 3106 -1472
rect 3202 1472 3272 1904
rect 3202 -1904 3272 -1472
rect 3368 1472 3438 1904
rect 3368 -1904 3438 -1472
rect 3534 1472 3604 1904
rect 3534 -1904 3604 -1472
rect 3700 1472 3770 1904
rect 3700 -1904 3770 -1472
rect 3866 1472 3936 1904
rect 3866 -1904 3936 -1472
rect 4032 1472 4102 1904
rect 4032 -1904 4102 -1472
rect 4198 1472 4268 1904
rect 4198 -1904 4268 -1472
rect 4364 1472 4434 1904
rect 4364 -1904 4434 -1472
rect 4530 1472 4600 1904
rect 4530 -1904 4600 -1472
rect 4696 1472 4766 1904
rect 4696 -1904 4766 -1472
rect 4862 1472 4932 1904
rect 4862 -1904 4932 -1472
rect 5028 1472 5098 1904
rect 5028 -1904 5098 -1472
rect 5194 1472 5264 1904
rect 5194 -1904 5264 -1472
rect 5360 1472 5430 1904
rect 5360 -1904 5430 -1472
rect 5526 1472 5596 1904
rect 5526 -1904 5596 -1472
rect 5692 1472 5762 1904
rect 5692 -1904 5762 -1472
rect 5858 1472 5928 1904
rect 5858 -1904 5928 -1472
rect 6024 1472 6094 1904
rect 6024 -1904 6094 -1472
rect 6190 1472 6260 1904
rect 6190 -1904 6260 -1472
rect 6356 1472 6426 1904
rect 6356 -1904 6426 -1472
rect 6522 1472 6592 1904
rect 6522 -1904 6592 -1472
rect 6688 1472 6758 1904
rect 6688 -1904 6758 -1472
rect 6854 1472 6924 1904
rect 6854 -1904 6924 -1472
rect 7020 1472 7090 1904
rect 7020 -1904 7090 -1472
rect 7186 1472 7256 1904
rect 7186 -1904 7256 -1472
rect 7352 1472 7422 1904
rect 7352 -1904 7422 -1472
rect 7518 1472 7588 1904
rect 7518 -1904 7588 -1472
rect 7684 1472 7754 1904
rect 7684 -1904 7754 -1472
rect 7850 1472 7920 1904
rect 7850 -1904 7920 -1472
rect 8016 1472 8086 1904
rect 8016 -1904 8086 -1472
rect 8182 1472 8252 1904
rect 8182 -1904 8252 -1472
rect 8348 1472 8418 1904
rect 8348 -1904 8418 -1472
rect 8514 1472 8584 1904
rect 8514 -1904 8584 -1472
rect 8680 1472 8750 1904
rect 8680 -1904 8750 -1472
rect 8846 1472 8916 1904
rect 8846 -1904 8916 -1472
rect 9012 1472 9082 1904
rect 9012 -1904 9082 -1472
rect 9178 1472 9248 1904
rect 9178 -1904 9248 -1472
rect 9344 1472 9414 1904
rect 9344 -1904 9414 -1472
rect 9510 1472 9580 1904
rect 9510 -1904 9580 -1472
rect 9676 1472 9746 1904
rect 9676 -1904 9746 -1472
rect 9842 1472 9912 1904
rect 9842 -1904 9912 -1472
rect 10008 1472 10078 1904
rect 10008 -1904 10078 -1472
rect 10174 1472 10244 1904
rect 10174 -1904 10244 -1472
rect 10340 1472 10410 1904
rect 10340 -1904 10410 -1472
rect 10506 1472 10576 1904
rect 10506 -1904 10576 -1472
rect 10672 1472 10742 1904
rect 10672 -1904 10742 -1472
rect 10838 1472 10908 1904
rect 10838 -1904 10908 -1472
rect 11004 1472 11074 1904
rect 11004 -1904 11074 -1472
rect 11170 1472 11240 1904
rect 11170 -1904 11240 -1472
rect 11336 1472 11406 1904
rect 11336 -1904 11406 -1472
rect 11502 1472 11572 1904
rect 11502 -1904 11572 -1472
rect 11668 1472 11738 1904
rect 11668 -1904 11738 -1472
rect 11834 1472 11904 1904
rect 11834 -1904 11904 -1472
rect 12000 1472 12070 1904
rect 12000 -1904 12070 -1472
rect 12166 1472 12236 1904
rect 12166 -1904 12236 -1472
rect 12332 1472 12402 1904
rect 12332 -1904 12402 -1472
rect 12498 1472 12568 1904
rect 12498 -1904 12568 -1472
rect 12664 1472 12734 1904
rect 12664 -1904 12734 -1472
rect 12830 1472 12900 1904
rect 12830 -1904 12900 -1472
rect 12996 1472 13066 1904
rect 12996 -1904 13066 -1472
rect 13162 1472 13232 1904
rect 13162 -1904 13232 -1472
rect 13328 1472 13398 1904
rect 13328 -1904 13398 -1472
rect 13494 1472 13564 1904
rect 13494 -1904 13564 -1472
rect 13660 1472 13730 1904
rect 13660 -1904 13730 -1472
rect 13826 1472 13896 1904
rect 13826 -1904 13896 -1472
rect 13992 1472 14062 1904
rect 13992 -1904 14062 -1472
rect 14158 1472 14228 1904
rect 14158 -1904 14228 -1472
<< xpolyres >>
rect -14228 -1472 -14158 1472
rect -14062 -1472 -13992 1472
rect -13896 -1472 -13826 1472
rect -13730 -1472 -13660 1472
rect -13564 -1472 -13494 1472
rect -13398 -1472 -13328 1472
rect -13232 -1472 -13162 1472
rect -13066 -1472 -12996 1472
rect -12900 -1472 -12830 1472
rect -12734 -1472 -12664 1472
rect -12568 -1472 -12498 1472
rect -12402 -1472 -12332 1472
rect -12236 -1472 -12166 1472
rect -12070 -1472 -12000 1472
rect -11904 -1472 -11834 1472
rect -11738 -1472 -11668 1472
rect -11572 -1472 -11502 1472
rect -11406 -1472 -11336 1472
rect -11240 -1472 -11170 1472
rect -11074 -1472 -11004 1472
rect -10908 -1472 -10838 1472
rect -10742 -1472 -10672 1472
rect -10576 -1472 -10506 1472
rect -10410 -1472 -10340 1472
rect -10244 -1472 -10174 1472
rect -10078 -1472 -10008 1472
rect -9912 -1472 -9842 1472
rect -9746 -1472 -9676 1472
rect -9580 -1472 -9510 1472
rect -9414 -1472 -9344 1472
rect -9248 -1472 -9178 1472
rect -9082 -1472 -9012 1472
rect -8916 -1472 -8846 1472
rect -8750 -1472 -8680 1472
rect -8584 -1472 -8514 1472
rect -8418 -1472 -8348 1472
rect -8252 -1472 -8182 1472
rect -8086 -1472 -8016 1472
rect -7920 -1472 -7850 1472
rect -7754 -1472 -7684 1472
rect -7588 -1472 -7518 1472
rect -7422 -1472 -7352 1472
rect -7256 -1472 -7186 1472
rect -7090 -1472 -7020 1472
rect -6924 -1472 -6854 1472
rect -6758 -1472 -6688 1472
rect -6592 -1472 -6522 1472
rect -6426 -1472 -6356 1472
rect -6260 -1472 -6190 1472
rect -6094 -1472 -6024 1472
rect -5928 -1472 -5858 1472
rect -5762 -1472 -5692 1472
rect -5596 -1472 -5526 1472
rect -5430 -1472 -5360 1472
rect -5264 -1472 -5194 1472
rect -5098 -1472 -5028 1472
rect -4932 -1472 -4862 1472
rect -4766 -1472 -4696 1472
rect -4600 -1472 -4530 1472
rect -4434 -1472 -4364 1472
rect -4268 -1472 -4198 1472
rect -4102 -1472 -4032 1472
rect -3936 -1472 -3866 1472
rect -3770 -1472 -3700 1472
rect -3604 -1472 -3534 1472
rect -3438 -1472 -3368 1472
rect -3272 -1472 -3202 1472
rect -3106 -1472 -3036 1472
rect -2940 -1472 -2870 1472
rect -2774 -1472 -2704 1472
rect -2608 -1472 -2538 1472
rect -2442 -1472 -2372 1472
rect -2276 -1472 -2206 1472
rect -2110 -1472 -2040 1472
rect -1944 -1472 -1874 1472
rect -1778 -1472 -1708 1472
rect -1612 -1472 -1542 1472
rect -1446 -1472 -1376 1472
rect -1280 -1472 -1210 1472
rect -1114 -1472 -1044 1472
rect -948 -1472 -878 1472
rect -782 -1472 -712 1472
rect -616 -1472 -546 1472
rect -450 -1472 -380 1472
rect -284 -1472 -214 1472
rect -118 -1472 -48 1472
rect 48 -1472 118 1472
rect 214 -1472 284 1472
rect 380 -1472 450 1472
rect 546 -1472 616 1472
rect 712 -1472 782 1472
rect 878 -1472 948 1472
rect 1044 -1472 1114 1472
rect 1210 -1472 1280 1472
rect 1376 -1472 1446 1472
rect 1542 -1472 1612 1472
rect 1708 -1472 1778 1472
rect 1874 -1472 1944 1472
rect 2040 -1472 2110 1472
rect 2206 -1472 2276 1472
rect 2372 -1472 2442 1472
rect 2538 -1472 2608 1472
rect 2704 -1472 2774 1472
rect 2870 -1472 2940 1472
rect 3036 -1472 3106 1472
rect 3202 -1472 3272 1472
rect 3368 -1472 3438 1472
rect 3534 -1472 3604 1472
rect 3700 -1472 3770 1472
rect 3866 -1472 3936 1472
rect 4032 -1472 4102 1472
rect 4198 -1472 4268 1472
rect 4364 -1472 4434 1472
rect 4530 -1472 4600 1472
rect 4696 -1472 4766 1472
rect 4862 -1472 4932 1472
rect 5028 -1472 5098 1472
rect 5194 -1472 5264 1472
rect 5360 -1472 5430 1472
rect 5526 -1472 5596 1472
rect 5692 -1472 5762 1472
rect 5858 -1472 5928 1472
rect 6024 -1472 6094 1472
rect 6190 -1472 6260 1472
rect 6356 -1472 6426 1472
rect 6522 -1472 6592 1472
rect 6688 -1472 6758 1472
rect 6854 -1472 6924 1472
rect 7020 -1472 7090 1472
rect 7186 -1472 7256 1472
rect 7352 -1472 7422 1472
rect 7518 -1472 7588 1472
rect 7684 -1472 7754 1472
rect 7850 -1472 7920 1472
rect 8016 -1472 8086 1472
rect 8182 -1472 8252 1472
rect 8348 -1472 8418 1472
rect 8514 -1472 8584 1472
rect 8680 -1472 8750 1472
rect 8846 -1472 8916 1472
rect 9012 -1472 9082 1472
rect 9178 -1472 9248 1472
rect 9344 -1472 9414 1472
rect 9510 -1472 9580 1472
rect 9676 -1472 9746 1472
rect 9842 -1472 9912 1472
rect 10008 -1472 10078 1472
rect 10174 -1472 10244 1472
rect 10340 -1472 10410 1472
rect 10506 -1472 10576 1472
rect 10672 -1472 10742 1472
rect 10838 -1472 10908 1472
rect 11004 -1472 11074 1472
rect 11170 -1472 11240 1472
rect 11336 -1472 11406 1472
rect 11502 -1472 11572 1472
rect 11668 -1472 11738 1472
rect 11834 -1472 11904 1472
rect 12000 -1472 12070 1472
rect 12166 -1472 12236 1472
rect 12332 -1472 12402 1472
rect 12498 -1472 12568 1472
rect 12664 -1472 12734 1472
rect 12830 -1472 12900 1472
rect 12996 -1472 13066 1472
rect 13162 -1472 13232 1472
rect 13328 -1472 13398 1472
rect 13494 -1472 13564 1472
rect 13660 -1472 13730 1472
rect 13826 -1472 13896 1472
rect 13992 -1472 14062 1472
rect 14158 -1472 14228 1472
<< locali >>
rect -14358 2000 -14262 2034
rect 14262 2000 14358 2034
rect -14358 1938 -14324 2000
rect 14324 1938 14358 2000
rect -14358 -2000 -14324 -1938
rect 14324 -2000 14358 -1938
rect -14358 -2034 -14262 -2000
rect 14262 -2034 14358 -2000
<< viali >>
rect -14212 1489 -14174 1886
rect -14046 1489 -14008 1886
rect -13880 1489 -13842 1886
rect -13714 1489 -13676 1886
rect -13548 1489 -13510 1886
rect -13382 1489 -13344 1886
rect -13216 1489 -13178 1886
rect -13050 1489 -13012 1886
rect -12884 1489 -12846 1886
rect -12718 1489 -12680 1886
rect -12552 1489 -12514 1886
rect -12386 1489 -12348 1886
rect -12220 1489 -12182 1886
rect -12054 1489 -12016 1886
rect -11888 1489 -11850 1886
rect -11722 1489 -11684 1886
rect -11556 1489 -11518 1886
rect -11390 1489 -11352 1886
rect -11224 1489 -11186 1886
rect -11058 1489 -11020 1886
rect -10892 1489 -10854 1886
rect -10726 1489 -10688 1886
rect -10560 1489 -10522 1886
rect -10394 1489 -10356 1886
rect -10228 1489 -10190 1886
rect -10062 1489 -10024 1886
rect -9896 1489 -9858 1886
rect -9730 1489 -9692 1886
rect -9564 1489 -9526 1886
rect -9398 1489 -9360 1886
rect -9232 1489 -9194 1886
rect -9066 1489 -9028 1886
rect -8900 1489 -8862 1886
rect -8734 1489 -8696 1886
rect -8568 1489 -8530 1886
rect -8402 1489 -8364 1886
rect -8236 1489 -8198 1886
rect -8070 1489 -8032 1886
rect -7904 1489 -7866 1886
rect -7738 1489 -7700 1886
rect -7572 1489 -7534 1886
rect -7406 1489 -7368 1886
rect -7240 1489 -7202 1886
rect -7074 1489 -7036 1886
rect -6908 1489 -6870 1886
rect -6742 1489 -6704 1886
rect -6576 1489 -6538 1886
rect -6410 1489 -6372 1886
rect -6244 1489 -6206 1886
rect -6078 1489 -6040 1886
rect -5912 1489 -5874 1886
rect -5746 1489 -5708 1886
rect -5580 1489 -5542 1886
rect -5414 1489 -5376 1886
rect -5248 1489 -5210 1886
rect -5082 1489 -5044 1886
rect -4916 1489 -4878 1886
rect -4750 1489 -4712 1886
rect -4584 1489 -4546 1886
rect -4418 1489 -4380 1886
rect -4252 1489 -4214 1886
rect -4086 1489 -4048 1886
rect -3920 1489 -3882 1886
rect -3754 1489 -3716 1886
rect -3588 1489 -3550 1886
rect -3422 1489 -3384 1886
rect -3256 1489 -3218 1886
rect -3090 1489 -3052 1886
rect -2924 1489 -2886 1886
rect -2758 1489 -2720 1886
rect -2592 1489 -2554 1886
rect -2426 1489 -2388 1886
rect -2260 1489 -2222 1886
rect -2094 1489 -2056 1886
rect -1928 1489 -1890 1886
rect -1762 1489 -1724 1886
rect -1596 1489 -1558 1886
rect -1430 1489 -1392 1886
rect -1264 1489 -1226 1886
rect -1098 1489 -1060 1886
rect -932 1489 -894 1886
rect -766 1489 -728 1886
rect -600 1489 -562 1886
rect -434 1489 -396 1886
rect -268 1489 -230 1886
rect -102 1489 -64 1886
rect 64 1489 102 1886
rect 230 1489 268 1886
rect 396 1489 434 1886
rect 562 1489 600 1886
rect 728 1489 766 1886
rect 894 1489 932 1886
rect 1060 1489 1098 1886
rect 1226 1489 1264 1886
rect 1392 1489 1430 1886
rect 1558 1489 1596 1886
rect 1724 1489 1762 1886
rect 1890 1489 1928 1886
rect 2056 1489 2094 1886
rect 2222 1489 2260 1886
rect 2388 1489 2426 1886
rect 2554 1489 2592 1886
rect 2720 1489 2758 1886
rect 2886 1489 2924 1886
rect 3052 1489 3090 1886
rect 3218 1489 3256 1886
rect 3384 1489 3422 1886
rect 3550 1489 3588 1886
rect 3716 1489 3754 1886
rect 3882 1489 3920 1886
rect 4048 1489 4086 1886
rect 4214 1489 4252 1886
rect 4380 1489 4418 1886
rect 4546 1489 4584 1886
rect 4712 1489 4750 1886
rect 4878 1489 4916 1886
rect 5044 1489 5082 1886
rect 5210 1489 5248 1886
rect 5376 1489 5414 1886
rect 5542 1489 5580 1886
rect 5708 1489 5746 1886
rect 5874 1489 5912 1886
rect 6040 1489 6078 1886
rect 6206 1489 6244 1886
rect 6372 1489 6410 1886
rect 6538 1489 6576 1886
rect 6704 1489 6742 1886
rect 6870 1489 6908 1886
rect 7036 1489 7074 1886
rect 7202 1489 7240 1886
rect 7368 1489 7406 1886
rect 7534 1489 7572 1886
rect 7700 1489 7738 1886
rect 7866 1489 7904 1886
rect 8032 1489 8070 1886
rect 8198 1489 8236 1886
rect 8364 1489 8402 1886
rect 8530 1489 8568 1886
rect 8696 1489 8734 1886
rect 8862 1489 8900 1886
rect 9028 1489 9066 1886
rect 9194 1489 9232 1886
rect 9360 1489 9398 1886
rect 9526 1489 9564 1886
rect 9692 1489 9730 1886
rect 9858 1489 9896 1886
rect 10024 1489 10062 1886
rect 10190 1489 10228 1886
rect 10356 1489 10394 1886
rect 10522 1489 10560 1886
rect 10688 1489 10726 1886
rect 10854 1489 10892 1886
rect 11020 1489 11058 1886
rect 11186 1489 11224 1886
rect 11352 1489 11390 1886
rect 11518 1489 11556 1886
rect 11684 1489 11722 1886
rect 11850 1489 11888 1886
rect 12016 1489 12054 1886
rect 12182 1489 12220 1886
rect 12348 1489 12386 1886
rect 12514 1489 12552 1886
rect 12680 1489 12718 1886
rect 12846 1489 12884 1886
rect 13012 1489 13050 1886
rect 13178 1489 13216 1886
rect 13344 1489 13382 1886
rect 13510 1489 13548 1886
rect 13676 1489 13714 1886
rect 13842 1489 13880 1886
rect 14008 1489 14046 1886
rect 14174 1489 14212 1886
rect -14212 -1886 -14174 -1489
rect -14046 -1886 -14008 -1489
rect -13880 -1886 -13842 -1489
rect -13714 -1886 -13676 -1489
rect -13548 -1886 -13510 -1489
rect -13382 -1886 -13344 -1489
rect -13216 -1886 -13178 -1489
rect -13050 -1886 -13012 -1489
rect -12884 -1886 -12846 -1489
rect -12718 -1886 -12680 -1489
rect -12552 -1886 -12514 -1489
rect -12386 -1886 -12348 -1489
rect -12220 -1886 -12182 -1489
rect -12054 -1886 -12016 -1489
rect -11888 -1886 -11850 -1489
rect -11722 -1886 -11684 -1489
rect -11556 -1886 -11518 -1489
rect -11390 -1886 -11352 -1489
rect -11224 -1886 -11186 -1489
rect -11058 -1886 -11020 -1489
rect -10892 -1886 -10854 -1489
rect -10726 -1886 -10688 -1489
rect -10560 -1886 -10522 -1489
rect -10394 -1886 -10356 -1489
rect -10228 -1886 -10190 -1489
rect -10062 -1886 -10024 -1489
rect -9896 -1886 -9858 -1489
rect -9730 -1886 -9692 -1489
rect -9564 -1886 -9526 -1489
rect -9398 -1886 -9360 -1489
rect -9232 -1886 -9194 -1489
rect -9066 -1886 -9028 -1489
rect -8900 -1886 -8862 -1489
rect -8734 -1886 -8696 -1489
rect -8568 -1886 -8530 -1489
rect -8402 -1886 -8364 -1489
rect -8236 -1886 -8198 -1489
rect -8070 -1886 -8032 -1489
rect -7904 -1886 -7866 -1489
rect -7738 -1886 -7700 -1489
rect -7572 -1886 -7534 -1489
rect -7406 -1886 -7368 -1489
rect -7240 -1886 -7202 -1489
rect -7074 -1886 -7036 -1489
rect -6908 -1886 -6870 -1489
rect -6742 -1886 -6704 -1489
rect -6576 -1886 -6538 -1489
rect -6410 -1886 -6372 -1489
rect -6244 -1886 -6206 -1489
rect -6078 -1886 -6040 -1489
rect -5912 -1886 -5874 -1489
rect -5746 -1886 -5708 -1489
rect -5580 -1886 -5542 -1489
rect -5414 -1886 -5376 -1489
rect -5248 -1886 -5210 -1489
rect -5082 -1886 -5044 -1489
rect -4916 -1886 -4878 -1489
rect -4750 -1886 -4712 -1489
rect -4584 -1886 -4546 -1489
rect -4418 -1886 -4380 -1489
rect -4252 -1886 -4214 -1489
rect -4086 -1886 -4048 -1489
rect -3920 -1886 -3882 -1489
rect -3754 -1886 -3716 -1489
rect -3588 -1886 -3550 -1489
rect -3422 -1886 -3384 -1489
rect -3256 -1886 -3218 -1489
rect -3090 -1886 -3052 -1489
rect -2924 -1886 -2886 -1489
rect -2758 -1886 -2720 -1489
rect -2592 -1886 -2554 -1489
rect -2426 -1886 -2388 -1489
rect -2260 -1886 -2222 -1489
rect -2094 -1886 -2056 -1489
rect -1928 -1886 -1890 -1489
rect -1762 -1886 -1724 -1489
rect -1596 -1886 -1558 -1489
rect -1430 -1886 -1392 -1489
rect -1264 -1886 -1226 -1489
rect -1098 -1886 -1060 -1489
rect -932 -1886 -894 -1489
rect -766 -1886 -728 -1489
rect -600 -1886 -562 -1489
rect -434 -1886 -396 -1489
rect -268 -1886 -230 -1489
rect -102 -1886 -64 -1489
rect 64 -1886 102 -1489
rect 230 -1886 268 -1489
rect 396 -1886 434 -1489
rect 562 -1886 600 -1489
rect 728 -1886 766 -1489
rect 894 -1886 932 -1489
rect 1060 -1886 1098 -1489
rect 1226 -1886 1264 -1489
rect 1392 -1886 1430 -1489
rect 1558 -1886 1596 -1489
rect 1724 -1886 1762 -1489
rect 1890 -1886 1928 -1489
rect 2056 -1886 2094 -1489
rect 2222 -1886 2260 -1489
rect 2388 -1886 2426 -1489
rect 2554 -1886 2592 -1489
rect 2720 -1886 2758 -1489
rect 2886 -1886 2924 -1489
rect 3052 -1886 3090 -1489
rect 3218 -1886 3256 -1489
rect 3384 -1886 3422 -1489
rect 3550 -1886 3588 -1489
rect 3716 -1886 3754 -1489
rect 3882 -1886 3920 -1489
rect 4048 -1886 4086 -1489
rect 4214 -1886 4252 -1489
rect 4380 -1886 4418 -1489
rect 4546 -1886 4584 -1489
rect 4712 -1886 4750 -1489
rect 4878 -1886 4916 -1489
rect 5044 -1886 5082 -1489
rect 5210 -1886 5248 -1489
rect 5376 -1886 5414 -1489
rect 5542 -1886 5580 -1489
rect 5708 -1886 5746 -1489
rect 5874 -1886 5912 -1489
rect 6040 -1886 6078 -1489
rect 6206 -1886 6244 -1489
rect 6372 -1886 6410 -1489
rect 6538 -1886 6576 -1489
rect 6704 -1886 6742 -1489
rect 6870 -1886 6908 -1489
rect 7036 -1886 7074 -1489
rect 7202 -1886 7240 -1489
rect 7368 -1886 7406 -1489
rect 7534 -1886 7572 -1489
rect 7700 -1886 7738 -1489
rect 7866 -1886 7904 -1489
rect 8032 -1886 8070 -1489
rect 8198 -1886 8236 -1489
rect 8364 -1886 8402 -1489
rect 8530 -1886 8568 -1489
rect 8696 -1886 8734 -1489
rect 8862 -1886 8900 -1489
rect 9028 -1886 9066 -1489
rect 9194 -1886 9232 -1489
rect 9360 -1886 9398 -1489
rect 9526 -1886 9564 -1489
rect 9692 -1886 9730 -1489
rect 9858 -1886 9896 -1489
rect 10024 -1886 10062 -1489
rect 10190 -1886 10228 -1489
rect 10356 -1886 10394 -1489
rect 10522 -1886 10560 -1489
rect 10688 -1886 10726 -1489
rect 10854 -1886 10892 -1489
rect 11020 -1886 11058 -1489
rect 11186 -1886 11224 -1489
rect 11352 -1886 11390 -1489
rect 11518 -1886 11556 -1489
rect 11684 -1886 11722 -1489
rect 11850 -1886 11888 -1489
rect 12016 -1886 12054 -1489
rect 12182 -1886 12220 -1489
rect 12348 -1886 12386 -1489
rect 12514 -1886 12552 -1489
rect 12680 -1886 12718 -1489
rect 12846 -1886 12884 -1489
rect 13012 -1886 13050 -1489
rect 13178 -1886 13216 -1489
rect 13344 -1886 13382 -1489
rect 13510 -1886 13548 -1489
rect 13676 -1886 13714 -1489
rect 13842 -1886 13880 -1489
rect 14008 -1886 14046 -1489
rect 14174 -1886 14212 -1489
<< metal1 >>
rect -14218 1886 -14168 1898
rect -14218 1489 -14212 1886
rect -14174 1489 -14168 1886
rect -14218 1477 -14168 1489
rect -14052 1886 -14002 1898
rect -14052 1489 -14046 1886
rect -14008 1489 -14002 1886
rect -14052 1477 -14002 1489
rect -13886 1886 -13836 1898
rect -13886 1489 -13880 1886
rect -13842 1489 -13836 1886
rect -13886 1477 -13836 1489
rect -13720 1886 -13670 1898
rect -13720 1489 -13714 1886
rect -13676 1489 -13670 1886
rect -13720 1477 -13670 1489
rect -13554 1886 -13504 1898
rect -13554 1489 -13548 1886
rect -13510 1489 -13504 1886
rect -13554 1477 -13504 1489
rect -13388 1886 -13338 1898
rect -13388 1489 -13382 1886
rect -13344 1489 -13338 1886
rect -13388 1477 -13338 1489
rect -13222 1886 -13172 1898
rect -13222 1489 -13216 1886
rect -13178 1489 -13172 1886
rect -13222 1477 -13172 1489
rect -13056 1886 -13006 1898
rect -13056 1489 -13050 1886
rect -13012 1489 -13006 1886
rect -13056 1477 -13006 1489
rect -12890 1886 -12840 1898
rect -12890 1489 -12884 1886
rect -12846 1489 -12840 1886
rect -12890 1477 -12840 1489
rect -12724 1886 -12674 1898
rect -12724 1489 -12718 1886
rect -12680 1489 -12674 1886
rect -12724 1477 -12674 1489
rect -12558 1886 -12508 1898
rect -12558 1489 -12552 1886
rect -12514 1489 -12508 1886
rect -12558 1477 -12508 1489
rect -12392 1886 -12342 1898
rect -12392 1489 -12386 1886
rect -12348 1489 -12342 1886
rect -12392 1477 -12342 1489
rect -12226 1886 -12176 1898
rect -12226 1489 -12220 1886
rect -12182 1489 -12176 1886
rect -12226 1477 -12176 1489
rect -12060 1886 -12010 1898
rect -12060 1489 -12054 1886
rect -12016 1489 -12010 1886
rect -12060 1477 -12010 1489
rect -11894 1886 -11844 1898
rect -11894 1489 -11888 1886
rect -11850 1489 -11844 1886
rect -11894 1477 -11844 1489
rect -11728 1886 -11678 1898
rect -11728 1489 -11722 1886
rect -11684 1489 -11678 1886
rect -11728 1477 -11678 1489
rect -11562 1886 -11512 1898
rect -11562 1489 -11556 1886
rect -11518 1489 -11512 1886
rect -11562 1477 -11512 1489
rect -11396 1886 -11346 1898
rect -11396 1489 -11390 1886
rect -11352 1489 -11346 1886
rect -11396 1477 -11346 1489
rect -11230 1886 -11180 1898
rect -11230 1489 -11224 1886
rect -11186 1489 -11180 1886
rect -11230 1477 -11180 1489
rect -11064 1886 -11014 1898
rect -11064 1489 -11058 1886
rect -11020 1489 -11014 1886
rect -11064 1477 -11014 1489
rect -10898 1886 -10848 1898
rect -10898 1489 -10892 1886
rect -10854 1489 -10848 1886
rect -10898 1477 -10848 1489
rect -10732 1886 -10682 1898
rect -10732 1489 -10726 1886
rect -10688 1489 -10682 1886
rect -10732 1477 -10682 1489
rect -10566 1886 -10516 1898
rect -10566 1489 -10560 1886
rect -10522 1489 -10516 1886
rect -10566 1477 -10516 1489
rect -10400 1886 -10350 1898
rect -10400 1489 -10394 1886
rect -10356 1489 -10350 1886
rect -10400 1477 -10350 1489
rect -10234 1886 -10184 1898
rect -10234 1489 -10228 1886
rect -10190 1489 -10184 1886
rect -10234 1477 -10184 1489
rect -10068 1886 -10018 1898
rect -10068 1489 -10062 1886
rect -10024 1489 -10018 1886
rect -10068 1477 -10018 1489
rect -9902 1886 -9852 1898
rect -9902 1489 -9896 1886
rect -9858 1489 -9852 1886
rect -9902 1477 -9852 1489
rect -9736 1886 -9686 1898
rect -9736 1489 -9730 1886
rect -9692 1489 -9686 1886
rect -9736 1477 -9686 1489
rect -9570 1886 -9520 1898
rect -9570 1489 -9564 1886
rect -9526 1489 -9520 1886
rect -9570 1477 -9520 1489
rect -9404 1886 -9354 1898
rect -9404 1489 -9398 1886
rect -9360 1489 -9354 1886
rect -9404 1477 -9354 1489
rect -9238 1886 -9188 1898
rect -9238 1489 -9232 1886
rect -9194 1489 -9188 1886
rect -9238 1477 -9188 1489
rect -9072 1886 -9022 1898
rect -9072 1489 -9066 1886
rect -9028 1489 -9022 1886
rect -9072 1477 -9022 1489
rect -8906 1886 -8856 1898
rect -8906 1489 -8900 1886
rect -8862 1489 -8856 1886
rect -8906 1477 -8856 1489
rect -8740 1886 -8690 1898
rect -8740 1489 -8734 1886
rect -8696 1489 -8690 1886
rect -8740 1477 -8690 1489
rect -8574 1886 -8524 1898
rect -8574 1489 -8568 1886
rect -8530 1489 -8524 1886
rect -8574 1477 -8524 1489
rect -8408 1886 -8358 1898
rect -8408 1489 -8402 1886
rect -8364 1489 -8358 1886
rect -8408 1477 -8358 1489
rect -8242 1886 -8192 1898
rect -8242 1489 -8236 1886
rect -8198 1489 -8192 1886
rect -8242 1477 -8192 1489
rect -8076 1886 -8026 1898
rect -8076 1489 -8070 1886
rect -8032 1489 -8026 1886
rect -8076 1477 -8026 1489
rect -7910 1886 -7860 1898
rect -7910 1489 -7904 1886
rect -7866 1489 -7860 1886
rect -7910 1477 -7860 1489
rect -7744 1886 -7694 1898
rect -7744 1489 -7738 1886
rect -7700 1489 -7694 1886
rect -7744 1477 -7694 1489
rect -7578 1886 -7528 1898
rect -7578 1489 -7572 1886
rect -7534 1489 -7528 1886
rect -7578 1477 -7528 1489
rect -7412 1886 -7362 1898
rect -7412 1489 -7406 1886
rect -7368 1489 -7362 1886
rect -7412 1477 -7362 1489
rect -7246 1886 -7196 1898
rect -7246 1489 -7240 1886
rect -7202 1489 -7196 1886
rect -7246 1477 -7196 1489
rect -7080 1886 -7030 1898
rect -7080 1489 -7074 1886
rect -7036 1489 -7030 1886
rect -7080 1477 -7030 1489
rect -6914 1886 -6864 1898
rect -6914 1489 -6908 1886
rect -6870 1489 -6864 1886
rect -6914 1477 -6864 1489
rect -6748 1886 -6698 1898
rect -6748 1489 -6742 1886
rect -6704 1489 -6698 1886
rect -6748 1477 -6698 1489
rect -6582 1886 -6532 1898
rect -6582 1489 -6576 1886
rect -6538 1489 -6532 1886
rect -6582 1477 -6532 1489
rect -6416 1886 -6366 1898
rect -6416 1489 -6410 1886
rect -6372 1489 -6366 1886
rect -6416 1477 -6366 1489
rect -6250 1886 -6200 1898
rect -6250 1489 -6244 1886
rect -6206 1489 -6200 1886
rect -6250 1477 -6200 1489
rect -6084 1886 -6034 1898
rect -6084 1489 -6078 1886
rect -6040 1489 -6034 1886
rect -6084 1477 -6034 1489
rect -5918 1886 -5868 1898
rect -5918 1489 -5912 1886
rect -5874 1489 -5868 1886
rect -5918 1477 -5868 1489
rect -5752 1886 -5702 1898
rect -5752 1489 -5746 1886
rect -5708 1489 -5702 1886
rect -5752 1477 -5702 1489
rect -5586 1886 -5536 1898
rect -5586 1489 -5580 1886
rect -5542 1489 -5536 1886
rect -5586 1477 -5536 1489
rect -5420 1886 -5370 1898
rect -5420 1489 -5414 1886
rect -5376 1489 -5370 1886
rect -5420 1477 -5370 1489
rect -5254 1886 -5204 1898
rect -5254 1489 -5248 1886
rect -5210 1489 -5204 1886
rect -5254 1477 -5204 1489
rect -5088 1886 -5038 1898
rect -5088 1489 -5082 1886
rect -5044 1489 -5038 1886
rect -5088 1477 -5038 1489
rect -4922 1886 -4872 1898
rect -4922 1489 -4916 1886
rect -4878 1489 -4872 1886
rect -4922 1477 -4872 1489
rect -4756 1886 -4706 1898
rect -4756 1489 -4750 1886
rect -4712 1489 -4706 1886
rect -4756 1477 -4706 1489
rect -4590 1886 -4540 1898
rect -4590 1489 -4584 1886
rect -4546 1489 -4540 1886
rect -4590 1477 -4540 1489
rect -4424 1886 -4374 1898
rect -4424 1489 -4418 1886
rect -4380 1489 -4374 1886
rect -4424 1477 -4374 1489
rect -4258 1886 -4208 1898
rect -4258 1489 -4252 1886
rect -4214 1489 -4208 1886
rect -4258 1477 -4208 1489
rect -4092 1886 -4042 1898
rect -4092 1489 -4086 1886
rect -4048 1489 -4042 1886
rect -4092 1477 -4042 1489
rect -3926 1886 -3876 1898
rect -3926 1489 -3920 1886
rect -3882 1489 -3876 1886
rect -3926 1477 -3876 1489
rect -3760 1886 -3710 1898
rect -3760 1489 -3754 1886
rect -3716 1489 -3710 1886
rect -3760 1477 -3710 1489
rect -3594 1886 -3544 1898
rect -3594 1489 -3588 1886
rect -3550 1489 -3544 1886
rect -3594 1477 -3544 1489
rect -3428 1886 -3378 1898
rect -3428 1489 -3422 1886
rect -3384 1489 -3378 1886
rect -3428 1477 -3378 1489
rect -3262 1886 -3212 1898
rect -3262 1489 -3256 1886
rect -3218 1489 -3212 1886
rect -3262 1477 -3212 1489
rect -3096 1886 -3046 1898
rect -3096 1489 -3090 1886
rect -3052 1489 -3046 1886
rect -3096 1477 -3046 1489
rect -2930 1886 -2880 1898
rect -2930 1489 -2924 1886
rect -2886 1489 -2880 1886
rect -2930 1477 -2880 1489
rect -2764 1886 -2714 1898
rect -2764 1489 -2758 1886
rect -2720 1489 -2714 1886
rect -2764 1477 -2714 1489
rect -2598 1886 -2548 1898
rect -2598 1489 -2592 1886
rect -2554 1489 -2548 1886
rect -2598 1477 -2548 1489
rect -2432 1886 -2382 1898
rect -2432 1489 -2426 1886
rect -2388 1489 -2382 1886
rect -2432 1477 -2382 1489
rect -2266 1886 -2216 1898
rect -2266 1489 -2260 1886
rect -2222 1489 -2216 1886
rect -2266 1477 -2216 1489
rect -2100 1886 -2050 1898
rect -2100 1489 -2094 1886
rect -2056 1489 -2050 1886
rect -2100 1477 -2050 1489
rect -1934 1886 -1884 1898
rect -1934 1489 -1928 1886
rect -1890 1489 -1884 1886
rect -1934 1477 -1884 1489
rect -1768 1886 -1718 1898
rect -1768 1489 -1762 1886
rect -1724 1489 -1718 1886
rect -1768 1477 -1718 1489
rect -1602 1886 -1552 1898
rect -1602 1489 -1596 1886
rect -1558 1489 -1552 1886
rect -1602 1477 -1552 1489
rect -1436 1886 -1386 1898
rect -1436 1489 -1430 1886
rect -1392 1489 -1386 1886
rect -1436 1477 -1386 1489
rect -1270 1886 -1220 1898
rect -1270 1489 -1264 1886
rect -1226 1489 -1220 1886
rect -1270 1477 -1220 1489
rect -1104 1886 -1054 1898
rect -1104 1489 -1098 1886
rect -1060 1489 -1054 1886
rect -1104 1477 -1054 1489
rect -938 1886 -888 1898
rect -938 1489 -932 1886
rect -894 1489 -888 1886
rect -938 1477 -888 1489
rect -772 1886 -722 1898
rect -772 1489 -766 1886
rect -728 1489 -722 1886
rect -772 1477 -722 1489
rect -606 1886 -556 1898
rect -606 1489 -600 1886
rect -562 1489 -556 1886
rect -606 1477 -556 1489
rect -440 1886 -390 1898
rect -440 1489 -434 1886
rect -396 1489 -390 1886
rect -440 1477 -390 1489
rect -274 1886 -224 1898
rect -274 1489 -268 1886
rect -230 1489 -224 1886
rect -274 1477 -224 1489
rect -108 1886 -58 1898
rect -108 1489 -102 1886
rect -64 1489 -58 1886
rect -108 1477 -58 1489
rect 58 1886 108 1898
rect 58 1489 64 1886
rect 102 1489 108 1886
rect 58 1477 108 1489
rect 224 1886 274 1898
rect 224 1489 230 1886
rect 268 1489 274 1886
rect 224 1477 274 1489
rect 390 1886 440 1898
rect 390 1489 396 1886
rect 434 1489 440 1886
rect 390 1477 440 1489
rect 556 1886 606 1898
rect 556 1489 562 1886
rect 600 1489 606 1886
rect 556 1477 606 1489
rect 722 1886 772 1898
rect 722 1489 728 1886
rect 766 1489 772 1886
rect 722 1477 772 1489
rect 888 1886 938 1898
rect 888 1489 894 1886
rect 932 1489 938 1886
rect 888 1477 938 1489
rect 1054 1886 1104 1898
rect 1054 1489 1060 1886
rect 1098 1489 1104 1886
rect 1054 1477 1104 1489
rect 1220 1886 1270 1898
rect 1220 1489 1226 1886
rect 1264 1489 1270 1886
rect 1220 1477 1270 1489
rect 1386 1886 1436 1898
rect 1386 1489 1392 1886
rect 1430 1489 1436 1886
rect 1386 1477 1436 1489
rect 1552 1886 1602 1898
rect 1552 1489 1558 1886
rect 1596 1489 1602 1886
rect 1552 1477 1602 1489
rect 1718 1886 1768 1898
rect 1718 1489 1724 1886
rect 1762 1489 1768 1886
rect 1718 1477 1768 1489
rect 1884 1886 1934 1898
rect 1884 1489 1890 1886
rect 1928 1489 1934 1886
rect 1884 1477 1934 1489
rect 2050 1886 2100 1898
rect 2050 1489 2056 1886
rect 2094 1489 2100 1886
rect 2050 1477 2100 1489
rect 2216 1886 2266 1898
rect 2216 1489 2222 1886
rect 2260 1489 2266 1886
rect 2216 1477 2266 1489
rect 2382 1886 2432 1898
rect 2382 1489 2388 1886
rect 2426 1489 2432 1886
rect 2382 1477 2432 1489
rect 2548 1886 2598 1898
rect 2548 1489 2554 1886
rect 2592 1489 2598 1886
rect 2548 1477 2598 1489
rect 2714 1886 2764 1898
rect 2714 1489 2720 1886
rect 2758 1489 2764 1886
rect 2714 1477 2764 1489
rect 2880 1886 2930 1898
rect 2880 1489 2886 1886
rect 2924 1489 2930 1886
rect 2880 1477 2930 1489
rect 3046 1886 3096 1898
rect 3046 1489 3052 1886
rect 3090 1489 3096 1886
rect 3046 1477 3096 1489
rect 3212 1886 3262 1898
rect 3212 1489 3218 1886
rect 3256 1489 3262 1886
rect 3212 1477 3262 1489
rect 3378 1886 3428 1898
rect 3378 1489 3384 1886
rect 3422 1489 3428 1886
rect 3378 1477 3428 1489
rect 3544 1886 3594 1898
rect 3544 1489 3550 1886
rect 3588 1489 3594 1886
rect 3544 1477 3594 1489
rect 3710 1886 3760 1898
rect 3710 1489 3716 1886
rect 3754 1489 3760 1886
rect 3710 1477 3760 1489
rect 3876 1886 3926 1898
rect 3876 1489 3882 1886
rect 3920 1489 3926 1886
rect 3876 1477 3926 1489
rect 4042 1886 4092 1898
rect 4042 1489 4048 1886
rect 4086 1489 4092 1886
rect 4042 1477 4092 1489
rect 4208 1886 4258 1898
rect 4208 1489 4214 1886
rect 4252 1489 4258 1886
rect 4208 1477 4258 1489
rect 4374 1886 4424 1898
rect 4374 1489 4380 1886
rect 4418 1489 4424 1886
rect 4374 1477 4424 1489
rect 4540 1886 4590 1898
rect 4540 1489 4546 1886
rect 4584 1489 4590 1886
rect 4540 1477 4590 1489
rect 4706 1886 4756 1898
rect 4706 1489 4712 1886
rect 4750 1489 4756 1886
rect 4706 1477 4756 1489
rect 4872 1886 4922 1898
rect 4872 1489 4878 1886
rect 4916 1489 4922 1886
rect 4872 1477 4922 1489
rect 5038 1886 5088 1898
rect 5038 1489 5044 1886
rect 5082 1489 5088 1886
rect 5038 1477 5088 1489
rect 5204 1886 5254 1898
rect 5204 1489 5210 1886
rect 5248 1489 5254 1886
rect 5204 1477 5254 1489
rect 5370 1886 5420 1898
rect 5370 1489 5376 1886
rect 5414 1489 5420 1886
rect 5370 1477 5420 1489
rect 5536 1886 5586 1898
rect 5536 1489 5542 1886
rect 5580 1489 5586 1886
rect 5536 1477 5586 1489
rect 5702 1886 5752 1898
rect 5702 1489 5708 1886
rect 5746 1489 5752 1886
rect 5702 1477 5752 1489
rect 5868 1886 5918 1898
rect 5868 1489 5874 1886
rect 5912 1489 5918 1886
rect 5868 1477 5918 1489
rect 6034 1886 6084 1898
rect 6034 1489 6040 1886
rect 6078 1489 6084 1886
rect 6034 1477 6084 1489
rect 6200 1886 6250 1898
rect 6200 1489 6206 1886
rect 6244 1489 6250 1886
rect 6200 1477 6250 1489
rect 6366 1886 6416 1898
rect 6366 1489 6372 1886
rect 6410 1489 6416 1886
rect 6366 1477 6416 1489
rect 6532 1886 6582 1898
rect 6532 1489 6538 1886
rect 6576 1489 6582 1886
rect 6532 1477 6582 1489
rect 6698 1886 6748 1898
rect 6698 1489 6704 1886
rect 6742 1489 6748 1886
rect 6698 1477 6748 1489
rect 6864 1886 6914 1898
rect 6864 1489 6870 1886
rect 6908 1489 6914 1886
rect 6864 1477 6914 1489
rect 7030 1886 7080 1898
rect 7030 1489 7036 1886
rect 7074 1489 7080 1886
rect 7030 1477 7080 1489
rect 7196 1886 7246 1898
rect 7196 1489 7202 1886
rect 7240 1489 7246 1886
rect 7196 1477 7246 1489
rect 7362 1886 7412 1898
rect 7362 1489 7368 1886
rect 7406 1489 7412 1886
rect 7362 1477 7412 1489
rect 7528 1886 7578 1898
rect 7528 1489 7534 1886
rect 7572 1489 7578 1886
rect 7528 1477 7578 1489
rect 7694 1886 7744 1898
rect 7694 1489 7700 1886
rect 7738 1489 7744 1886
rect 7694 1477 7744 1489
rect 7860 1886 7910 1898
rect 7860 1489 7866 1886
rect 7904 1489 7910 1886
rect 7860 1477 7910 1489
rect 8026 1886 8076 1898
rect 8026 1489 8032 1886
rect 8070 1489 8076 1886
rect 8026 1477 8076 1489
rect 8192 1886 8242 1898
rect 8192 1489 8198 1886
rect 8236 1489 8242 1886
rect 8192 1477 8242 1489
rect 8358 1886 8408 1898
rect 8358 1489 8364 1886
rect 8402 1489 8408 1886
rect 8358 1477 8408 1489
rect 8524 1886 8574 1898
rect 8524 1489 8530 1886
rect 8568 1489 8574 1886
rect 8524 1477 8574 1489
rect 8690 1886 8740 1898
rect 8690 1489 8696 1886
rect 8734 1489 8740 1886
rect 8690 1477 8740 1489
rect 8856 1886 8906 1898
rect 8856 1489 8862 1886
rect 8900 1489 8906 1886
rect 8856 1477 8906 1489
rect 9022 1886 9072 1898
rect 9022 1489 9028 1886
rect 9066 1489 9072 1886
rect 9022 1477 9072 1489
rect 9188 1886 9238 1898
rect 9188 1489 9194 1886
rect 9232 1489 9238 1886
rect 9188 1477 9238 1489
rect 9354 1886 9404 1898
rect 9354 1489 9360 1886
rect 9398 1489 9404 1886
rect 9354 1477 9404 1489
rect 9520 1886 9570 1898
rect 9520 1489 9526 1886
rect 9564 1489 9570 1886
rect 9520 1477 9570 1489
rect 9686 1886 9736 1898
rect 9686 1489 9692 1886
rect 9730 1489 9736 1886
rect 9686 1477 9736 1489
rect 9852 1886 9902 1898
rect 9852 1489 9858 1886
rect 9896 1489 9902 1886
rect 9852 1477 9902 1489
rect 10018 1886 10068 1898
rect 10018 1489 10024 1886
rect 10062 1489 10068 1886
rect 10018 1477 10068 1489
rect 10184 1886 10234 1898
rect 10184 1489 10190 1886
rect 10228 1489 10234 1886
rect 10184 1477 10234 1489
rect 10350 1886 10400 1898
rect 10350 1489 10356 1886
rect 10394 1489 10400 1886
rect 10350 1477 10400 1489
rect 10516 1886 10566 1898
rect 10516 1489 10522 1886
rect 10560 1489 10566 1886
rect 10516 1477 10566 1489
rect 10682 1886 10732 1898
rect 10682 1489 10688 1886
rect 10726 1489 10732 1886
rect 10682 1477 10732 1489
rect 10848 1886 10898 1898
rect 10848 1489 10854 1886
rect 10892 1489 10898 1886
rect 10848 1477 10898 1489
rect 11014 1886 11064 1898
rect 11014 1489 11020 1886
rect 11058 1489 11064 1886
rect 11014 1477 11064 1489
rect 11180 1886 11230 1898
rect 11180 1489 11186 1886
rect 11224 1489 11230 1886
rect 11180 1477 11230 1489
rect 11346 1886 11396 1898
rect 11346 1489 11352 1886
rect 11390 1489 11396 1886
rect 11346 1477 11396 1489
rect 11512 1886 11562 1898
rect 11512 1489 11518 1886
rect 11556 1489 11562 1886
rect 11512 1477 11562 1489
rect 11678 1886 11728 1898
rect 11678 1489 11684 1886
rect 11722 1489 11728 1886
rect 11678 1477 11728 1489
rect 11844 1886 11894 1898
rect 11844 1489 11850 1886
rect 11888 1489 11894 1886
rect 11844 1477 11894 1489
rect 12010 1886 12060 1898
rect 12010 1489 12016 1886
rect 12054 1489 12060 1886
rect 12010 1477 12060 1489
rect 12176 1886 12226 1898
rect 12176 1489 12182 1886
rect 12220 1489 12226 1886
rect 12176 1477 12226 1489
rect 12342 1886 12392 1898
rect 12342 1489 12348 1886
rect 12386 1489 12392 1886
rect 12342 1477 12392 1489
rect 12508 1886 12558 1898
rect 12508 1489 12514 1886
rect 12552 1489 12558 1886
rect 12508 1477 12558 1489
rect 12674 1886 12724 1898
rect 12674 1489 12680 1886
rect 12718 1489 12724 1886
rect 12674 1477 12724 1489
rect 12840 1886 12890 1898
rect 12840 1489 12846 1886
rect 12884 1489 12890 1886
rect 12840 1477 12890 1489
rect 13006 1886 13056 1898
rect 13006 1489 13012 1886
rect 13050 1489 13056 1886
rect 13006 1477 13056 1489
rect 13172 1886 13222 1898
rect 13172 1489 13178 1886
rect 13216 1489 13222 1886
rect 13172 1477 13222 1489
rect 13338 1886 13388 1898
rect 13338 1489 13344 1886
rect 13382 1489 13388 1886
rect 13338 1477 13388 1489
rect 13504 1886 13554 1898
rect 13504 1489 13510 1886
rect 13548 1489 13554 1886
rect 13504 1477 13554 1489
rect 13670 1886 13720 1898
rect 13670 1489 13676 1886
rect 13714 1489 13720 1886
rect 13670 1477 13720 1489
rect 13836 1886 13886 1898
rect 13836 1489 13842 1886
rect 13880 1489 13886 1886
rect 13836 1477 13886 1489
rect 14002 1886 14052 1898
rect 14002 1489 14008 1886
rect 14046 1489 14052 1886
rect 14002 1477 14052 1489
rect 14168 1886 14218 1898
rect 14168 1489 14174 1886
rect 14212 1489 14218 1886
rect 14168 1477 14218 1489
rect -14218 -1489 -14168 -1477
rect -14218 -1886 -14212 -1489
rect -14174 -1886 -14168 -1489
rect -14218 -1898 -14168 -1886
rect -14052 -1489 -14002 -1477
rect -14052 -1886 -14046 -1489
rect -14008 -1886 -14002 -1489
rect -14052 -1898 -14002 -1886
rect -13886 -1489 -13836 -1477
rect -13886 -1886 -13880 -1489
rect -13842 -1886 -13836 -1489
rect -13886 -1898 -13836 -1886
rect -13720 -1489 -13670 -1477
rect -13720 -1886 -13714 -1489
rect -13676 -1886 -13670 -1489
rect -13720 -1898 -13670 -1886
rect -13554 -1489 -13504 -1477
rect -13554 -1886 -13548 -1489
rect -13510 -1886 -13504 -1489
rect -13554 -1898 -13504 -1886
rect -13388 -1489 -13338 -1477
rect -13388 -1886 -13382 -1489
rect -13344 -1886 -13338 -1489
rect -13388 -1898 -13338 -1886
rect -13222 -1489 -13172 -1477
rect -13222 -1886 -13216 -1489
rect -13178 -1886 -13172 -1489
rect -13222 -1898 -13172 -1886
rect -13056 -1489 -13006 -1477
rect -13056 -1886 -13050 -1489
rect -13012 -1886 -13006 -1489
rect -13056 -1898 -13006 -1886
rect -12890 -1489 -12840 -1477
rect -12890 -1886 -12884 -1489
rect -12846 -1886 -12840 -1489
rect -12890 -1898 -12840 -1886
rect -12724 -1489 -12674 -1477
rect -12724 -1886 -12718 -1489
rect -12680 -1886 -12674 -1489
rect -12724 -1898 -12674 -1886
rect -12558 -1489 -12508 -1477
rect -12558 -1886 -12552 -1489
rect -12514 -1886 -12508 -1489
rect -12558 -1898 -12508 -1886
rect -12392 -1489 -12342 -1477
rect -12392 -1886 -12386 -1489
rect -12348 -1886 -12342 -1489
rect -12392 -1898 -12342 -1886
rect -12226 -1489 -12176 -1477
rect -12226 -1886 -12220 -1489
rect -12182 -1886 -12176 -1489
rect -12226 -1898 -12176 -1886
rect -12060 -1489 -12010 -1477
rect -12060 -1886 -12054 -1489
rect -12016 -1886 -12010 -1489
rect -12060 -1898 -12010 -1886
rect -11894 -1489 -11844 -1477
rect -11894 -1886 -11888 -1489
rect -11850 -1886 -11844 -1489
rect -11894 -1898 -11844 -1886
rect -11728 -1489 -11678 -1477
rect -11728 -1886 -11722 -1489
rect -11684 -1886 -11678 -1489
rect -11728 -1898 -11678 -1886
rect -11562 -1489 -11512 -1477
rect -11562 -1886 -11556 -1489
rect -11518 -1886 -11512 -1489
rect -11562 -1898 -11512 -1886
rect -11396 -1489 -11346 -1477
rect -11396 -1886 -11390 -1489
rect -11352 -1886 -11346 -1489
rect -11396 -1898 -11346 -1886
rect -11230 -1489 -11180 -1477
rect -11230 -1886 -11224 -1489
rect -11186 -1886 -11180 -1489
rect -11230 -1898 -11180 -1886
rect -11064 -1489 -11014 -1477
rect -11064 -1886 -11058 -1489
rect -11020 -1886 -11014 -1489
rect -11064 -1898 -11014 -1886
rect -10898 -1489 -10848 -1477
rect -10898 -1886 -10892 -1489
rect -10854 -1886 -10848 -1489
rect -10898 -1898 -10848 -1886
rect -10732 -1489 -10682 -1477
rect -10732 -1886 -10726 -1489
rect -10688 -1886 -10682 -1489
rect -10732 -1898 -10682 -1886
rect -10566 -1489 -10516 -1477
rect -10566 -1886 -10560 -1489
rect -10522 -1886 -10516 -1489
rect -10566 -1898 -10516 -1886
rect -10400 -1489 -10350 -1477
rect -10400 -1886 -10394 -1489
rect -10356 -1886 -10350 -1489
rect -10400 -1898 -10350 -1886
rect -10234 -1489 -10184 -1477
rect -10234 -1886 -10228 -1489
rect -10190 -1886 -10184 -1489
rect -10234 -1898 -10184 -1886
rect -10068 -1489 -10018 -1477
rect -10068 -1886 -10062 -1489
rect -10024 -1886 -10018 -1489
rect -10068 -1898 -10018 -1886
rect -9902 -1489 -9852 -1477
rect -9902 -1886 -9896 -1489
rect -9858 -1886 -9852 -1489
rect -9902 -1898 -9852 -1886
rect -9736 -1489 -9686 -1477
rect -9736 -1886 -9730 -1489
rect -9692 -1886 -9686 -1489
rect -9736 -1898 -9686 -1886
rect -9570 -1489 -9520 -1477
rect -9570 -1886 -9564 -1489
rect -9526 -1886 -9520 -1489
rect -9570 -1898 -9520 -1886
rect -9404 -1489 -9354 -1477
rect -9404 -1886 -9398 -1489
rect -9360 -1886 -9354 -1489
rect -9404 -1898 -9354 -1886
rect -9238 -1489 -9188 -1477
rect -9238 -1886 -9232 -1489
rect -9194 -1886 -9188 -1489
rect -9238 -1898 -9188 -1886
rect -9072 -1489 -9022 -1477
rect -9072 -1886 -9066 -1489
rect -9028 -1886 -9022 -1489
rect -9072 -1898 -9022 -1886
rect -8906 -1489 -8856 -1477
rect -8906 -1886 -8900 -1489
rect -8862 -1886 -8856 -1489
rect -8906 -1898 -8856 -1886
rect -8740 -1489 -8690 -1477
rect -8740 -1886 -8734 -1489
rect -8696 -1886 -8690 -1489
rect -8740 -1898 -8690 -1886
rect -8574 -1489 -8524 -1477
rect -8574 -1886 -8568 -1489
rect -8530 -1886 -8524 -1489
rect -8574 -1898 -8524 -1886
rect -8408 -1489 -8358 -1477
rect -8408 -1886 -8402 -1489
rect -8364 -1886 -8358 -1489
rect -8408 -1898 -8358 -1886
rect -8242 -1489 -8192 -1477
rect -8242 -1886 -8236 -1489
rect -8198 -1886 -8192 -1489
rect -8242 -1898 -8192 -1886
rect -8076 -1489 -8026 -1477
rect -8076 -1886 -8070 -1489
rect -8032 -1886 -8026 -1489
rect -8076 -1898 -8026 -1886
rect -7910 -1489 -7860 -1477
rect -7910 -1886 -7904 -1489
rect -7866 -1886 -7860 -1489
rect -7910 -1898 -7860 -1886
rect -7744 -1489 -7694 -1477
rect -7744 -1886 -7738 -1489
rect -7700 -1886 -7694 -1489
rect -7744 -1898 -7694 -1886
rect -7578 -1489 -7528 -1477
rect -7578 -1886 -7572 -1489
rect -7534 -1886 -7528 -1489
rect -7578 -1898 -7528 -1886
rect -7412 -1489 -7362 -1477
rect -7412 -1886 -7406 -1489
rect -7368 -1886 -7362 -1489
rect -7412 -1898 -7362 -1886
rect -7246 -1489 -7196 -1477
rect -7246 -1886 -7240 -1489
rect -7202 -1886 -7196 -1489
rect -7246 -1898 -7196 -1886
rect -7080 -1489 -7030 -1477
rect -7080 -1886 -7074 -1489
rect -7036 -1886 -7030 -1489
rect -7080 -1898 -7030 -1886
rect -6914 -1489 -6864 -1477
rect -6914 -1886 -6908 -1489
rect -6870 -1886 -6864 -1489
rect -6914 -1898 -6864 -1886
rect -6748 -1489 -6698 -1477
rect -6748 -1886 -6742 -1489
rect -6704 -1886 -6698 -1489
rect -6748 -1898 -6698 -1886
rect -6582 -1489 -6532 -1477
rect -6582 -1886 -6576 -1489
rect -6538 -1886 -6532 -1489
rect -6582 -1898 -6532 -1886
rect -6416 -1489 -6366 -1477
rect -6416 -1886 -6410 -1489
rect -6372 -1886 -6366 -1489
rect -6416 -1898 -6366 -1886
rect -6250 -1489 -6200 -1477
rect -6250 -1886 -6244 -1489
rect -6206 -1886 -6200 -1489
rect -6250 -1898 -6200 -1886
rect -6084 -1489 -6034 -1477
rect -6084 -1886 -6078 -1489
rect -6040 -1886 -6034 -1489
rect -6084 -1898 -6034 -1886
rect -5918 -1489 -5868 -1477
rect -5918 -1886 -5912 -1489
rect -5874 -1886 -5868 -1489
rect -5918 -1898 -5868 -1886
rect -5752 -1489 -5702 -1477
rect -5752 -1886 -5746 -1489
rect -5708 -1886 -5702 -1489
rect -5752 -1898 -5702 -1886
rect -5586 -1489 -5536 -1477
rect -5586 -1886 -5580 -1489
rect -5542 -1886 -5536 -1489
rect -5586 -1898 -5536 -1886
rect -5420 -1489 -5370 -1477
rect -5420 -1886 -5414 -1489
rect -5376 -1886 -5370 -1489
rect -5420 -1898 -5370 -1886
rect -5254 -1489 -5204 -1477
rect -5254 -1886 -5248 -1489
rect -5210 -1886 -5204 -1489
rect -5254 -1898 -5204 -1886
rect -5088 -1489 -5038 -1477
rect -5088 -1886 -5082 -1489
rect -5044 -1886 -5038 -1489
rect -5088 -1898 -5038 -1886
rect -4922 -1489 -4872 -1477
rect -4922 -1886 -4916 -1489
rect -4878 -1886 -4872 -1489
rect -4922 -1898 -4872 -1886
rect -4756 -1489 -4706 -1477
rect -4756 -1886 -4750 -1489
rect -4712 -1886 -4706 -1489
rect -4756 -1898 -4706 -1886
rect -4590 -1489 -4540 -1477
rect -4590 -1886 -4584 -1489
rect -4546 -1886 -4540 -1489
rect -4590 -1898 -4540 -1886
rect -4424 -1489 -4374 -1477
rect -4424 -1886 -4418 -1489
rect -4380 -1886 -4374 -1489
rect -4424 -1898 -4374 -1886
rect -4258 -1489 -4208 -1477
rect -4258 -1886 -4252 -1489
rect -4214 -1886 -4208 -1489
rect -4258 -1898 -4208 -1886
rect -4092 -1489 -4042 -1477
rect -4092 -1886 -4086 -1489
rect -4048 -1886 -4042 -1489
rect -4092 -1898 -4042 -1886
rect -3926 -1489 -3876 -1477
rect -3926 -1886 -3920 -1489
rect -3882 -1886 -3876 -1489
rect -3926 -1898 -3876 -1886
rect -3760 -1489 -3710 -1477
rect -3760 -1886 -3754 -1489
rect -3716 -1886 -3710 -1489
rect -3760 -1898 -3710 -1886
rect -3594 -1489 -3544 -1477
rect -3594 -1886 -3588 -1489
rect -3550 -1886 -3544 -1489
rect -3594 -1898 -3544 -1886
rect -3428 -1489 -3378 -1477
rect -3428 -1886 -3422 -1489
rect -3384 -1886 -3378 -1489
rect -3428 -1898 -3378 -1886
rect -3262 -1489 -3212 -1477
rect -3262 -1886 -3256 -1489
rect -3218 -1886 -3212 -1489
rect -3262 -1898 -3212 -1886
rect -3096 -1489 -3046 -1477
rect -3096 -1886 -3090 -1489
rect -3052 -1886 -3046 -1489
rect -3096 -1898 -3046 -1886
rect -2930 -1489 -2880 -1477
rect -2930 -1886 -2924 -1489
rect -2886 -1886 -2880 -1489
rect -2930 -1898 -2880 -1886
rect -2764 -1489 -2714 -1477
rect -2764 -1886 -2758 -1489
rect -2720 -1886 -2714 -1489
rect -2764 -1898 -2714 -1886
rect -2598 -1489 -2548 -1477
rect -2598 -1886 -2592 -1489
rect -2554 -1886 -2548 -1489
rect -2598 -1898 -2548 -1886
rect -2432 -1489 -2382 -1477
rect -2432 -1886 -2426 -1489
rect -2388 -1886 -2382 -1489
rect -2432 -1898 -2382 -1886
rect -2266 -1489 -2216 -1477
rect -2266 -1886 -2260 -1489
rect -2222 -1886 -2216 -1489
rect -2266 -1898 -2216 -1886
rect -2100 -1489 -2050 -1477
rect -2100 -1886 -2094 -1489
rect -2056 -1886 -2050 -1489
rect -2100 -1898 -2050 -1886
rect -1934 -1489 -1884 -1477
rect -1934 -1886 -1928 -1489
rect -1890 -1886 -1884 -1489
rect -1934 -1898 -1884 -1886
rect -1768 -1489 -1718 -1477
rect -1768 -1886 -1762 -1489
rect -1724 -1886 -1718 -1489
rect -1768 -1898 -1718 -1886
rect -1602 -1489 -1552 -1477
rect -1602 -1886 -1596 -1489
rect -1558 -1886 -1552 -1489
rect -1602 -1898 -1552 -1886
rect -1436 -1489 -1386 -1477
rect -1436 -1886 -1430 -1489
rect -1392 -1886 -1386 -1489
rect -1436 -1898 -1386 -1886
rect -1270 -1489 -1220 -1477
rect -1270 -1886 -1264 -1489
rect -1226 -1886 -1220 -1489
rect -1270 -1898 -1220 -1886
rect -1104 -1489 -1054 -1477
rect -1104 -1886 -1098 -1489
rect -1060 -1886 -1054 -1489
rect -1104 -1898 -1054 -1886
rect -938 -1489 -888 -1477
rect -938 -1886 -932 -1489
rect -894 -1886 -888 -1489
rect -938 -1898 -888 -1886
rect -772 -1489 -722 -1477
rect -772 -1886 -766 -1489
rect -728 -1886 -722 -1489
rect -772 -1898 -722 -1886
rect -606 -1489 -556 -1477
rect -606 -1886 -600 -1489
rect -562 -1886 -556 -1489
rect -606 -1898 -556 -1886
rect -440 -1489 -390 -1477
rect -440 -1886 -434 -1489
rect -396 -1886 -390 -1489
rect -440 -1898 -390 -1886
rect -274 -1489 -224 -1477
rect -274 -1886 -268 -1489
rect -230 -1886 -224 -1489
rect -274 -1898 -224 -1886
rect -108 -1489 -58 -1477
rect -108 -1886 -102 -1489
rect -64 -1886 -58 -1489
rect -108 -1898 -58 -1886
rect 58 -1489 108 -1477
rect 58 -1886 64 -1489
rect 102 -1886 108 -1489
rect 58 -1898 108 -1886
rect 224 -1489 274 -1477
rect 224 -1886 230 -1489
rect 268 -1886 274 -1489
rect 224 -1898 274 -1886
rect 390 -1489 440 -1477
rect 390 -1886 396 -1489
rect 434 -1886 440 -1489
rect 390 -1898 440 -1886
rect 556 -1489 606 -1477
rect 556 -1886 562 -1489
rect 600 -1886 606 -1489
rect 556 -1898 606 -1886
rect 722 -1489 772 -1477
rect 722 -1886 728 -1489
rect 766 -1886 772 -1489
rect 722 -1898 772 -1886
rect 888 -1489 938 -1477
rect 888 -1886 894 -1489
rect 932 -1886 938 -1489
rect 888 -1898 938 -1886
rect 1054 -1489 1104 -1477
rect 1054 -1886 1060 -1489
rect 1098 -1886 1104 -1489
rect 1054 -1898 1104 -1886
rect 1220 -1489 1270 -1477
rect 1220 -1886 1226 -1489
rect 1264 -1886 1270 -1489
rect 1220 -1898 1270 -1886
rect 1386 -1489 1436 -1477
rect 1386 -1886 1392 -1489
rect 1430 -1886 1436 -1489
rect 1386 -1898 1436 -1886
rect 1552 -1489 1602 -1477
rect 1552 -1886 1558 -1489
rect 1596 -1886 1602 -1489
rect 1552 -1898 1602 -1886
rect 1718 -1489 1768 -1477
rect 1718 -1886 1724 -1489
rect 1762 -1886 1768 -1489
rect 1718 -1898 1768 -1886
rect 1884 -1489 1934 -1477
rect 1884 -1886 1890 -1489
rect 1928 -1886 1934 -1489
rect 1884 -1898 1934 -1886
rect 2050 -1489 2100 -1477
rect 2050 -1886 2056 -1489
rect 2094 -1886 2100 -1489
rect 2050 -1898 2100 -1886
rect 2216 -1489 2266 -1477
rect 2216 -1886 2222 -1489
rect 2260 -1886 2266 -1489
rect 2216 -1898 2266 -1886
rect 2382 -1489 2432 -1477
rect 2382 -1886 2388 -1489
rect 2426 -1886 2432 -1489
rect 2382 -1898 2432 -1886
rect 2548 -1489 2598 -1477
rect 2548 -1886 2554 -1489
rect 2592 -1886 2598 -1489
rect 2548 -1898 2598 -1886
rect 2714 -1489 2764 -1477
rect 2714 -1886 2720 -1489
rect 2758 -1886 2764 -1489
rect 2714 -1898 2764 -1886
rect 2880 -1489 2930 -1477
rect 2880 -1886 2886 -1489
rect 2924 -1886 2930 -1489
rect 2880 -1898 2930 -1886
rect 3046 -1489 3096 -1477
rect 3046 -1886 3052 -1489
rect 3090 -1886 3096 -1489
rect 3046 -1898 3096 -1886
rect 3212 -1489 3262 -1477
rect 3212 -1886 3218 -1489
rect 3256 -1886 3262 -1489
rect 3212 -1898 3262 -1886
rect 3378 -1489 3428 -1477
rect 3378 -1886 3384 -1489
rect 3422 -1886 3428 -1489
rect 3378 -1898 3428 -1886
rect 3544 -1489 3594 -1477
rect 3544 -1886 3550 -1489
rect 3588 -1886 3594 -1489
rect 3544 -1898 3594 -1886
rect 3710 -1489 3760 -1477
rect 3710 -1886 3716 -1489
rect 3754 -1886 3760 -1489
rect 3710 -1898 3760 -1886
rect 3876 -1489 3926 -1477
rect 3876 -1886 3882 -1489
rect 3920 -1886 3926 -1489
rect 3876 -1898 3926 -1886
rect 4042 -1489 4092 -1477
rect 4042 -1886 4048 -1489
rect 4086 -1886 4092 -1489
rect 4042 -1898 4092 -1886
rect 4208 -1489 4258 -1477
rect 4208 -1886 4214 -1489
rect 4252 -1886 4258 -1489
rect 4208 -1898 4258 -1886
rect 4374 -1489 4424 -1477
rect 4374 -1886 4380 -1489
rect 4418 -1886 4424 -1489
rect 4374 -1898 4424 -1886
rect 4540 -1489 4590 -1477
rect 4540 -1886 4546 -1489
rect 4584 -1886 4590 -1489
rect 4540 -1898 4590 -1886
rect 4706 -1489 4756 -1477
rect 4706 -1886 4712 -1489
rect 4750 -1886 4756 -1489
rect 4706 -1898 4756 -1886
rect 4872 -1489 4922 -1477
rect 4872 -1886 4878 -1489
rect 4916 -1886 4922 -1489
rect 4872 -1898 4922 -1886
rect 5038 -1489 5088 -1477
rect 5038 -1886 5044 -1489
rect 5082 -1886 5088 -1489
rect 5038 -1898 5088 -1886
rect 5204 -1489 5254 -1477
rect 5204 -1886 5210 -1489
rect 5248 -1886 5254 -1489
rect 5204 -1898 5254 -1886
rect 5370 -1489 5420 -1477
rect 5370 -1886 5376 -1489
rect 5414 -1886 5420 -1489
rect 5370 -1898 5420 -1886
rect 5536 -1489 5586 -1477
rect 5536 -1886 5542 -1489
rect 5580 -1886 5586 -1489
rect 5536 -1898 5586 -1886
rect 5702 -1489 5752 -1477
rect 5702 -1886 5708 -1489
rect 5746 -1886 5752 -1489
rect 5702 -1898 5752 -1886
rect 5868 -1489 5918 -1477
rect 5868 -1886 5874 -1489
rect 5912 -1886 5918 -1489
rect 5868 -1898 5918 -1886
rect 6034 -1489 6084 -1477
rect 6034 -1886 6040 -1489
rect 6078 -1886 6084 -1489
rect 6034 -1898 6084 -1886
rect 6200 -1489 6250 -1477
rect 6200 -1886 6206 -1489
rect 6244 -1886 6250 -1489
rect 6200 -1898 6250 -1886
rect 6366 -1489 6416 -1477
rect 6366 -1886 6372 -1489
rect 6410 -1886 6416 -1489
rect 6366 -1898 6416 -1886
rect 6532 -1489 6582 -1477
rect 6532 -1886 6538 -1489
rect 6576 -1886 6582 -1489
rect 6532 -1898 6582 -1886
rect 6698 -1489 6748 -1477
rect 6698 -1886 6704 -1489
rect 6742 -1886 6748 -1489
rect 6698 -1898 6748 -1886
rect 6864 -1489 6914 -1477
rect 6864 -1886 6870 -1489
rect 6908 -1886 6914 -1489
rect 6864 -1898 6914 -1886
rect 7030 -1489 7080 -1477
rect 7030 -1886 7036 -1489
rect 7074 -1886 7080 -1489
rect 7030 -1898 7080 -1886
rect 7196 -1489 7246 -1477
rect 7196 -1886 7202 -1489
rect 7240 -1886 7246 -1489
rect 7196 -1898 7246 -1886
rect 7362 -1489 7412 -1477
rect 7362 -1886 7368 -1489
rect 7406 -1886 7412 -1489
rect 7362 -1898 7412 -1886
rect 7528 -1489 7578 -1477
rect 7528 -1886 7534 -1489
rect 7572 -1886 7578 -1489
rect 7528 -1898 7578 -1886
rect 7694 -1489 7744 -1477
rect 7694 -1886 7700 -1489
rect 7738 -1886 7744 -1489
rect 7694 -1898 7744 -1886
rect 7860 -1489 7910 -1477
rect 7860 -1886 7866 -1489
rect 7904 -1886 7910 -1489
rect 7860 -1898 7910 -1886
rect 8026 -1489 8076 -1477
rect 8026 -1886 8032 -1489
rect 8070 -1886 8076 -1489
rect 8026 -1898 8076 -1886
rect 8192 -1489 8242 -1477
rect 8192 -1886 8198 -1489
rect 8236 -1886 8242 -1489
rect 8192 -1898 8242 -1886
rect 8358 -1489 8408 -1477
rect 8358 -1886 8364 -1489
rect 8402 -1886 8408 -1489
rect 8358 -1898 8408 -1886
rect 8524 -1489 8574 -1477
rect 8524 -1886 8530 -1489
rect 8568 -1886 8574 -1489
rect 8524 -1898 8574 -1886
rect 8690 -1489 8740 -1477
rect 8690 -1886 8696 -1489
rect 8734 -1886 8740 -1489
rect 8690 -1898 8740 -1886
rect 8856 -1489 8906 -1477
rect 8856 -1886 8862 -1489
rect 8900 -1886 8906 -1489
rect 8856 -1898 8906 -1886
rect 9022 -1489 9072 -1477
rect 9022 -1886 9028 -1489
rect 9066 -1886 9072 -1489
rect 9022 -1898 9072 -1886
rect 9188 -1489 9238 -1477
rect 9188 -1886 9194 -1489
rect 9232 -1886 9238 -1489
rect 9188 -1898 9238 -1886
rect 9354 -1489 9404 -1477
rect 9354 -1886 9360 -1489
rect 9398 -1886 9404 -1489
rect 9354 -1898 9404 -1886
rect 9520 -1489 9570 -1477
rect 9520 -1886 9526 -1489
rect 9564 -1886 9570 -1489
rect 9520 -1898 9570 -1886
rect 9686 -1489 9736 -1477
rect 9686 -1886 9692 -1489
rect 9730 -1886 9736 -1489
rect 9686 -1898 9736 -1886
rect 9852 -1489 9902 -1477
rect 9852 -1886 9858 -1489
rect 9896 -1886 9902 -1489
rect 9852 -1898 9902 -1886
rect 10018 -1489 10068 -1477
rect 10018 -1886 10024 -1489
rect 10062 -1886 10068 -1489
rect 10018 -1898 10068 -1886
rect 10184 -1489 10234 -1477
rect 10184 -1886 10190 -1489
rect 10228 -1886 10234 -1489
rect 10184 -1898 10234 -1886
rect 10350 -1489 10400 -1477
rect 10350 -1886 10356 -1489
rect 10394 -1886 10400 -1489
rect 10350 -1898 10400 -1886
rect 10516 -1489 10566 -1477
rect 10516 -1886 10522 -1489
rect 10560 -1886 10566 -1489
rect 10516 -1898 10566 -1886
rect 10682 -1489 10732 -1477
rect 10682 -1886 10688 -1489
rect 10726 -1886 10732 -1489
rect 10682 -1898 10732 -1886
rect 10848 -1489 10898 -1477
rect 10848 -1886 10854 -1489
rect 10892 -1886 10898 -1489
rect 10848 -1898 10898 -1886
rect 11014 -1489 11064 -1477
rect 11014 -1886 11020 -1489
rect 11058 -1886 11064 -1489
rect 11014 -1898 11064 -1886
rect 11180 -1489 11230 -1477
rect 11180 -1886 11186 -1489
rect 11224 -1886 11230 -1489
rect 11180 -1898 11230 -1886
rect 11346 -1489 11396 -1477
rect 11346 -1886 11352 -1489
rect 11390 -1886 11396 -1489
rect 11346 -1898 11396 -1886
rect 11512 -1489 11562 -1477
rect 11512 -1886 11518 -1489
rect 11556 -1886 11562 -1489
rect 11512 -1898 11562 -1886
rect 11678 -1489 11728 -1477
rect 11678 -1886 11684 -1489
rect 11722 -1886 11728 -1489
rect 11678 -1898 11728 -1886
rect 11844 -1489 11894 -1477
rect 11844 -1886 11850 -1489
rect 11888 -1886 11894 -1489
rect 11844 -1898 11894 -1886
rect 12010 -1489 12060 -1477
rect 12010 -1886 12016 -1489
rect 12054 -1886 12060 -1489
rect 12010 -1898 12060 -1886
rect 12176 -1489 12226 -1477
rect 12176 -1886 12182 -1489
rect 12220 -1886 12226 -1489
rect 12176 -1898 12226 -1886
rect 12342 -1489 12392 -1477
rect 12342 -1886 12348 -1489
rect 12386 -1886 12392 -1489
rect 12342 -1898 12392 -1886
rect 12508 -1489 12558 -1477
rect 12508 -1886 12514 -1489
rect 12552 -1886 12558 -1489
rect 12508 -1898 12558 -1886
rect 12674 -1489 12724 -1477
rect 12674 -1886 12680 -1489
rect 12718 -1886 12724 -1489
rect 12674 -1898 12724 -1886
rect 12840 -1489 12890 -1477
rect 12840 -1886 12846 -1489
rect 12884 -1886 12890 -1489
rect 12840 -1898 12890 -1886
rect 13006 -1489 13056 -1477
rect 13006 -1886 13012 -1489
rect 13050 -1886 13056 -1489
rect 13006 -1898 13056 -1886
rect 13172 -1489 13222 -1477
rect 13172 -1886 13178 -1489
rect 13216 -1886 13222 -1489
rect 13172 -1898 13222 -1886
rect 13338 -1489 13388 -1477
rect 13338 -1886 13344 -1489
rect 13382 -1886 13388 -1489
rect 13338 -1898 13388 -1886
rect 13504 -1489 13554 -1477
rect 13504 -1886 13510 -1489
rect 13548 -1886 13554 -1489
rect 13504 -1898 13554 -1886
rect 13670 -1489 13720 -1477
rect 13670 -1886 13676 -1489
rect 13714 -1886 13720 -1489
rect 13670 -1898 13720 -1886
rect 13836 -1489 13886 -1477
rect 13836 -1886 13842 -1489
rect 13880 -1886 13886 -1489
rect 13836 -1898 13886 -1886
rect 14002 -1489 14052 -1477
rect 14002 -1886 14008 -1489
rect 14046 -1886 14052 -1489
rect 14002 -1898 14052 -1886
rect 14168 -1489 14218 -1477
rect 14168 -1886 14174 -1489
rect 14212 -1886 14218 -1489
rect 14168 -1898 14218 -1886
<< properties >>
string FIXED_BBOX -14341 -2017 14341 2017
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 14.88 m 1 nx 172 wmin 0.350 lmin 0.50 class resistor rho 2000 val 86.104k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
