magic
tech sky130A
magscale 1 2
timestamp 1730992408
<< pwell >>
rect -3295 -2978 3295 2978
<< mvnmos >>
rect -3067 1720 -2867 2720
rect -2809 1720 -2609 2720
rect -2551 1720 -2351 2720
rect -2293 1720 -2093 2720
rect -2035 1720 -1835 2720
rect -1777 1720 -1577 2720
rect -1519 1720 -1319 2720
rect -1261 1720 -1061 2720
rect -1003 1720 -803 2720
rect -745 1720 -545 2720
rect -487 1720 -287 2720
rect -229 1720 -29 2720
rect 29 1720 229 2720
rect 287 1720 487 2720
rect 545 1720 745 2720
rect 803 1720 1003 2720
rect 1061 1720 1261 2720
rect 1319 1720 1519 2720
rect 1577 1720 1777 2720
rect 1835 1720 2035 2720
rect 2093 1720 2293 2720
rect 2351 1720 2551 2720
rect 2609 1720 2809 2720
rect 2867 1720 3067 2720
rect -3067 610 -2867 1610
rect -2809 610 -2609 1610
rect -2551 610 -2351 1610
rect -2293 610 -2093 1610
rect -2035 610 -1835 1610
rect -1777 610 -1577 1610
rect -1519 610 -1319 1610
rect -1261 610 -1061 1610
rect -1003 610 -803 1610
rect -745 610 -545 1610
rect -487 610 -287 1610
rect -229 610 -29 1610
rect 29 610 229 1610
rect 287 610 487 1610
rect 545 610 745 1610
rect 803 610 1003 1610
rect 1061 610 1261 1610
rect 1319 610 1519 1610
rect 1577 610 1777 1610
rect 1835 610 2035 1610
rect 2093 610 2293 1610
rect 2351 610 2551 1610
rect 2609 610 2809 1610
rect 2867 610 3067 1610
rect -3067 -500 -2867 500
rect -2809 -500 -2609 500
rect -2551 -500 -2351 500
rect -2293 -500 -2093 500
rect -2035 -500 -1835 500
rect -1777 -500 -1577 500
rect -1519 -500 -1319 500
rect -1261 -500 -1061 500
rect -1003 -500 -803 500
rect -745 -500 -545 500
rect -487 -500 -287 500
rect -229 -500 -29 500
rect 29 -500 229 500
rect 287 -500 487 500
rect 545 -500 745 500
rect 803 -500 1003 500
rect 1061 -500 1261 500
rect 1319 -500 1519 500
rect 1577 -500 1777 500
rect 1835 -500 2035 500
rect 2093 -500 2293 500
rect 2351 -500 2551 500
rect 2609 -500 2809 500
rect 2867 -500 3067 500
rect -3067 -1610 -2867 -610
rect -2809 -1610 -2609 -610
rect -2551 -1610 -2351 -610
rect -2293 -1610 -2093 -610
rect -2035 -1610 -1835 -610
rect -1777 -1610 -1577 -610
rect -1519 -1610 -1319 -610
rect -1261 -1610 -1061 -610
rect -1003 -1610 -803 -610
rect -745 -1610 -545 -610
rect -487 -1610 -287 -610
rect -229 -1610 -29 -610
rect 29 -1610 229 -610
rect 287 -1610 487 -610
rect 545 -1610 745 -610
rect 803 -1610 1003 -610
rect 1061 -1610 1261 -610
rect 1319 -1610 1519 -610
rect 1577 -1610 1777 -610
rect 1835 -1610 2035 -610
rect 2093 -1610 2293 -610
rect 2351 -1610 2551 -610
rect 2609 -1610 2809 -610
rect 2867 -1610 3067 -610
rect -3067 -2720 -2867 -1720
rect -2809 -2720 -2609 -1720
rect -2551 -2720 -2351 -1720
rect -2293 -2720 -2093 -1720
rect -2035 -2720 -1835 -1720
rect -1777 -2720 -1577 -1720
rect -1519 -2720 -1319 -1720
rect -1261 -2720 -1061 -1720
rect -1003 -2720 -803 -1720
rect -745 -2720 -545 -1720
rect -487 -2720 -287 -1720
rect -229 -2720 -29 -1720
rect 29 -2720 229 -1720
rect 287 -2720 487 -1720
rect 545 -2720 745 -1720
rect 803 -2720 1003 -1720
rect 1061 -2720 1261 -1720
rect 1319 -2720 1519 -1720
rect 1577 -2720 1777 -1720
rect 1835 -2720 2035 -1720
rect 2093 -2720 2293 -1720
rect 2351 -2720 2551 -1720
rect 2609 -2720 2809 -1720
rect 2867 -2720 3067 -1720
<< mvndiff >>
rect -3125 2708 -3067 2720
rect -3125 1732 -3113 2708
rect -3079 1732 -3067 2708
rect -3125 1720 -3067 1732
rect -2867 2708 -2809 2720
rect -2867 1732 -2855 2708
rect -2821 1732 -2809 2708
rect -2867 1720 -2809 1732
rect -2609 2708 -2551 2720
rect -2609 1732 -2597 2708
rect -2563 1732 -2551 2708
rect -2609 1720 -2551 1732
rect -2351 2708 -2293 2720
rect -2351 1732 -2339 2708
rect -2305 1732 -2293 2708
rect -2351 1720 -2293 1732
rect -2093 2708 -2035 2720
rect -2093 1732 -2081 2708
rect -2047 1732 -2035 2708
rect -2093 1720 -2035 1732
rect -1835 2708 -1777 2720
rect -1835 1732 -1823 2708
rect -1789 1732 -1777 2708
rect -1835 1720 -1777 1732
rect -1577 2708 -1519 2720
rect -1577 1732 -1565 2708
rect -1531 1732 -1519 2708
rect -1577 1720 -1519 1732
rect -1319 2708 -1261 2720
rect -1319 1732 -1307 2708
rect -1273 1732 -1261 2708
rect -1319 1720 -1261 1732
rect -1061 2708 -1003 2720
rect -1061 1732 -1049 2708
rect -1015 1732 -1003 2708
rect -1061 1720 -1003 1732
rect -803 2708 -745 2720
rect -803 1732 -791 2708
rect -757 1732 -745 2708
rect -803 1720 -745 1732
rect -545 2708 -487 2720
rect -545 1732 -533 2708
rect -499 1732 -487 2708
rect -545 1720 -487 1732
rect -287 2708 -229 2720
rect -287 1732 -275 2708
rect -241 1732 -229 2708
rect -287 1720 -229 1732
rect -29 2708 29 2720
rect -29 1732 -17 2708
rect 17 1732 29 2708
rect -29 1720 29 1732
rect 229 2708 287 2720
rect 229 1732 241 2708
rect 275 1732 287 2708
rect 229 1720 287 1732
rect 487 2708 545 2720
rect 487 1732 499 2708
rect 533 1732 545 2708
rect 487 1720 545 1732
rect 745 2708 803 2720
rect 745 1732 757 2708
rect 791 1732 803 2708
rect 745 1720 803 1732
rect 1003 2708 1061 2720
rect 1003 1732 1015 2708
rect 1049 1732 1061 2708
rect 1003 1720 1061 1732
rect 1261 2708 1319 2720
rect 1261 1732 1273 2708
rect 1307 1732 1319 2708
rect 1261 1720 1319 1732
rect 1519 2708 1577 2720
rect 1519 1732 1531 2708
rect 1565 1732 1577 2708
rect 1519 1720 1577 1732
rect 1777 2708 1835 2720
rect 1777 1732 1789 2708
rect 1823 1732 1835 2708
rect 1777 1720 1835 1732
rect 2035 2708 2093 2720
rect 2035 1732 2047 2708
rect 2081 1732 2093 2708
rect 2035 1720 2093 1732
rect 2293 2708 2351 2720
rect 2293 1732 2305 2708
rect 2339 1732 2351 2708
rect 2293 1720 2351 1732
rect 2551 2708 2609 2720
rect 2551 1732 2563 2708
rect 2597 1732 2609 2708
rect 2551 1720 2609 1732
rect 2809 2708 2867 2720
rect 2809 1732 2821 2708
rect 2855 1732 2867 2708
rect 2809 1720 2867 1732
rect 3067 2708 3125 2720
rect 3067 1732 3079 2708
rect 3113 1732 3125 2708
rect 3067 1720 3125 1732
rect -3125 1598 -3067 1610
rect -3125 622 -3113 1598
rect -3079 622 -3067 1598
rect -3125 610 -3067 622
rect -2867 1598 -2809 1610
rect -2867 622 -2855 1598
rect -2821 622 -2809 1598
rect -2867 610 -2809 622
rect -2609 1598 -2551 1610
rect -2609 622 -2597 1598
rect -2563 622 -2551 1598
rect -2609 610 -2551 622
rect -2351 1598 -2293 1610
rect -2351 622 -2339 1598
rect -2305 622 -2293 1598
rect -2351 610 -2293 622
rect -2093 1598 -2035 1610
rect -2093 622 -2081 1598
rect -2047 622 -2035 1598
rect -2093 610 -2035 622
rect -1835 1598 -1777 1610
rect -1835 622 -1823 1598
rect -1789 622 -1777 1598
rect -1835 610 -1777 622
rect -1577 1598 -1519 1610
rect -1577 622 -1565 1598
rect -1531 622 -1519 1598
rect -1577 610 -1519 622
rect -1319 1598 -1261 1610
rect -1319 622 -1307 1598
rect -1273 622 -1261 1598
rect -1319 610 -1261 622
rect -1061 1598 -1003 1610
rect -1061 622 -1049 1598
rect -1015 622 -1003 1598
rect -1061 610 -1003 622
rect -803 1598 -745 1610
rect -803 622 -791 1598
rect -757 622 -745 1598
rect -803 610 -745 622
rect -545 1598 -487 1610
rect -545 622 -533 1598
rect -499 622 -487 1598
rect -545 610 -487 622
rect -287 1598 -229 1610
rect -287 622 -275 1598
rect -241 622 -229 1598
rect -287 610 -229 622
rect -29 1598 29 1610
rect -29 622 -17 1598
rect 17 622 29 1598
rect -29 610 29 622
rect 229 1598 287 1610
rect 229 622 241 1598
rect 275 622 287 1598
rect 229 610 287 622
rect 487 1598 545 1610
rect 487 622 499 1598
rect 533 622 545 1598
rect 487 610 545 622
rect 745 1598 803 1610
rect 745 622 757 1598
rect 791 622 803 1598
rect 745 610 803 622
rect 1003 1598 1061 1610
rect 1003 622 1015 1598
rect 1049 622 1061 1598
rect 1003 610 1061 622
rect 1261 1598 1319 1610
rect 1261 622 1273 1598
rect 1307 622 1319 1598
rect 1261 610 1319 622
rect 1519 1598 1577 1610
rect 1519 622 1531 1598
rect 1565 622 1577 1598
rect 1519 610 1577 622
rect 1777 1598 1835 1610
rect 1777 622 1789 1598
rect 1823 622 1835 1598
rect 1777 610 1835 622
rect 2035 1598 2093 1610
rect 2035 622 2047 1598
rect 2081 622 2093 1598
rect 2035 610 2093 622
rect 2293 1598 2351 1610
rect 2293 622 2305 1598
rect 2339 622 2351 1598
rect 2293 610 2351 622
rect 2551 1598 2609 1610
rect 2551 622 2563 1598
rect 2597 622 2609 1598
rect 2551 610 2609 622
rect 2809 1598 2867 1610
rect 2809 622 2821 1598
rect 2855 622 2867 1598
rect 2809 610 2867 622
rect 3067 1598 3125 1610
rect 3067 622 3079 1598
rect 3113 622 3125 1598
rect 3067 610 3125 622
rect -3125 488 -3067 500
rect -3125 -488 -3113 488
rect -3079 -488 -3067 488
rect -3125 -500 -3067 -488
rect -2867 488 -2809 500
rect -2867 -488 -2855 488
rect -2821 -488 -2809 488
rect -2867 -500 -2809 -488
rect -2609 488 -2551 500
rect -2609 -488 -2597 488
rect -2563 -488 -2551 488
rect -2609 -500 -2551 -488
rect -2351 488 -2293 500
rect -2351 -488 -2339 488
rect -2305 -488 -2293 488
rect -2351 -500 -2293 -488
rect -2093 488 -2035 500
rect -2093 -488 -2081 488
rect -2047 -488 -2035 488
rect -2093 -500 -2035 -488
rect -1835 488 -1777 500
rect -1835 -488 -1823 488
rect -1789 -488 -1777 488
rect -1835 -500 -1777 -488
rect -1577 488 -1519 500
rect -1577 -488 -1565 488
rect -1531 -488 -1519 488
rect -1577 -500 -1519 -488
rect -1319 488 -1261 500
rect -1319 -488 -1307 488
rect -1273 -488 -1261 488
rect -1319 -500 -1261 -488
rect -1061 488 -1003 500
rect -1061 -488 -1049 488
rect -1015 -488 -1003 488
rect -1061 -500 -1003 -488
rect -803 488 -745 500
rect -803 -488 -791 488
rect -757 -488 -745 488
rect -803 -500 -745 -488
rect -545 488 -487 500
rect -545 -488 -533 488
rect -499 -488 -487 488
rect -545 -500 -487 -488
rect -287 488 -229 500
rect -287 -488 -275 488
rect -241 -488 -229 488
rect -287 -500 -229 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 229 488 287 500
rect 229 -488 241 488
rect 275 -488 287 488
rect 229 -500 287 -488
rect 487 488 545 500
rect 487 -488 499 488
rect 533 -488 545 488
rect 487 -500 545 -488
rect 745 488 803 500
rect 745 -488 757 488
rect 791 -488 803 488
rect 745 -500 803 -488
rect 1003 488 1061 500
rect 1003 -488 1015 488
rect 1049 -488 1061 488
rect 1003 -500 1061 -488
rect 1261 488 1319 500
rect 1261 -488 1273 488
rect 1307 -488 1319 488
rect 1261 -500 1319 -488
rect 1519 488 1577 500
rect 1519 -488 1531 488
rect 1565 -488 1577 488
rect 1519 -500 1577 -488
rect 1777 488 1835 500
rect 1777 -488 1789 488
rect 1823 -488 1835 488
rect 1777 -500 1835 -488
rect 2035 488 2093 500
rect 2035 -488 2047 488
rect 2081 -488 2093 488
rect 2035 -500 2093 -488
rect 2293 488 2351 500
rect 2293 -488 2305 488
rect 2339 -488 2351 488
rect 2293 -500 2351 -488
rect 2551 488 2609 500
rect 2551 -488 2563 488
rect 2597 -488 2609 488
rect 2551 -500 2609 -488
rect 2809 488 2867 500
rect 2809 -488 2821 488
rect 2855 -488 2867 488
rect 2809 -500 2867 -488
rect 3067 488 3125 500
rect 3067 -488 3079 488
rect 3113 -488 3125 488
rect 3067 -500 3125 -488
rect -3125 -622 -3067 -610
rect -3125 -1598 -3113 -622
rect -3079 -1598 -3067 -622
rect -3125 -1610 -3067 -1598
rect -2867 -622 -2809 -610
rect -2867 -1598 -2855 -622
rect -2821 -1598 -2809 -622
rect -2867 -1610 -2809 -1598
rect -2609 -622 -2551 -610
rect -2609 -1598 -2597 -622
rect -2563 -1598 -2551 -622
rect -2609 -1610 -2551 -1598
rect -2351 -622 -2293 -610
rect -2351 -1598 -2339 -622
rect -2305 -1598 -2293 -622
rect -2351 -1610 -2293 -1598
rect -2093 -622 -2035 -610
rect -2093 -1598 -2081 -622
rect -2047 -1598 -2035 -622
rect -2093 -1610 -2035 -1598
rect -1835 -622 -1777 -610
rect -1835 -1598 -1823 -622
rect -1789 -1598 -1777 -622
rect -1835 -1610 -1777 -1598
rect -1577 -622 -1519 -610
rect -1577 -1598 -1565 -622
rect -1531 -1598 -1519 -622
rect -1577 -1610 -1519 -1598
rect -1319 -622 -1261 -610
rect -1319 -1598 -1307 -622
rect -1273 -1598 -1261 -622
rect -1319 -1610 -1261 -1598
rect -1061 -622 -1003 -610
rect -1061 -1598 -1049 -622
rect -1015 -1598 -1003 -622
rect -1061 -1610 -1003 -1598
rect -803 -622 -745 -610
rect -803 -1598 -791 -622
rect -757 -1598 -745 -622
rect -803 -1610 -745 -1598
rect -545 -622 -487 -610
rect -545 -1598 -533 -622
rect -499 -1598 -487 -622
rect -545 -1610 -487 -1598
rect -287 -622 -229 -610
rect -287 -1598 -275 -622
rect -241 -1598 -229 -622
rect -287 -1610 -229 -1598
rect -29 -622 29 -610
rect -29 -1598 -17 -622
rect 17 -1598 29 -622
rect -29 -1610 29 -1598
rect 229 -622 287 -610
rect 229 -1598 241 -622
rect 275 -1598 287 -622
rect 229 -1610 287 -1598
rect 487 -622 545 -610
rect 487 -1598 499 -622
rect 533 -1598 545 -622
rect 487 -1610 545 -1598
rect 745 -622 803 -610
rect 745 -1598 757 -622
rect 791 -1598 803 -622
rect 745 -1610 803 -1598
rect 1003 -622 1061 -610
rect 1003 -1598 1015 -622
rect 1049 -1598 1061 -622
rect 1003 -1610 1061 -1598
rect 1261 -622 1319 -610
rect 1261 -1598 1273 -622
rect 1307 -1598 1319 -622
rect 1261 -1610 1319 -1598
rect 1519 -622 1577 -610
rect 1519 -1598 1531 -622
rect 1565 -1598 1577 -622
rect 1519 -1610 1577 -1598
rect 1777 -622 1835 -610
rect 1777 -1598 1789 -622
rect 1823 -1598 1835 -622
rect 1777 -1610 1835 -1598
rect 2035 -622 2093 -610
rect 2035 -1598 2047 -622
rect 2081 -1598 2093 -622
rect 2035 -1610 2093 -1598
rect 2293 -622 2351 -610
rect 2293 -1598 2305 -622
rect 2339 -1598 2351 -622
rect 2293 -1610 2351 -1598
rect 2551 -622 2609 -610
rect 2551 -1598 2563 -622
rect 2597 -1598 2609 -622
rect 2551 -1610 2609 -1598
rect 2809 -622 2867 -610
rect 2809 -1598 2821 -622
rect 2855 -1598 2867 -622
rect 2809 -1610 2867 -1598
rect 3067 -622 3125 -610
rect 3067 -1598 3079 -622
rect 3113 -1598 3125 -622
rect 3067 -1610 3125 -1598
rect -3125 -1732 -3067 -1720
rect -3125 -2708 -3113 -1732
rect -3079 -2708 -3067 -1732
rect -3125 -2720 -3067 -2708
rect -2867 -1732 -2809 -1720
rect -2867 -2708 -2855 -1732
rect -2821 -2708 -2809 -1732
rect -2867 -2720 -2809 -2708
rect -2609 -1732 -2551 -1720
rect -2609 -2708 -2597 -1732
rect -2563 -2708 -2551 -1732
rect -2609 -2720 -2551 -2708
rect -2351 -1732 -2293 -1720
rect -2351 -2708 -2339 -1732
rect -2305 -2708 -2293 -1732
rect -2351 -2720 -2293 -2708
rect -2093 -1732 -2035 -1720
rect -2093 -2708 -2081 -1732
rect -2047 -2708 -2035 -1732
rect -2093 -2720 -2035 -2708
rect -1835 -1732 -1777 -1720
rect -1835 -2708 -1823 -1732
rect -1789 -2708 -1777 -1732
rect -1835 -2720 -1777 -2708
rect -1577 -1732 -1519 -1720
rect -1577 -2708 -1565 -1732
rect -1531 -2708 -1519 -1732
rect -1577 -2720 -1519 -2708
rect -1319 -1732 -1261 -1720
rect -1319 -2708 -1307 -1732
rect -1273 -2708 -1261 -1732
rect -1319 -2720 -1261 -2708
rect -1061 -1732 -1003 -1720
rect -1061 -2708 -1049 -1732
rect -1015 -2708 -1003 -1732
rect -1061 -2720 -1003 -2708
rect -803 -1732 -745 -1720
rect -803 -2708 -791 -1732
rect -757 -2708 -745 -1732
rect -803 -2720 -745 -2708
rect -545 -1732 -487 -1720
rect -545 -2708 -533 -1732
rect -499 -2708 -487 -1732
rect -545 -2720 -487 -2708
rect -287 -1732 -229 -1720
rect -287 -2708 -275 -1732
rect -241 -2708 -229 -1732
rect -287 -2720 -229 -2708
rect -29 -1732 29 -1720
rect -29 -2708 -17 -1732
rect 17 -2708 29 -1732
rect -29 -2720 29 -2708
rect 229 -1732 287 -1720
rect 229 -2708 241 -1732
rect 275 -2708 287 -1732
rect 229 -2720 287 -2708
rect 487 -1732 545 -1720
rect 487 -2708 499 -1732
rect 533 -2708 545 -1732
rect 487 -2720 545 -2708
rect 745 -1732 803 -1720
rect 745 -2708 757 -1732
rect 791 -2708 803 -1732
rect 745 -2720 803 -2708
rect 1003 -1732 1061 -1720
rect 1003 -2708 1015 -1732
rect 1049 -2708 1061 -1732
rect 1003 -2720 1061 -2708
rect 1261 -1732 1319 -1720
rect 1261 -2708 1273 -1732
rect 1307 -2708 1319 -1732
rect 1261 -2720 1319 -2708
rect 1519 -1732 1577 -1720
rect 1519 -2708 1531 -1732
rect 1565 -2708 1577 -1732
rect 1519 -2720 1577 -2708
rect 1777 -1732 1835 -1720
rect 1777 -2708 1789 -1732
rect 1823 -2708 1835 -1732
rect 1777 -2720 1835 -2708
rect 2035 -1732 2093 -1720
rect 2035 -2708 2047 -1732
rect 2081 -2708 2093 -1732
rect 2035 -2720 2093 -2708
rect 2293 -1732 2351 -1720
rect 2293 -2708 2305 -1732
rect 2339 -2708 2351 -1732
rect 2293 -2720 2351 -2708
rect 2551 -1732 2609 -1720
rect 2551 -2708 2563 -1732
rect 2597 -2708 2609 -1732
rect 2551 -2720 2609 -2708
rect 2809 -1732 2867 -1720
rect 2809 -2708 2821 -1732
rect 2855 -2708 2867 -1732
rect 2809 -2720 2867 -2708
rect 3067 -1732 3125 -1720
rect 3067 -2708 3079 -1732
rect 3113 -2708 3125 -1732
rect 3067 -2720 3125 -2708
<< mvndiffc >>
rect -3113 1732 -3079 2708
rect -2855 1732 -2821 2708
rect -2597 1732 -2563 2708
rect -2339 1732 -2305 2708
rect -2081 1732 -2047 2708
rect -1823 1732 -1789 2708
rect -1565 1732 -1531 2708
rect -1307 1732 -1273 2708
rect -1049 1732 -1015 2708
rect -791 1732 -757 2708
rect -533 1732 -499 2708
rect -275 1732 -241 2708
rect -17 1732 17 2708
rect 241 1732 275 2708
rect 499 1732 533 2708
rect 757 1732 791 2708
rect 1015 1732 1049 2708
rect 1273 1732 1307 2708
rect 1531 1732 1565 2708
rect 1789 1732 1823 2708
rect 2047 1732 2081 2708
rect 2305 1732 2339 2708
rect 2563 1732 2597 2708
rect 2821 1732 2855 2708
rect 3079 1732 3113 2708
rect -3113 622 -3079 1598
rect -2855 622 -2821 1598
rect -2597 622 -2563 1598
rect -2339 622 -2305 1598
rect -2081 622 -2047 1598
rect -1823 622 -1789 1598
rect -1565 622 -1531 1598
rect -1307 622 -1273 1598
rect -1049 622 -1015 1598
rect -791 622 -757 1598
rect -533 622 -499 1598
rect -275 622 -241 1598
rect -17 622 17 1598
rect 241 622 275 1598
rect 499 622 533 1598
rect 757 622 791 1598
rect 1015 622 1049 1598
rect 1273 622 1307 1598
rect 1531 622 1565 1598
rect 1789 622 1823 1598
rect 2047 622 2081 1598
rect 2305 622 2339 1598
rect 2563 622 2597 1598
rect 2821 622 2855 1598
rect 3079 622 3113 1598
rect -3113 -488 -3079 488
rect -2855 -488 -2821 488
rect -2597 -488 -2563 488
rect -2339 -488 -2305 488
rect -2081 -488 -2047 488
rect -1823 -488 -1789 488
rect -1565 -488 -1531 488
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
rect 1531 -488 1565 488
rect 1789 -488 1823 488
rect 2047 -488 2081 488
rect 2305 -488 2339 488
rect 2563 -488 2597 488
rect 2821 -488 2855 488
rect 3079 -488 3113 488
rect -3113 -1598 -3079 -622
rect -2855 -1598 -2821 -622
rect -2597 -1598 -2563 -622
rect -2339 -1598 -2305 -622
rect -2081 -1598 -2047 -622
rect -1823 -1598 -1789 -622
rect -1565 -1598 -1531 -622
rect -1307 -1598 -1273 -622
rect -1049 -1598 -1015 -622
rect -791 -1598 -757 -622
rect -533 -1598 -499 -622
rect -275 -1598 -241 -622
rect -17 -1598 17 -622
rect 241 -1598 275 -622
rect 499 -1598 533 -622
rect 757 -1598 791 -622
rect 1015 -1598 1049 -622
rect 1273 -1598 1307 -622
rect 1531 -1598 1565 -622
rect 1789 -1598 1823 -622
rect 2047 -1598 2081 -622
rect 2305 -1598 2339 -622
rect 2563 -1598 2597 -622
rect 2821 -1598 2855 -622
rect 3079 -1598 3113 -622
rect -3113 -2708 -3079 -1732
rect -2855 -2708 -2821 -1732
rect -2597 -2708 -2563 -1732
rect -2339 -2708 -2305 -1732
rect -2081 -2708 -2047 -1732
rect -1823 -2708 -1789 -1732
rect -1565 -2708 -1531 -1732
rect -1307 -2708 -1273 -1732
rect -1049 -2708 -1015 -1732
rect -791 -2708 -757 -1732
rect -533 -2708 -499 -1732
rect -275 -2708 -241 -1732
rect -17 -2708 17 -1732
rect 241 -2708 275 -1732
rect 499 -2708 533 -1732
rect 757 -2708 791 -1732
rect 1015 -2708 1049 -1732
rect 1273 -2708 1307 -1732
rect 1531 -2708 1565 -1732
rect 1789 -2708 1823 -1732
rect 2047 -2708 2081 -1732
rect 2305 -2708 2339 -1732
rect 2563 -2708 2597 -1732
rect 2821 -2708 2855 -1732
rect 3079 -2708 3113 -1732
<< mvpsubdiff >>
rect -3259 2930 3259 2942
rect -3259 2896 -3151 2930
rect 3151 2896 3259 2930
rect -3259 2884 3259 2896
rect -3259 2834 -3201 2884
rect -3259 -2834 -3247 2834
rect -3213 -2834 -3201 2834
rect 3201 2834 3259 2884
rect -3259 -2884 -3201 -2834
rect 3201 -2834 3213 2834
rect 3247 -2834 3259 2834
rect 3201 -2884 3259 -2834
rect -3259 -2896 3259 -2884
rect -3259 -2930 -3151 -2896
rect 3151 -2930 3259 -2896
rect -3259 -2942 3259 -2930
<< mvpsubdiffcont >>
rect -3151 2896 3151 2930
rect -3247 -2834 -3213 2834
rect 3213 -2834 3247 2834
rect -3151 -2930 3151 -2896
<< poly >>
rect -3067 2792 -2867 2808
rect -3067 2758 -3051 2792
rect -2883 2758 -2867 2792
rect -3067 2720 -2867 2758
rect -2809 2792 -2609 2808
rect -2809 2758 -2793 2792
rect -2625 2758 -2609 2792
rect -2809 2720 -2609 2758
rect -2551 2792 -2351 2808
rect -2551 2758 -2535 2792
rect -2367 2758 -2351 2792
rect -2551 2720 -2351 2758
rect -2293 2792 -2093 2808
rect -2293 2758 -2277 2792
rect -2109 2758 -2093 2792
rect -2293 2720 -2093 2758
rect -2035 2792 -1835 2808
rect -2035 2758 -2019 2792
rect -1851 2758 -1835 2792
rect -2035 2720 -1835 2758
rect -1777 2792 -1577 2808
rect -1777 2758 -1761 2792
rect -1593 2758 -1577 2792
rect -1777 2720 -1577 2758
rect -1519 2792 -1319 2808
rect -1519 2758 -1503 2792
rect -1335 2758 -1319 2792
rect -1519 2720 -1319 2758
rect -1261 2792 -1061 2808
rect -1261 2758 -1245 2792
rect -1077 2758 -1061 2792
rect -1261 2720 -1061 2758
rect -1003 2792 -803 2808
rect -1003 2758 -987 2792
rect -819 2758 -803 2792
rect -1003 2720 -803 2758
rect -745 2792 -545 2808
rect -745 2758 -729 2792
rect -561 2758 -545 2792
rect -745 2720 -545 2758
rect -487 2792 -287 2808
rect -487 2758 -471 2792
rect -303 2758 -287 2792
rect -487 2720 -287 2758
rect -229 2792 -29 2808
rect -229 2758 -213 2792
rect -45 2758 -29 2792
rect -229 2720 -29 2758
rect 29 2792 229 2808
rect 29 2758 45 2792
rect 213 2758 229 2792
rect 29 2720 229 2758
rect 287 2792 487 2808
rect 287 2758 303 2792
rect 471 2758 487 2792
rect 287 2720 487 2758
rect 545 2792 745 2808
rect 545 2758 561 2792
rect 729 2758 745 2792
rect 545 2720 745 2758
rect 803 2792 1003 2808
rect 803 2758 819 2792
rect 987 2758 1003 2792
rect 803 2720 1003 2758
rect 1061 2792 1261 2808
rect 1061 2758 1077 2792
rect 1245 2758 1261 2792
rect 1061 2720 1261 2758
rect 1319 2792 1519 2808
rect 1319 2758 1335 2792
rect 1503 2758 1519 2792
rect 1319 2720 1519 2758
rect 1577 2792 1777 2808
rect 1577 2758 1593 2792
rect 1761 2758 1777 2792
rect 1577 2720 1777 2758
rect 1835 2792 2035 2808
rect 1835 2758 1851 2792
rect 2019 2758 2035 2792
rect 1835 2720 2035 2758
rect 2093 2792 2293 2808
rect 2093 2758 2109 2792
rect 2277 2758 2293 2792
rect 2093 2720 2293 2758
rect 2351 2792 2551 2808
rect 2351 2758 2367 2792
rect 2535 2758 2551 2792
rect 2351 2720 2551 2758
rect 2609 2792 2809 2808
rect 2609 2758 2625 2792
rect 2793 2758 2809 2792
rect 2609 2720 2809 2758
rect 2867 2792 3067 2808
rect 2867 2758 2883 2792
rect 3051 2758 3067 2792
rect 2867 2720 3067 2758
rect -3067 1682 -2867 1720
rect -3067 1648 -3051 1682
rect -2883 1648 -2867 1682
rect -3067 1610 -2867 1648
rect -2809 1682 -2609 1720
rect -2809 1648 -2793 1682
rect -2625 1648 -2609 1682
rect -2809 1610 -2609 1648
rect -2551 1682 -2351 1720
rect -2551 1648 -2535 1682
rect -2367 1648 -2351 1682
rect -2551 1610 -2351 1648
rect -2293 1682 -2093 1720
rect -2293 1648 -2277 1682
rect -2109 1648 -2093 1682
rect -2293 1610 -2093 1648
rect -2035 1682 -1835 1720
rect -2035 1648 -2019 1682
rect -1851 1648 -1835 1682
rect -2035 1610 -1835 1648
rect -1777 1682 -1577 1720
rect -1777 1648 -1761 1682
rect -1593 1648 -1577 1682
rect -1777 1610 -1577 1648
rect -1519 1682 -1319 1720
rect -1519 1648 -1503 1682
rect -1335 1648 -1319 1682
rect -1519 1610 -1319 1648
rect -1261 1682 -1061 1720
rect -1261 1648 -1245 1682
rect -1077 1648 -1061 1682
rect -1261 1610 -1061 1648
rect -1003 1682 -803 1720
rect -1003 1648 -987 1682
rect -819 1648 -803 1682
rect -1003 1610 -803 1648
rect -745 1682 -545 1720
rect -745 1648 -729 1682
rect -561 1648 -545 1682
rect -745 1610 -545 1648
rect -487 1682 -287 1720
rect -487 1648 -471 1682
rect -303 1648 -287 1682
rect -487 1610 -287 1648
rect -229 1682 -29 1720
rect -229 1648 -213 1682
rect -45 1648 -29 1682
rect -229 1610 -29 1648
rect 29 1682 229 1720
rect 29 1648 45 1682
rect 213 1648 229 1682
rect 29 1610 229 1648
rect 287 1682 487 1720
rect 287 1648 303 1682
rect 471 1648 487 1682
rect 287 1610 487 1648
rect 545 1682 745 1720
rect 545 1648 561 1682
rect 729 1648 745 1682
rect 545 1610 745 1648
rect 803 1682 1003 1720
rect 803 1648 819 1682
rect 987 1648 1003 1682
rect 803 1610 1003 1648
rect 1061 1682 1261 1720
rect 1061 1648 1077 1682
rect 1245 1648 1261 1682
rect 1061 1610 1261 1648
rect 1319 1682 1519 1720
rect 1319 1648 1335 1682
rect 1503 1648 1519 1682
rect 1319 1610 1519 1648
rect 1577 1682 1777 1720
rect 1577 1648 1593 1682
rect 1761 1648 1777 1682
rect 1577 1610 1777 1648
rect 1835 1682 2035 1720
rect 1835 1648 1851 1682
rect 2019 1648 2035 1682
rect 1835 1610 2035 1648
rect 2093 1682 2293 1720
rect 2093 1648 2109 1682
rect 2277 1648 2293 1682
rect 2093 1610 2293 1648
rect 2351 1682 2551 1720
rect 2351 1648 2367 1682
rect 2535 1648 2551 1682
rect 2351 1610 2551 1648
rect 2609 1682 2809 1720
rect 2609 1648 2625 1682
rect 2793 1648 2809 1682
rect 2609 1610 2809 1648
rect 2867 1682 3067 1720
rect 2867 1648 2883 1682
rect 3051 1648 3067 1682
rect 2867 1610 3067 1648
rect -3067 572 -2867 610
rect -3067 538 -3051 572
rect -2883 538 -2867 572
rect -3067 500 -2867 538
rect -2809 572 -2609 610
rect -2809 538 -2793 572
rect -2625 538 -2609 572
rect -2809 500 -2609 538
rect -2551 572 -2351 610
rect -2551 538 -2535 572
rect -2367 538 -2351 572
rect -2551 500 -2351 538
rect -2293 572 -2093 610
rect -2293 538 -2277 572
rect -2109 538 -2093 572
rect -2293 500 -2093 538
rect -2035 572 -1835 610
rect -2035 538 -2019 572
rect -1851 538 -1835 572
rect -2035 500 -1835 538
rect -1777 572 -1577 610
rect -1777 538 -1761 572
rect -1593 538 -1577 572
rect -1777 500 -1577 538
rect -1519 572 -1319 610
rect -1519 538 -1503 572
rect -1335 538 -1319 572
rect -1519 500 -1319 538
rect -1261 572 -1061 610
rect -1261 538 -1245 572
rect -1077 538 -1061 572
rect -1261 500 -1061 538
rect -1003 572 -803 610
rect -1003 538 -987 572
rect -819 538 -803 572
rect -1003 500 -803 538
rect -745 572 -545 610
rect -745 538 -729 572
rect -561 538 -545 572
rect -745 500 -545 538
rect -487 572 -287 610
rect -487 538 -471 572
rect -303 538 -287 572
rect -487 500 -287 538
rect -229 572 -29 610
rect -229 538 -213 572
rect -45 538 -29 572
rect -229 500 -29 538
rect 29 572 229 610
rect 29 538 45 572
rect 213 538 229 572
rect 29 500 229 538
rect 287 572 487 610
rect 287 538 303 572
rect 471 538 487 572
rect 287 500 487 538
rect 545 572 745 610
rect 545 538 561 572
rect 729 538 745 572
rect 545 500 745 538
rect 803 572 1003 610
rect 803 538 819 572
rect 987 538 1003 572
rect 803 500 1003 538
rect 1061 572 1261 610
rect 1061 538 1077 572
rect 1245 538 1261 572
rect 1061 500 1261 538
rect 1319 572 1519 610
rect 1319 538 1335 572
rect 1503 538 1519 572
rect 1319 500 1519 538
rect 1577 572 1777 610
rect 1577 538 1593 572
rect 1761 538 1777 572
rect 1577 500 1777 538
rect 1835 572 2035 610
rect 1835 538 1851 572
rect 2019 538 2035 572
rect 1835 500 2035 538
rect 2093 572 2293 610
rect 2093 538 2109 572
rect 2277 538 2293 572
rect 2093 500 2293 538
rect 2351 572 2551 610
rect 2351 538 2367 572
rect 2535 538 2551 572
rect 2351 500 2551 538
rect 2609 572 2809 610
rect 2609 538 2625 572
rect 2793 538 2809 572
rect 2609 500 2809 538
rect 2867 572 3067 610
rect 2867 538 2883 572
rect 3051 538 3067 572
rect 2867 500 3067 538
rect -3067 -538 -2867 -500
rect -3067 -572 -3051 -538
rect -2883 -572 -2867 -538
rect -3067 -610 -2867 -572
rect -2809 -538 -2609 -500
rect -2809 -572 -2793 -538
rect -2625 -572 -2609 -538
rect -2809 -610 -2609 -572
rect -2551 -538 -2351 -500
rect -2551 -572 -2535 -538
rect -2367 -572 -2351 -538
rect -2551 -610 -2351 -572
rect -2293 -538 -2093 -500
rect -2293 -572 -2277 -538
rect -2109 -572 -2093 -538
rect -2293 -610 -2093 -572
rect -2035 -538 -1835 -500
rect -2035 -572 -2019 -538
rect -1851 -572 -1835 -538
rect -2035 -610 -1835 -572
rect -1777 -538 -1577 -500
rect -1777 -572 -1761 -538
rect -1593 -572 -1577 -538
rect -1777 -610 -1577 -572
rect -1519 -538 -1319 -500
rect -1519 -572 -1503 -538
rect -1335 -572 -1319 -538
rect -1519 -610 -1319 -572
rect -1261 -538 -1061 -500
rect -1261 -572 -1245 -538
rect -1077 -572 -1061 -538
rect -1261 -610 -1061 -572
rect -1003 -538 -803 -500
rect -1003 -572 -987 -538
rect -819 -572 -803 -538
rect -1003 -610 -803 -572
rect -745 -538 -545 -500
rect -745 -572 -729 -538
rect -561 -572 -545 -538
rect -745 -610 -545 -572
rect -487 -538 -287 -500
rect -487 -572 -471 -538
rect -303 -572 -287 -538
rect -487 -610 -287 -572
rect -229 -538 -29 -500
rect -229 -572 -213 -538
rect -45 -572 -29 -538
rect -229 -610 -29 -572
rect 29 -538 229 -500
rect 29 -572 45 -538
rect 213 -572 229 -538
rect 29 -610 229 -572
rect 287 -538 487 -500
rect 287 -572 303 -538
rect 471 -572 487 -538
rect 287 -610 487 -572
rect 545 -538 745 -500
rect 545 -572 561 -538
rect 729 -572 745 -538
rect 545 -610 745 -572
rect 803 -538 1003 -500
rect 803 -572 819 -538
rect 987 -572 1003 -538
rect 803 -610 1003 -572
rect 1061 -538 1261 -500
rect 1061 -572 1077 -538
rect 1245 -572 1261 -538
rect 1061 -610 1261 -572
rect 1319 -538 1519 -500
rect 1319 -572 1335 -538
rect 1503 -572 1519 -538
rect 1319 -610 1519 -572
rect 1577 -538 1777 -500
rect 1577 -572 1593 -538
rect 1761 -572 1777 -538
rect 1577 -610 1777 -572
rect 1835 -538 2035 -500
rect 1835 -572 1851 -538
rect 2019 -572 2035 -538
rect 1835 -610 2035 -572
rect 2093 -538 2293 -500
rect 2093 -572 2109 -538
rect 2277 -572 2293 -538
rect 2093 -610 2293 -572
rect 2351 -538 2551 -500
rect 2351 -572 2367 -538
rect 2535 -572 2551 -538
rect 2351 -610 2551 -572
rect 2609 -538 2809 -500
rect 2609 -572 2625 -538
rect 2793 -572 2809 -538
rect 2609 -610 2809 -572
rect 2867 -538 3067 -500
rect 2867 -572 2883 -538
rect 3051 -572 3067 -538
rect 2867 -610 3067 -572
rect -3067 -1648 -2867 -1610
rect -3067 -1682 -3051 -1648
rect -2883 -1682 -2867 -1648
rect -3067 -1720 -2867 -1682
rect -2809 -1648 -2609 -1610
rect -2809 -1682 -2793 -1648
rect -2625 -1682 -2609 -1648
rect -2809 -1720 -2609 -1682
rect -2551 -1648 -2351 -1610
rect -2551 -1682 -2535 -1648
rect -2367 -1682 -2351 -1648
rect -2551 -1720 -2351 -1682
rect -2293 -1648 -2093 -1610
rect -2293 -1682 -2277 -1648
rect -2109 -1682 -2093 -1648
rect -2293 -1720 -2093 -1682
rect -2035 -1648 -1835 -1610
rect -2035 -1682 -2019 -1648
rect -1851 -1682 -1835 -1648
rect -2035 -1720 -1835 -1682
rect -1777 -1648 -1577 -1610
rect -1777 -1682 -1761 -1648
rect -1593 -1682 -1577 -1648
rect -1777 -1720 -1577 -1682
rect -1519 -1648 -1319 -1610
rect -1519 -1682 -1503 -1648
rect -1335 -1682 -1319 -1648
rect -1519 -1720 -1319 -1682
rect -1261 -1648 -1061 -1610
rect -1261 -1682 -1245 -1648
rect -1077 -1682 -1061 -1648
rect -1261 -1720 -1061 -1682
rect -1003 -1648 -803 -1610
rect -1003 -1682 -987 -1648
rect -819 -1682 -803 -1648
rect -1003 -1720 -803 -1682
rect -745 -1648 -545 -1610
rect -745 -1682 -729 -1648
rect -561 -1682 -545 -1648
rect -745 -1720 -545 -1682
rect -487 -1648 -287 -1610
rect -487 -1682 -471 -1648
rect -303 -1682 -287 -1648
rect -487 -1720 -287 -1682
rect -229 -1648 -29 -1610
rect -229 -1682 -213 -1648
rect -45 -1682 -29 -1648
rect -229 -1720 -29 -1682
rect 29 -1648 229 -1610
rect 29 -1682 45 -1648
rect 213 -1682 229 -1648
rect 29 -1720 229 -1682
rect 287 -1648 487 -1610
rect 287 -1682 303 -1648
rect 471 -1682 487 -1648
rect 287 -1720 487 -1682
rect 545 -1648 745 -1610
rect 545 -1682 561 -1648
rect 729 -1682 745 -1648
rect 545 -1720 745 -1682
rect 803 -1648 1003 -1610
rect 803 -1682 819 -1648
rect 987 -1682 1003 -1648
rect 803 -1720 1003 -1682
rect 1061 -1648 1261 -1610
rect 1061 -1682 1077 -1648
rect 1245 -1682 1261 -1648
rect 1061 -1720 1261 -1682
rect 1319 -1648 1519 -1610
rect 1319 -1682 1335 -1648
rect 1503 -1682 1519 -1648
rect 1319 -1720 1519 -1682
rect 1577 -1648 1777 -1610
rect 1577 -1682 1593 -1648
rect 1761 -1682 1777 -1648
rect 1577 -1720 1777 -1682
rect 1835 -1648 2035 -1610
rect 1835 -1682 1851 -1648
rect 2019 -1682 2035 -1648
rect 1835 -1720 2035 -1682
rect 2093 -1648 2293 -1610
rect 2093 -1682 2109 -1648
rect 2277 -1682 2293 -1648
rect 2093 -1720 2293 -1682
rect 2351 -1648 2551 -1610
rect 2351 -1682 2367 -1648
rect 2535 -1682 2551 -1648
rect 2351 -1720 2551 -1682
rect 2609 -1648 2809 -1610
rect 2609 -1682 2625 -1648
rect 2793 -1682 2809 -1648
rect 2609 -1720 2809 -1682
rect 2867 -1648 3067 -1610
rect 2867 -1682 2883 -1648
rect 3051 -1682 3067 -1648
rect 2867 -1720 3067 -1682
rect -3067 -2758 -2867 -2720
rect -3067 -2792 -3051 -2758
rect -2883 -2792 -2867 -2758
rect -3067 -2808 -2867 -2792
rect -2809 -2758 -2609 -2720
rect -2809 -2792 -2793 -2758
rect -2625 -2792 -2609 -2758
rect -2809 -2808 -2609 -2792
rect -2551 -2758 -2351 -2720
rect -2551 -2792 -2535 -2758
rect -2367 -2792 -2351 -2758
rect -2551 -2808 -2351 -2792
rect -2293 -2758 -2093 -2720
rect -2293 -2792 -2277 -2758
rect -2109 -2792 -2093 -2758
rect -2293 -2808 -2093 -2792
rect -2035 -2758 -1835 -2720
rect -2035 -2792 -2019 -2758
rect -1851 -2792 -1835 -2758
rect -2035 -2808 -1835 -2792
rect -1777 -2758 -1577 -2720
rect -1777 -2792 -1761 -2758
rect -1593 -2792 -1577 -2758
rect -1777 -2808 -1577 -2792
rect -1519 -2758 -1319 -2720
rect -1519 -2792 -1503 -2758
rect -1335 -2792 -1319 -2758
rect -1519 -2808 -1319 -2792
rect -1261 -2758 -1061 -2720
rect -1261 -2792 -1245 -2758
rect -1077 -2792 -1061 -2758
rect -1261 -2808 -1061 -2792
rect -1003 -2758 -803 -2720
rect -1003 -2792 -987 -2758
rect -819 -2792 -803 -2758
rect -1003 -2808 -803 -2792
rect -745 -2758 -545 -2720
rect -745 -2792 -729 -2758
rect -561 -2792 -545 -2758
rect -745 -2808 -545 -2792
rect -487 -2758 -287 -2720
rect -487 -2792 -471 -2758
rect -303 -2792 -287 -2758
rect -487 -2808 -287 -2792
rect -229 -2758 -29 -2720
rect -229 -2792 -213 -2758
rect -45 -2792 -29 -2758
rect -229 -2808 -29 -2792
rect 29 -2758 229 -2720
rect 29 -2792 45 -2758
rect 213 -2792 229 -2758
rect 29 -2808 229 -2792
rect 287 -2758 487 -2720
rect 287 -2792 303 -2758
rect 471 -2792 487 -2758
rect 287 -2808 487 -2792
rect 545 -2758 745 -2720
rect 545 -2792 561 -2758
rect 729 -2792 745 -2758
rect 545 -2808 745 -2792
rect 803 -2758 1003 -2720
rect 803 -2792 819 -2758
rect 987 -2792 1003 -2758
rect 803 -2808 1003 -2792
rect 1061 -2758 1261 -2720
rect 1061 -2792 1077 -2758
rect 1245 -2792 1261 -2758
rect 1061 -2808 1261 -2792
rect 1319 -2758 1519 -2720
rect 1319 -2792 1335 -2758
rect 1503 -2792 1519 -2758
rect 1319 -2808 1519 -2792
rect 1577 -2758 1777 -2720
rect 1577 -2792 1593 -2758
rect 1761 -2792 1777 -2758
rect 1577 -2808 1777 -2792
rect 1835 -2758 2035 -2720
rect 1835 -2792 1851 -2758
rect 2019 -2792 2035 -2758
rect 1835 -2808 2035 -2792
rect 2093 -2758 2293 -2720
rect 2093 -2792 2109 -2758
rect 2277 -2792 2293 -2758
rect 2093 -2808 2293 -2792
rect 2351 -2758 2551 -2720
rect 2351 -2792 2367 -2758
rect 2535 -2792 2551 -2758
rect 2351 -2808 2551 -2792
rect 2609 -2758 2809 -2720
rect 2609 -2792 2625 -2758
rect 2793 -2792 2809 -2758
rect 2609 -2808 2809 -2792
rect 2867 -2758 3067 -2720
rect 2867 -2792 2883 -2758
rect 3051 -2792 3067 -2758
rect 2867 -2808 3067 -2792
<< polycont >>
rect -3051 2758 -2883 2792
rect -2793 2758 -2625 2792
rect -2535 2758 -2367 2792
rect -2277 2758 -2109 2792
rect -2019 2758 -1851 2792
rect -1761 2758 -1593 2792
rect -1503 2758 -1335 2792
rect -1245 2758 -1077 2792
rect -987 2758 -819 2792
rect -729 2758 -561 2792
rect -471 2758 -303 2792
rect -213 2758 -45 2792
rect 45 2758 213 2792
rect 303 2758 471 2792
rect 561 2758 729 2792
rect 819 2758 987 2792
rect 1077 2758 1245 2792
rect 1335 2758 1503 2792
rect 1593 2758 1761 2792
rect 1851 2758 2019 2792
rect 2109 2758 2277 2792
rect 2367 2758 2535 2792
rect 2625 2758 2793 2792
rect 2883 2758 3051 2792
rect -3051 1648 -2883 1682
rect -2793 1648 -2625 1682
rect -2535 1648 -2367 1682
rect -2277 1648 -2109 1682
rect -2019 1648 -1851 1682
rect -1761 1648 -1593 1682
rect -1503 1648 -1335 1682
rect -1245 1648 -1077 1682
rect -987 1648 -819 1682
rect -729 1648 -561 1682
rect -471 1648 -303 1682
rect -213 1648 -45 1682
rect 45 1648 213 1682
rect 303 1648 471 1682
rect 561 1648 729 1682
rect 819 1648 987 1682
rect 1077 1648 1245 1682
rect 1335 1648 1503 1682
rect 1593 1648 1761 1682
rect 1851 1648 2019 1682
rect 2109 1648 2277 1682
rect 2367 1648 2535 1682
rect 2625 1648 2793 1682
rect 2883 1648 3051 1682
rect -3051 538 -2883 572
rect -2793 538 -2625 572
rect -2535 538 -2367 572
rect -2277 538 -2109 572
rect -2019 538 -1851 572
rect -1761 538 -1593 572
rect -1503 538 -1335 572
rect -1245 538 -1077 572
rect -987 538 -819 572
rect -729 538 -561 572
rect -471 538 -303 572
rect -213 538 -45 572
rect 45 538 213 572
rect 303 538 471 572
rect 561 538 729 572
rect 819 538 987 572
rect 1077 538 1245 572
rect 1335 538 1503 572
rect 1593 538 1761 572
rect 1851 538 2019 572
rect 2109 538 2277 572
rect 2367 538 2535 572
rect 2625 538 2793 572
rect 2883 538 3051 572
rect -3051 -572 -2883 -538
rect -2793 -572 -2625 -538
rect -2535 -572 -2367 -538
rect -2277 -572 -2109 -538
rect -2019 -572 -1851 -538
rect -1761 -572 -1593 -538
rect -1503 -572 -1335 -538
rect -1245 -572 -1077 -538
rect -987 -572 -819 -538
rect -729 -572 -561 -538
rect -471 -572 -303 -538
rect -213 -572 -45 -538
rect 45 -572 213 -538
rect 303 -572 471 -538
rect 561 -572 729 -538
rect 819 -572 987 -538
rect 1077 -572 1245 -538
rect 1335 -572 1503 -538
rect 1593 -572 1761 -538
rect 1851 -572 2019 -538
rect 2109 -572 2277 -538
rect 2367 -572 2535 -538
rect 2625 -572 2793 -538
rect 2883 -572 3051 -538
rect -3051 -1682 -2883 -1648
rect -2793 -1682 -2625 -1648
rect -2535 -1682 -2367 -1648
rect -2277 -1682 -2109 -1648
rect -2019 -1682 -1851 -1648
rect -1761 -1682 -1593 -1648
rect -1503 -1682 -1335 -1648
rect -1245 -1682 -1077 -1648
rect -987 -1682 -819 -1648
rect -729 -1682 -561 -1648
rect -471 -1682 -303 -1648
rect -213 -1682 -45 -1648
rect 45 -1682 213 -1648
rect 303 -1682 471 -1648
rect 561 -1682 729 -1648
rect 819 -1682 987 -1648
rect 1077 -1682 1245 -1648
rect 1335 -1682 1503 -1648
rect 1593 -1682 1761 -1648
rect 1851 -1682 2019 -1648
rect 2109 -1682 2277 -1648
rect 2367 -1682 2535 -1648
rect 2625 -1682 2793 -1648
rect 2883 -1682 3051 -1648
rect -3051 -2792 -2883 -2758
rect -2793 -2792 -2625 -2758
rect -2535 -2792 -2367 -2758
rect -2277 -2792 -2109 -2758
rect -2019 -2792 -1851 -2758
rect -1761 -2792 -1593 -2758
rect -1503 -2792 -1335 -2758
rect -1245 -2792 -1077 -2758
rect -987 -2792 -819 -2758
rect -729 -2792 -561 -2758
rect -471 -2792 -303 -2758
rect -213 -2792 -45 -2758
rect 45 -2792 213 -2758
rect 303 -2792 471 -2758
rect 561 -2792 729 -2758
rect 819 -2792 987 -2758
rect 1077 -2792 1245 -2758
rect 1335 -2792 1503 -2758
rect 1593 -2792 1761 -2758
rect 1851 -2792 2019 -2758
rect 2109 -2792 2277 -2758
rect 2367 -2792 2535 -2758
rect 2625 -2792 2793 -2758
rect 2883 -2792 3051 -2758
<< locali >>
rect -3247 2896 -3151 2930
rect 3151 2896 3247 2930
rect -3247 2834 -3213 2896
rect 3213 2834 3247 2896
rect -3067 2758 -3051 2792
rect -2883 2758 -2867 2792
rect -2809 2758 -2793 2792
rect -2625 2758 -2609 2792
rect -2551 2758 -2535 2792
rect -2367 2758 -2351 2792
rect -2293 2758 -2277 2792
rect -2109 2758 -2093 2792
rect -2035 2758 -2019 2792
rect -1851 2758 -1835 2792
rect -1777 2758 -1761 2792
rect -1593 2758 -1577 2792
rect -1519 2758 -1503 2792
rect -1335 2758 -1319 2792
rect -1261 2758 -1245 2792
rect -1077 2758 -1061 2792
rect -1003 2758 -987 2792
rect -819 2758 -803 2792
rect -745 2758 -729 2792
rect -561 2758 -545 2792
rect -487 2758 -471 2792
rect -303 2758 -287 2792
rect -229 2758 -213 2792
rect -45 2758 -29 2792
rect 29 2758 45 2792
rect 213 2758 229 2792
rect 287 2758 303 2792
rect 471 2758 487 2792
rect 545 2758 561 2792
rect 729 2758 745 2792
rect 803 2758 819 2792
rect 987 2758 1003 2792
rect 1061 2758 1077 2792
rect 1245 2758 1261 2792
rect 1319 2758 1335 2792
rect 1503 2758 1519 2792
rect 1577 2758 1593 2792
rect 1761 2758 1777 2792
rect 1835 2758 1851 2792
rect 2019 2758 2035 2792
rect 2093 2758 2109 2792
rect 2277 2758 2293 2792
rect 2351 2758 2367 2792
rect 2535 2758 2551 2792
rect 2609 2758 2625 2792
rect 2793 2758 2809 2792
rect 2867 2758 2883 2792
rect 3051 2758 3067 2792
rect -3113 2708 -3079 2724
rect -3113 1716 -3079 1732
rect -2855 2708 -2821 2724
rect -2855 1716 -2821 1732
rect -2597 2708 -2563 2724
rect -2597 1716 -2563 1732
rect -2339 2708 -2305 2724
rect -2339 1716 -2305 1732
rect -2081 2708 -2047 2724
rect -2081 1716 -2047 1732
rect -1823 2708 -1789 2724
rect -1823 1716 -1789 1732
rect -1565 2708 -1531 2724
rect -1565 1716 -1531 1732
rect -1307 2708 -1273 2724
rect -1307 1716 -1273 1732
rect -1049 2708 -1015 2724
rect -1049 1716 -1015 1732
rect -791 2708 -757 2724
rect -791 1716 -757 1732
rect -533 2708 -499 2724
rect -533 1716 -499 1732
rect -275 2708 -241 2724
rect -275 1716 -241 1732
rect -17 2708 17 2724
rect -17 1716 17 1732
rect 241 2708 275 2724
rect 241 1716 275 1732
rect 499 2708 533 2724
rect 499 1716 533 1732
rect 757 2708 791 2724
rect 757 1716 791 1732
rect 1015 2708 1049 2724
rect 1015 1716 1049 1732
rect 1273 2708 1307 2724
rect 1273 1716 1307 1732
rect 1531 2708 1565 2724
rect 1531 1716 1565 1732
rect 1789 2708 1823 2724
rect 1789 1716 1823 1732
rect 2047 2708 2081 2724
rect 2047 1716 2081 1732
rect 2305 2708 2339 2724
rect 2305 1716 2339 1732
rect 2563 2708 2597 2724
rect 2563 1716 2597 1732
rect 2821 2708 2855 2724
rect 2821 1716 2855 1732
rect 3079 2708 3113 2724
rect 3079 1716 3113 1732
rect -3067 1648 -3051 1682
rect -2883 1648 -2867 1682
rect -2809 1648 -2793 1682
rect -2625 1648 -2609 1682
rect -2551 1648 -2535 1682
rect -2367 1648 -2351 1682
rect -2293 1648 -2277 1682
rect -2109 1648 -2093 1682
rect -2035 1648 -2019 1682
rect -1851 1648 -1835 1682
rect -1777 1648 -1761 1682
rect -1593 1648 -1577 1682
rect -1519 1648 -1503 1682
rect -1335 1648 -1319 1682
rect -1261 1648 -1245 1682
rect -1077 1648 -1061 1682
rect -1003 1648 -987 1682
rect -819 1648 -803 1682
rect -745 1648 -729 1682
rect -561 1648 -545 1682
rect -487 1648 -471 1682
rect -303 1648 -287 1682
rect -229 1648 -213 1682
rect -45 1648 -29 1682
rect 29 1648 45 1682
rect 213 1648 229 1682
rect 287 1648 303 1682
rect 471 1648 487 1682
rect 545 1648 561 1682
rect 729 1648 745 1682
rect 803 1648 819 1682
rect 987 1648 1003 1682
rect 1061 1648 1077 1682
rect 1245 1648 1261 1682
rect 1319 1648 1335 1682
rect 1503 1648 1519 1682
rect 1577 1648 1593 1682
rect 1761 1648 1777 1682
rect 1835 1648 1851 1682
rect 2019 1648 2035 1682
rect 2093 1648 2109 1682
rect 2277 1648 2293 1682
rect 2351 1648 2367 1682
rect 2535 1648 2551 1682
rect 2609 1648 2625 1682
rect 2793 1648 2809 1682
rect 2867 1648 2883 1682
rect 3051 1648 3067 1682
rect -3113 1598 -3079 1614
rect -3113 606 -3079 622
rect -2855 1598 -2821 1614
rect -2855 606 -2821 622
rect -2597 1598 -2563 1614
rect -2597 606 -2563 622
rect -2339 1598 -2305 1614
rect -2339 606 -2305 622
rect -2081 1598 -2047 1614
rect -2081 606 -2047 622
rect -1823 1598 -1789 1614
rect -1823 606 -1789 622
rect -1565 1598 -1531 1614
rect -1565 606 -1531 622
rect -1307 1598 -1273 1614
rect -1307 606 -1273 622
rect -1049 1598 -1015 1614
rect -1049 606 -1015 622
rect -791 1598 -757 1614
rect -791 606 -757 622
rect -533 1598 -499 1614
rect -533 606 -499 622
rect -275 1598 -241 1614
rect -275 606 -241 622
rect -17 1598 17 1614
rect -17 606 17 622
rect 241 1598 275 1614
rect 241 606 275 622
rect 499 1598 533 1614
rect 499 606 533 622
rect 757 1598 791 1614
rect 757 606 791 622
rect 1015 1598 1049 1614
rect 1015 606 1049 622
rect 1273 1598 1307 1614
rect 1273 606 1307 622
rect 1531 1598 1565 1614
rect 1531 606 1565 622
rect 1789 1598 1823 1614
rect 1789 606 1823 622
rect 2047 1598 2081 1614
rect 2047 606 2081 622
rect 2305 1598 2339 1614
rect 2305 606 2339 622
rect 2563 1598 2597 1614
rect 2563 606 2597 622
rect 2821 1598 2855 1614
rect 2821 606 2855 622
rect 3079 1598 3113 1614
rect 3079 606 3113 622
rect -3067 538 -3051 572
rect -2883 538 -2867 572
rect -2809 538 -2793 572
rect -2625 538 -2609 572
rect -2551 538 -2535 572
rect -2367 538 -2351 572
rect -2293 538 -2277 572
rect -2109 538 -2093 572
rect -2035 538 -2019 572
rect -1851 538 -1835 572
rect -1777 538 -1761 572
rect -1593 538 -1577 572
rect -1519 538 -1503 572
rect -1335 538 -1319 572
rect -1261 538 -1245 572
rect -1077 538 -1061 572
rect -1003 538 -987 572
rect -819 538 -803 572
rect -745 538 -729 572
rect -561 538 -545 572
rect -487 538 -471 572
rect -303 538 -287 572
rect -229 538 -213 572
rect -45 538 -29 572
rect 29 538 45 572
rect 213 538 229 572
rect 287 538 303 572
rect 471 538 487 572
rect 545 538 561 572
rect 729 538 745 572
rect 803 538 819 572
rect 987 538 1003 572
rect 1061 538 1077 572
rect 1245 538 1261 572
rect 1319 538 1335 572
rect 1503 538 1519 572
rect 1577 538 1593 572
rect 1761 538 1777 572
rect 1835 538 1851 572
rect 2019 538 2035 572
rect 2093 538 2109 572
rect 2277 538 2293 572
rect 2351 538 2367 572
rect 2535 538 2551 572
rect 2609 538 2625 572
rect 2793 538 2809 572
rect 2867 538 2883 572
rect 3051 538 3067 572
rect -3113 488 -3079 504
rect -3113 -504 -3079 -488
rect -2855 488 -2821 504
rect -2855 -504 -2821 -488
rect -2597 488 -2563 504
rect -2597 -504 -2563 -488
rect -2339 488 -2305 504
rect -2339 -504 -2305 -488
rect -2081 488 -2047 504
rect -2081 -504 -2047 -488
rect -1823 488 -1789 504
rect -1823 -504 -1789 -488
rect -1565 488 -1531 504
rect -1565 -504 -1531 -488
rect -1307 488 -1273 504
rect -1307 -504 -1273 -488
rect -1049 488 -1015 504
rect -1049 -504 -1015 -488
rect -791 488 -757 504
rect -791 -504 -757 -488
rect -533 488 -499 504
rect -533 -504 -499 -488
rect -275 488 -241 504
rect -275 -504 -241 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 241 488 275 504
rect 241 -504 275 -488
rect 499 488 533 504
rect 499 -504 533 -488
rect 757 488 791 504
rect 757 -504 791 -488
rect 1015 488 1049 504
rect 1015 -504 1049 -488
rect 1273 488 1307 504
rect 1273 -504 1307 -488
rect 1531 488 1565 504
rect 1531 -504 1565 -488
rect 1789 488 1823 504
rect 1789 -504 1823 -488
rect 2047 488 2081 504
rect 2047 -504 2081 -488
rect 2305 488 2339 504
rect 2305 -504 2339 -488
rect 2563 488 2597 504
rect 2563 -504 2597 -488
rect 2821 488 2855 504
rect 2821 -504 2855 -488
rect 3079 488 3113 504
rect 3079 -504 3113 -488
rect -3067 -572 -3051 -538
rect -2883 -572 -2867 -538
rect -2809 -572 -2793 -538
rect -2625 -572 -2609 -538
rect -2551 -572 -2535 -538
rect -2367 -572 -2351 -538
rect -2293 -572 -2277 -538
rect -2109 -572 -2093 -538
rect -2035 -572 -2019 -538
rect -1851 -572 -1835 -538
rect -1777 -572 -1761 -538
rect -1593 -572 -1577 -538
rect -1519 -572 -1503 -538
rect -1335 -572 -1319 -538
rect -1261 -572 -1245 -538
rect -1077 -572 -1061 -538
rect -1003 -572 -987 -538
rect -819 -572 -803 -538
rect -745 -572 -729 -538
rect -561 -572 -545 -538
rect -487 -572 -471 -538
rect -303 -572 -287 -538
rect -229 -572 -213 -538
rect -45 -572 -29 -538
rect 29 -572 45 -538
rect 213 -572 229 -538
rect 287 -572 303 -538
rect 471 -572 487 -538
rect 545 -572 561 -538
rect 729 -572 745 -538
rect 803 -572 819 -538
rect 987 -572 1003 -538
rect 1061 -572 1077 -538
rect 1245 -572 1261 -538
rect 1319 -572 1335 -538
rect 1503 -572 1519 -538
rect 1577 -572 1593 -538
rect 1761 -572 1777 -538
rect 1835 -572 1851 -538
rect 2019 -572 2035 -538
rect 2093 -572 2109 -538
rect 2277 -572 2293 -538
rect 2351 -572 2367 -538
rect 2535 -572 2551 -538
rect 2609 -572 2625 -538
rect 2793 -572 2809 -538
rect 2867 -572 2883 -538
rect 3051 -572 3067 -538
rect -3113 -622 -3079 -606
rect -3113 -1614 -3079 -1598
rect -2855 -622 -2821 -606
rect -2855 -1614 -2821 -1598
rect -2597 -622 -2563 -606
rect -2597 -1614 -2563 -1598
rect -2339 -622 -2305 -606
rect -2339 -1614 -2305 -1598
rect -2081 -622 -2047 -606
rect -2081 -1614 -2047 -1598
rect -1823 -622 -1789 -606
rect -1823 -1614 -1789 -1598
rect -1565 -622 -1531 -606
rect -1565 -1614 -1531 -1598
rect -1307 -622 -1273 -606
rect -1307 -1614 -1273 -1598
rect -1049 -622 -1015 -606
rect -1049 -1614 -1015 -1598
rect -791 -622 -757 -606
rect -791 -1614 -757 -1598
rect -533 -622 -499 -606
rect -533 -1614 -499 -1598
rect -275 -622 -241 -606
rect -275 -1614 -241 -1598
rect -17 -622 17 -606
rect -17 -1614 17 -1598
rect 241 -622 275 -606
rect 241 -1614 275 -1598
rect 499 -622 533 -606
rect 499 -1614 533 -1598
rect 757 -622 791 -606
rect 757 -1614 791 -1598
rect 1015 -622 1049 -606
rect 1015 -1614 1049 -1598
rect 1273 -622 1307 -606
rect 1273 -1614 1307 -1598
rect 1531 -622 1565 -606
rect 1531 -1614 1565 -1598
rect 1789 -622 1823 -606
rect 1789 -1614 1823 -1598
rect 2047 -622 2081 -606
rect 2047 -1614 2081 -1598
rect 2305 -622 2339 -606
rect 2305 -1614 2339 -1598
rect 2563 -622 2597 -606
rect 2563 -1614 2597 -1598
rect 2821 -622 2855 -606
rect 2821 -1614 2855 -1598
rect 3079 -622 3113 -606
rect 3079 -1614 3113 -1598
rect -3067 -1682 -3051 -1648
rect -2883 -1682 -2867 -1648
rect -2809 -1682 -2793 -1648
rect -2625 -1682 -2609 -1648
rect -2551 -1682 -2535 -1648
rect -2367 -1682 -2351 -1648
rect -2293 -1682 -2277 -1648
rect -2109 -1682 -2093 -1648
rect -2035 -1682 -2019 -1648
rect -1851 -1682 -1835 -1648
rect -1777 -1682 -1761 -1648
rect -1593 -1682 -1577 -1648
rect -1519 -1682 -1503 -1648
rect -1335 -1682 -1319 -1648
rect -1261 -1682 -1245 -1648
rect -1077 -1682 -1061 -1648
rect -1003 -1682 -987 -1648
rect -819 -1682 -803 -1648
rect -745 -1682 -729 -1648
rect -561 -1682 -545 -1648
rect -487 -1682 -471 -1648
rect -303 -1682 -287 -1648
rect -229 -1682 -213 -1648
rect -45 -1682 -29 -1648
rect 29 -1682 45 -1648
rect 213 -1682 229 -1648
rect 287 -1682 303 -1648
rect 471 -1682 487 -1648
rect 545 -1682 561 -1648
rect 729 -1682 745 -1648
rect 803 -1682 819 -1648
rect 987 -1682 1003 -1648
rect 1061 -1682 1077 -1648
rect 1245 -1682 1261 -1648
rect 1319 -1682 1335 -1648
rect 1503 -1682 1519 -1648
rect 1577 -1682 1593 -1648
rect 1761 -1682 1777 -1648
rect 1835 -1682 1851 -1648
rect 2019 -1682 2035 -1648
rect 2093 -1682 2109 -1648
rect 2277 -1682 2293 -1648
rect 2351 -1682 2367 -1648
rect 2535 -1682 2551 -1648
rect 2609 -1682 2625 -1648
rect 2793 -1682 2809 -1648
rect 2867 -1682 2883 -1648
rect 3051 -1682 3067 -1648
rect -3113 -1732 -3079 -1716
rect -3113 -2724 -3079 -2708
rect -2855 -1732 -2821 -1716
rect -2855 -2724 -2821 -2708
rect -2597 -1732 -2563 -1716
rect -2597 -2724 -2563 -2708
rect -2339 -1732 -2305 -1716
rect -2339 -2724 -2305 -2708
rect -2081 -1732 -2047 -1716
rect -2081 -2724 -2047 -2708
rect -1823 -1732 -1789 -1716
rect -1823 -2724 -1789 -2708
rect -1565 -1732 -1531 -1716
rect -1565 -2724 -1531 -2708
rect -1307 -1732 -1273 -1716
rect -1307 -2724 -1273 -2708
rect -1049 -1732 -1015 -1716
rect -1049 -2724 -1015 -2708
rect -791 -1732 -757 -1716
rect -791 -2724 -757 -2708
rect -533 -1732 -499 -1716
rect -533 -2724 -499 -2708
rect -275 -1732 -241 -1716
rect -275 -2724 -241 -2708
rect -17 -1732 17 -1716
rect -17 -2724 17 -2708
rect 241 -1732 275 -1716
rect 241 -2724 275 -2708
rect 499 -1732 533 -1716
rect 499 -2724 533 -2708
rect 757 -1732 791 -1716
rect 757 -2724 791 -2708
rect 1015 -1732 1049 -1716
rect 1015 -2724 1049 -2708
rect 1273 -1732 1307 -1716
rect 1273 -2724 1307 -2708
rect 1531 -1732 1565 -1716
rect 1531 -2724 1565 -2708
rect 1789 -1732 1823 -1716
rect 1789 -2724 1823 -2708
rect 2047 -1732 2081 -1716
rect 2047 -2724 2081 -2708
rect 2305 -1732 2339 -1716
rect 2305 -2724 2339 -2708
rect 2563 -1732 2597 -1716
rect 2563 -2724 2597 -2708
rect 2821 -1732 2855 -1716
rect 2821 -2724 2855 -2708
rect 3079 -1732 3113 -1716
rect 3079 -2724 3113 -2708
rect -3067 -2792 -3051 -2758
rect -2883 -2792 -2867 -2758
rect -2809 -2792 -2793 -2758
rect -2625 -2792 -2609 -2758
rect -2551 -2792 -2535 -2758
rect -2367 -2792 -2351 -2758
rect -2293 -2792 -2277 -2758
rect -2109 -2792 -2093 -2758
rect -2035 -2792 -2019 -2758
rect -1851 -2792 -1835 -2758
rect -1777 -2792 -1761 -2758
rect -1593 -2792 -1577 -2758
rect -1519 -2792 -1503 -2758
rect -1335 -2792 -1319 -2758
rect -1261 -2792 -1245 -2758
rect -1077 -2792 -1061 -2758
rect -1003 -2792 -987 -2758
rect -819 -2792 -803 -2758
rect -745 -2792 -729 -2758
rect -561 -2792 -545 -2758
rect -487 -2792 -471 -2758
rect -303 -2792 -287 -2758
rect -229 -2792 -213 -2758
rect -45 -2792 -29 -2758
rect 29 -2792 45 -2758
rect 213 -2792 229 -2758
rect 287 -2792 303 -2758
rect 471 -2792 487 -2758
rect 545 -2792 561 -2758
rect 729 -2792 745 -2758
rect 803 -2792 819 -2758
rect 987 -2792 1003 -2758
rect 1061 -2792 1077 -2758
rect 1245 -2792 1261 -2758
rect 1319 -2792 1335 -2758
rect 1503 -2792 1519 -2758
rect 1577 -2792 1593 -2758
rect 1761 -2792 1777 -2758
rect 1835 -2792 1851 -2758
rect 2019 -2792 2035 -2758
rect 2093 -2792 2109 -2758
rect 2277 -2792 2293 -2758
rect 2351 -2792 2367 -2758
rect 2535 -2792 2551 -2758
rect 2609 -2792 2625 -2758
rect 2793 -2792 2809 -2758
rect 2867 -2792 2883 -2758
rect 3051 -2792 3067 -2758
rect -3247 -2896 -3213 -2834
rect 3213 -2896 3247 -2834
rect -3247 -2930 -3151 -2896
rect 3151 -2930 3247 -2896
<< viali >>
rect -3051 2758 -2883 2792
rect -2793 2758 -2625 2792
rect -2535 2758 -2367 2792
rect -2277 2758 -2109 2792
rect -2019 2758 -1851 2792
rect -1761 2758 -1593 2792
rect -1503 2758 -1335 2792
rect -1245 2758 -1077 2792
rect -987 2758 -819 2792
rect -729 2758 -561 2792
rect -471 2758 -303 2792
rect -213 2758 -45 2792
rect 45 2758 213 2792
rect 303 2758 471 2792
rect 561 2758 729 2792
rect 819 2758 987 2792
rect 1077 2758 1245 2792
rect 1335 2758 1503 2792
rect 1593 2758 1761 2792
rect 1851 2758 2019 2792
rect 2109 2758 2277 2792
rect 2367 2758 2535 2792
rect 2625 2758 2793 2792
rect 2883 2758 3051 2792
rect -3113 1732 -3079 2708
rect -2855 1732 -2821 2708
rect -2597 1732 -2563 2708
rect -2339 1732 -2305 2708
rect -2081 1732 -2047 2708
rect -1823 1732 -1789 2708
rect -1565 1732 -1531 2708
rect -1307 1732 -1273 2708
rect -1049 1732 -1015 2708
rect -791 1732 -757 2708
rect -533 1732 -499 2708
rect -275 1732 -241 2708
rect -17 1732 17 2708
rect 241 1732 275 2708
rect 499 1732 533 2708
rect 757 1732 791 2708
rect 1015 1732 1049 2708
rect 1273 1732 1307 2708
rect 1531 1732 1565 2708
rect 1789 1732 1823 2708
rect 2047 1732 2081 2708
rect 2305 1732 2339 2708
rect 2563 1732 2597 2708
rect 2821 1732 2855 2708
rect 3079 1732 3113 2708
rect -3051 1648 -2883 1682
rect -2793 1648 -2625 1682
rect -2535 1648 -2367 1682
rect -2277 1648 -2109 1682
rect -2019 1648 -1851 1682
rect -1761 1648 -1593 1682
rect -1503 1648 -1335 1682
rect -1245 1648 -1077 1682
rect -987 1648 -819 1682
rect -729 1648 -561 1682
rect -471 1648 -303 1682
rect -213 1648 -45 1682
rect 45 1648 213 1682
rect 303 1648 471 1682
rect 561 1648 729 1682
rect 819 1648 987 1682
rect 1077 1648 1245 1682
rect 1335 1648 1503 1682
rect 1593 1648 1761 1682
rect 1851 1648 2019 1682
rect 2109 1648 2277 1682
rect 2367 1648 2535 1682
rect 2625 1648 2793 1682
rect 2883 1648 3051 1682
rect -3113 622 -3079 1598
rect -2855 622 -2821 1598
rect -2597 622 -2563 1598
rect -2339 622 -2305 1598
rect -2081 622 -2047 1598
rect -1823 622 -1789 1598
rect -1565 622 -1531 1598
rect -1307 622 -1273 1598
rect -1049 622 -1015 1598
rect -791 622 -757 1598
rect -533 622 -499 1598
rect -275 622 -241 1598
rect -17 622 17 1598
rect 241 622 275 1598
rect 499 622 533 1598
rect 757 622 791 1598
rect 1015 622 1049 1598
rect 1273 622 1307 1598
rect 1531 622 1565 1598
rect 1789 622 1823 1598
rect 2047 622 2081 1598
rect 2305 622 2339 1598
rect 2563 622 2597 1598
rect 2821 622 2855 1598
rect 3079 622 3113 1598
rect -3051 538 -2883 572
rect -2793 538 -2625 572
rect -2535 538 -2367 572
rect -2277 538 -2109 572
rect -2019 538 -1851 572
rect -1761 538 -1593 572
rect -1503 538 -1335 572
rect -1245 538 -1077 572
rect -987 538 -819 572
rect -729 538 -561 572
rect -471 538 -303 572
rect -213 538 -45 572
rect 45 538 213 572
rect 303 538 471 572
rect 561 538 729 572
rect 819 538 987 572
rect 1077 538 1245 572
rect 1335 538 1503 572
rect 1593 538 1761 572
rect 1851 538 2019 572
rect 2109 538 2277 572
rect 2367 538 2535 572
rect 2625 538 2793 572
rect 2883 538 3051 572
rect -3113 -488 -3079 488
rect -2855 -488 -2821 488
rect -2597 -488 -2563 488
rect -2339 -488 -2305 488
rect -2081 -488 -2047 488
rect -1823 -488 -1789 488
rect -1565 -488 -1531 488
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
rect 1531 -488 1565 488
rect 1789 -488 1823 488
rect 2047 -488 2081 488
rect 2305 -488 2339 488
rect 2563 -488 2597 488
rect 2821 -488 2855 488
rect 3079 -488 3113 488
rect -3051 -572 -2883 -538
rect -2793 -572 -2625 -538
rect -2535 -572 -2367 -538
rect -2277 -572 -2109 -538
rect -2019 -572 -1851 -538
rect -1761 -572 -1593 -538
rect -1503 -572 -1335 -538
rect -1245 -572 -1077 -538
rect -987 -572 -819 -538
rect -729 -572 -561 -538
rect -471 -572 -303 -538
rect -213 -572 -45 -538
rect 45 -572 213 -538
rect 303 -572 471 -538
rect 561 -572 729 -538
rect 819 -572 987 -538
rect 1077 -572 1245 -538
rect 1335 -572 1503 -538
rect 1593 -572 1761 -538
rect 1851 -572 2019 -538
rect 2109 -572 2277 -538
rect 2367 -572 2535 -538
rect 2625 -572 2793 -538
rect 2883 -572 3051 -538
rect -3113 -1598 -3079 -622
rect -2855 -1598 -2821 -622
rect -2597 -1598 -2563 -622
rect -2339 -1598 -2305 -622
rect -2081 -1598 -2047 -622
rect -1823 -1598 -1789 -622
rect -1565 -1598 -1531 -622
rect -1307 -1598 -1273 -622
rect -1049 -1598 -1015 -622
rect -791 -1598 -757 -622
rect -533 -1598 -499 -622
rect -275 -1598 -241 -622
rect -17 -1598 17 -622
rect 241 -1598 275 -622
rect 499 -1598 533 -622
rect 757 -1598 791 -622
rect 1015 -1598 1049 -622
rect 1273 -1598 1307 -622
rect 1531 -1598 1565 -622
rect 1789 -1598 1823 -622
rect 2047 -1598 2081 -622
rect 2305 -1598 2339 -622
rect 2563 -1598 2597 -622
rect 2821 -1598 2855 -622
rect 3079 -1598 3113 -622
rect -3051 -1682 -2883 -1648
rect -2793 -1682 -2625 -1648
rect -2535 -1682 -2367 -1648
rect -2277 -1682 -2109 -1648
rect -2019 -1682 -1851 -1648
rect -1761 -1682 -1593 -1648
rect -1503 -1682 -1335 -1648
rect -1245 -1682 -1077 -1648
rect -987 -1682 -819 -1648
rect -729 -1682 -561 -1648
rect -471 -1682 -303 -1648
rect -213 -1682 -45 -1648
rect 45 -1682 213 -1648
rect 303 -1682 471 -1648
rect 561 -1682 729 -1648
rect 819 -1682 987 -1648
rect 1077 -1682 1245 -1648
rect 1335 -1682 1503 -1648
rect 1593 -1682 1761 -1648
rect 1851 -1682 2019 -1648
rect 2109 -1682 2277 -1648
rect 2367 -1682 2535 -1648
rect 2625 -1682 2793 -1648
rect 2883 -1682 3051 -1648
rect -3113 -2708 -3079 -1732
rect -2855 -2708 -2821 -1732
rect -2597 -2708 -2563 -1732
rect -2339 -2708 -2305 -1732
rect -2081 -2708 -2047 -1732
rect -1823 -2708 -1789 -1732
rect -1565 -2708 -1531 -1732
rect -1307 -2708 -1273 -1732
rect -1049 -2708 -1015 -1732
rect -791 -2708 -757 -1732
rect -533 -2708 -499 -1732
rect -275 -2708 -241 -1732
rect -17 -2708 17 -1732
rect 241 -2708 275 -1732
rect 499 -2708 533 -1732
rect 757 -2708 791 -1732
rect 1015 -2708 1049 -1732
rect 1273 -2708 1307 -1732
rect 1531 -2708 1565 -1732
rect 1789 -2708 1823 -1732
rect 2047 -2708 2081 -1732
rect 2305 -2708 2339 -1732
rect 2563 -2708 2597 -1732
rect 2821 -2708 2855 -1732
rect 3079 -2708 3113 -1732
rect -3051 -2792 -2883 -2758
rect -2793 -2792 -2625 -2758
rect -2535 -2792 -2367 -2758
rect -2277 -2792 -2109 -2758
rect -2019 -2792 -1851 -2758
rect -1761 -2792 -1593 -2758
rect -1503 -2792 -1335 -2758
rect -1245 -2792 -1077 -2758
rect -987 -2792 -819 -2758
rect -729 -2792 -561 -2758
rect -471 -2792 -303 -2758
rect -213 -2792 -45 -2758
rect 45 -2792 213 -2758
rect 303 -2792 471 -2758
rect 561 -2792 729 -2758
rect 819 -2792 987 -2758
rect 1077 -2792 1245 -2758
rect 1335 -2792 1503 -2758
rect 1593 -2792 1761 -2758
rect 1851 -2792 2019 -2758
rect 2109 -2792 2277 -2758
rect 2367 -2792 2535 -2758
rect 2625 -2792 2793 -2758
rect 2883 -2792 3051 -2758
<< metal1 >>
rect -3063 2792 -2871 2798
rect -3063 2758 -3051 2792
rect -2883 2758 -2871 2792
rect -3063 2752 -2871 2758
rect -2805 2792 -2613 2798
rect -2805 2758 -2793 2792
rect -2625 2758 -2613 2792
rect -2805 2752 -2613 2758
rect -2547 2792 -2355 2798
rect -2547 2758 -2535 2792
rect -2367 2758 -2355 2792
rect -2547 2752 -2355 2758
rect -2289 2792 -2097 2798
rect -2289 2758 -2277 2792
rect -2109 2758 -2097 2792
rect -2289 2752 -2097 2758
rect -2031 2792 -1839 2798
rect -2031 2758 -2019 2792
rect -1851 2758 -1839 2792
rect -2031 2752 -1839 2758
rect -1773 2792 -1581 2798
rect -1773 2758 -1761 2792
rect -1593 2758 -1581 2792
rect -1773 2752 -1581 2758
rect -1515 2792 -1323 2798
rect -1515 2758 -1503 2792
rect -1335 2758 -1323 2792
rect -1515 2752 -1323 2758
rect -1257 2792 -1065 2798
rect -1257 2758 -1245 2792
rect -1077 2758 -1065 2792
rect -1257 2752 -1065 2758
rect -999 2792 -807 2798
rect -999 2758 -987 2792
rect -819 2758 -807 2792
rect -999 2752 -807 2758
rect -741 2792 -549 2798
rect -741 2758 -729 2792
rect -561 2758 -549 2792
rect -741 2752 -549 2758
rect -483 2792 -291 2798
rect -483 2758 -471 2792
rect -303 2758 -291 2792
rect -483 2752 -291 2758
rect -225 2792 -33 2798
rect -225 2758 -213 2792
rect -45 2758 -33 2792
rect -225 2752 -33 2758
rect 33 2792 225 2798
rect 33 2758 45 2792
rect 213 2758 225 2792
rect 33 2752 225 2758
rect 291 2792 483 2798
rect 291 2758 303 2792
rect 471 2758 483 2792
rect 291 2752 483 2758
rect 549 2792 741 2798
rect 549 2758 561 2792
rect 729 2758 741 2792
rect 549 2752 741 2758
rect 807 2792 999 2798
rect 807 2758 819 2792
rect 987 2758 999 2792
rect 807 2752 999 2758
rect 1065 2792 1257 2798
rect 1065 2758 1077 2792
rect 1245 2758 1257 2792
rect 1065 2752 1257 2758
rect 1323 2792 1515 2798
rect 1323 2758 1335 2792
rect 1503 2758 1515 2792
rect 1323 2752 1515 2758
rect 1581 2792 1773 2798
rect 1581 2758 1593 2792
rect 1761 2758 1773 2792
rect 1581 2752 1773 2758
rect 1839 2792 2031 2798
rect 1839 2758 1851 2792
rect 2019 2758 2031 2792
rect 1839 2752 2031 2758
rect 2097 2792 2289 2798
rect 2097 2758 2109 2792
rect 2277 2758 2289 2792
rect 2097 2752 2289 2758
rect 2355 2792 2547 2798
rect 2355 2758 2367 2792
rect 2535 2758 2547 2792
rect 2355 2752 2547 2758
rect 2613 2792 2805 2798
rect 2613 2758 2625 2792
rect 2793 2758 2805 2792
rect 2613 2752 2805 2758
rect 2871 2792 3063 2798
rect 2871 2758 2883 2792
rect 3051 2758 3063 2792
rect 2871 2752 3063 2758
rect -3119 2708 -3073 2720
rect -3119 1732 -3113 2708
rect -3079 1732 -3073 2708
rect -3119 1720 -3073 1732
rect -2861 2708 -2815 2720
rect -2861 1732 -2855 2708
rect -2821 1732 -2815 2708
rect -2861 1720 -2815 1732
rect -2603 2708 -2557 2720
rect -2603 1732 -2597 2708
rect -2563 1732 -2557 2708
rect -2603 1720 -2557 1732
rect -2345 2708 -2299 2720
rect -2345 1732 -2339 2708
rect -2305 1732 -2299 2708
rect -2345 1720 -2299 1732
rect -2087 2708 -2041 2720
rect -2087 1732 -2081 2708
rect -2047 1732 -2041 2708
rect -2087 1720 -2041 1732
rect -1829 2708 -1783 2720
rect -1829 1732 -1823 2708
rect -1789 1732 -1783 2708
rect -1829 1720 -1783 1732
rect -1571 2708 -1525 2720
rect -1571 1732 -1565 2708
rect -1531 1732 -1525 2708
rect -1571 1720 -1525 1732
rect -1313 2708 -1267 2720
rect -1313 1732 -1307 2708
rect -1273 1732 -1267 2708
rect -1313 1720 -1267 1732
rect -1055 2708 -1009 2720
rect -1055 1732 -1049 2708
rect -1015 1732 -1009 2708
rect -1055 1720 -1009 1732
rect -797 2708 -751 2720
rect -797 1732 -791 2708
rect -757 1732 -751 2708
rect -797 1720 -751 1732
rect -539 2708 -493 2720
rect -539 1732 -533 2708
rect -499 1732 -493 2708
rect -539 1720 -493 1732
rect -281 2708 -235 2720
rect -281 1732 -275 2708
rect -241 1732 -235 2708
rect -281 1720 -235 1732
rect -23 2708 23 2720
rect -23 1732 -17 2708
rect 17 1732 23 2708
rect -23 1720 23 1732
rect 235 2708 281 2720
rect 235 1732 241 2708
rect 275 1732 281 2708
rect 235 1720 281 1732
rect 493 2708 539 2720
rect 493 1732 499 2708
rect 533 1732 539 2708
rect 493 1720 539 1732
rect 751 2708 797 2720
rect 751 1732 757 2708
rect 791 1732 797 2708
rect 751 1720 797 1732
rect 1009 2708 1055 2720
rect 1009 1732 1015 2708
rect 1049 1732 1055 2708
rect 1009 1720 1055 1732
rect 1267 2708 1313 2720
rect 1267 1732 1273 2708
rect 1307 1732 1313 2708
rect 1267 1720 1313 1732
rect 1525 2708 1571 2720
rect 1525 1732 1531 2708
rect 1565 1732 1571 2708
rect 1525 1720 1571 1732
rect 1783 2708 1829 2720
rect 1783 1732 1789 2708
rect 1823 1732 1829 2708
rect 1783 1720 1829 1732
rect 2041 2708 2087 2720
rect 2041 1732 2047 2708
rect 2081 1732 2087 2708
rect 2041 1720 2087 1732
rect 2299 2708 2345 2720
rect 2299 1732 2305 2708
rect 2339 1732 2345 2708
rect 2299 1720 2345 1732
rect 2557 2708 2603 2720
rect 2557 1732 2563 2708
rect 2597 1732 2603 2708
rect 2557 1720 2603 1732
rect 2815 2708 2861 2720
rect 2815 1732 2821 2708
rect 2855 1732 2861 2708
rect 2815 1720 2861 1732
rect 3073 2708 3119 2720
rect 3073 1732 3079 2708
rect 3113 1732 3119 2708
rect 3073 1720 3119 1732
rect -3063 1682 -2871 1688
rect -3063 1648 -3051 1682
rect -2883 1648 -2871 1682
rect -3063 1642 -2871 1648
rect -2805 1682 -2613 1688
rect -2805 1648 -2793 1682
rect -2625 1648 -2613 1682
rect -2805 1642 -2613 1648
rect -2547 1682 -2355 1688
rect -2547 1648 -2535 1682
rect -2367 1648 -2355 1682
rect -2547 1642 -2355 1648
rect -2289 1682 -2097 1688
rect -2289 1648 -2277 1682
rect -2109 1648 -2097 1682
rect -2289 1642 -2097 1648
rect -2031 1682 -1839 1688
rect -2031 1648 -2019 1682
rect -1851 1648 -1839 1682
rect -2031 1642 -1839 1648
rect -1773 1682 -1581 1688
rect -1773 1648 -1761 1682
rect -1593 1648 -1581 1682
rect -1773 1642 -1581 1648
rect -1515 1682 -1323 1688
rect -1515 1648 -1503 1682
rect -1335 1648 -1323 1682
rect -1515 1642 -1323 1648
rect -1257 1682 -1065 1688
rect -1257 1648 -1245 1682
rect -1077 1648 -1065 1682
rect -1257 1642 -1065 1648
rect -999 1682 -807 1688
rect -999 1648 -987 1682
rect -819 1648 -807 1682
rect -999 1642 -807 1648
rect -741 1682 -549 1688
rect -741 1648 -729 1682
rect -561 1648 -549 1682
rect -741 1642 -549 1648
rect -483 1682 -291 1688
rect -483 1648 -471 1682
rect -303 1648 -291 1682
rect -483 1642 -291 1648
rect -225 1682 -33 1688
rect -225 1648 -213 1682
rect -45 1648 -33 1682
rect -225 1642 -33 1648
rect 33 1682 225 1688
rect 33 1648 45 1682
rect 213 1648 225 1682
rect 33 1642 225 1648
rect 291 1682 483 1688
rect 291 1648 303 1682
rect 471 1648 483 1682
rect 291 1642 483 1648
rect 549 1682 741 1688
rect 549 1648 561 1682
rect 729 1648 741 1682
rect 549 1642 741 1648
rect 807 1682 999 1688
rect 807 1648 819 1682
rect 987 1648 999 1682
rect 807 1642 999 1648
rect 1065 1682 1257 1688
rect 1065 1648 1077 1682
rect 1245 1648 1257 1682
rect 1065 1642 1257 1648
rect 1323 1682 1515 1688
rect 1323 1648 1335 1682
rect 1503 1648 1515 1682
rect 1323 1642 1515 1648
rect 1581 1682 1773 1688
rect 1581 1648 1593 1682
rect 1761 1648 1773 1682
rect 1581 1642 1773 1648
rect 1839 1682 2031 1688
rect 1839 1648 1851 1682
rect 2019 1648 2031 1682
rect 1839 1642 2031 1648
rect 2097 1682 2289 1688
rect 2097 1648 2109 1682
rect 2277 1648 2289 1682
rect 2097 1642 2289 1648
rect 2355 1682 2547 1688
rect 2355 1648 2367 1682
rect 2535 1648 2547 1682
rect 2355 1642 2547 1648
rect 2613 1682 2805 1688
rect 2613 1648 2625 1682
rect 2793 1648 2805 1682
rect 2613 1642 2805 1648
rect 2871 1682 3063 1688
rect 2871 1648 2883 1682
rect 3051 1648 3063 1682
rect 2871 1642 3063 1648
rect -3119 1598 -3073 1610
rect -3119 622 -3113 1598
rect -3079 622 -3073 1598
rect -3119 610 -3073 622
rect -2861 1598 -2815 1610
rect -2861 622 -2855 1598
rect -2821 622 -2815 1598
rect -2861 610 -2815 622
rect -2603 1598 -2557 1610
rect -2603 622 -2597 1598
rect -2563 622 -2557 1598
rect -2603 610 -2557 622
rect -2345 1598 -2299 1610
rect -2345 622 -2339 1598
rect -2305 622 -2299 1598
rect -2345 610 -2299 622
rect -2087 1598 -2041 1610
rect -2087 622 -2081 1598
rect -2047 622 -2041 1598
rect -2087 610 -2041 622
rect -1829 1598 -1783 1610
rect -1829 622 -1823 1598
rect -1789 622 -1783 1598
rect -1829 610 -1783 622
rect -1571 1598 -1525 1610
rect -1571 622 -1565 1598
rect -1531 622 -1525 1598
rect -1571 610 -1525 622
rect -1313 1598 -1267 1610
rect -1313 622 -1307 1598
rect -1273 622 -1267 1598
rect -1313 610 -1267 622
rect -1055 1598 -1009 1610
rect -1055 622 -1049 1598
rect -1015 622 -1009 1598
rect -1055 610 -1009 622
rect -797 1598 -751 1610
rect -797 622 -791 1598
rect -757 622 -751 1598
rect -797 610 -751 622
rect -539 1598 -493 1610
rect -539 622 -533 1598
rect -499 622 -493 1598
rect -539 610 -493 622
rect -281 1598 -235 1610
rect -281 622 -275 1598
rect -241 622 -235 1598
rect -281 610 -235 622
rect -23 1598 23 1610
rect -23 622 -17 1598
rect 17 622 23 1598
rect -23 610 23 622
rect 235 1598 281 1610
rect 235 622 241 1598
rect 275 622 281 1598
rect 235 610 281 622
rect 493 1598 539 1610
rect 493 622 499 1598
rect 533 622 539 1598
rect 493 610 539 622
rect 751 1598 797 1610
rect 751 622 757 1598
rect 791 622 797 1598
rect 751 610 797 622
rect 1009 1598 1055 1610
rect 1009 622 1015 1598
rect 1049 622 1055 1598
rect 1009 610 1055 622
rect 1267 1598 1313 1610
rect 1267 622 1273 1598
rect 1307 622 1313 1598
rect 1267 610 1313 622
rect 1525 1598 1571 1610
rect 1525 622 1531 1598
rect 1565 622 1571 1598
rect 1525 610 1571 622
rect 1783 1598 1829 1610
rect 1783 622 1789 1598
rect 1823 622 1829 1598
rect 1783 610 1829 622
rect 2041 1598 2087 1610
rect 2041 622 2047 1598
rect 2081 622 2087 1598
rect 2041 610 2087 622
rect 2299 1598 2345 1610
rect 2299 622 2305 1598
rect 2339 622 2345 1598
rect 2299 610 2345 622
rect 2557 1598 2603 1610
rect 2557 622 2563 1598
rect 2597 622 2603 1598
rect 2557 610 2603 622
rect 2815 1598 2861 1610
rect 2815 622 2821 1598
rect 2855 622 2861 1598
rect 2815 610 2861 622
rect 3073 1598 3119 1610
rect 3073 622 3079 1598
rect 3113 622 3119 1598
rect 3073 610 3119 622
rect -3063 572 -2871 578
rect -3063 538 -3051 572
rect -2883 538 -2871 572
rect -3063 532 -2871 538
rect -2805 572 -2613 578
rect -2805 538 -2793 572
rect -2625 538 -2613 572
rect -2805 532 -2613 538
rect -2547 572 -2355 578
rect -2547 538 -2535 572
rect -2367 538 -2355 572
rect -2547 532 -2355 538
rect -2289 572 -2097 578
rect -2289 538 -2277 572
rect -2109 538 -2097 572
rect -2289 532 -2097 538
rect -2031 572 -1839 578
rect -2031 538 -2019 572
rect -1851 538 -1839 572
rect -2031 532 -1839 538
rect -1773 572 -1581 578
rect -1773 538 -1761 572
rect -1593 538 -1581 572
rect -1773 532 -1581 538
rect -1515 572 -1323 578
rect -1515 538 -1503 572
rect -1335 538 -1323 572
rect -1515 532 -1323 538
rect -1257 572 -1065 578
rect -1257 538 -1245 572
rect -1077 538 -1065 572
rect -1257 532 -1065 538
rect -999 572 -807 578
rect -999 538 -987 572
rect -819 538 -807 572
rect -999 532 -807 538
rect -741 572 -549 578
rect -741 538 -729 572
rect -561 538 -549 572
rect -741 532 -549 538
rect -483 572 -291 578
rect -483 538 -471 572
rect -303 538 -291 572
rect -483 532 -291 538
rect -225 572 -33 578
rect -225 538 -213 572
rect -45 538 -33 572
rect -225 532 -33 538
rect 33 572 225 578
rect 33 538 45 572
rect 213 538 225 572
rect 33 532 225 538
rect 291 572 483 578
rect 291 538 303 572
rect 471 538 483 572
rect 291 532 483 538
rect 549 572 741 578
rect 549 538 561 572
rect 729 538 741 572
rect 549 532 741 538
rect 807 572 999 578
rect 807 538 819 572
rect 987 538 999 572
rect 807 532 999 538
rect 1065 572 1257 578
rect 1065 538 1077 572
rect 1245 538 1257 572
rect 1065 532 1257 538
rect 1323 572 1515 578
rect 1323 538 1335 572
rect 1503 538 1515 572
rect 1323 532 1515 538
rect 1581 572 1773 578
rect 1581 538 1593 572
rect 1761 538 1773 572
rect 1581 532 1773 538
rect 1839 572 2031 578
rect 1839 538 1851 572
rect 2019 538 2031 572
rect 1839 532 2031 538
rect 2097 572 2289 578
rect 2097 538 2109 572
rect 2277 538 2289 572
rect 2097 532 2289 538
rect 2355 572 2547 578
rect 2355 538 2367 572
rect 2535 538 2547 572
rect 2355 532 2547 538
rect 2613 572 2805 578
rect 2613 538 2625 572
rect 2793 538 2805 572
rect 2613 532 2805 538
rect 2871 572 3063 578
rect 2871 538 2883 572
rect 3051 538 3063 572
rect 2871 532 3063 538
rect -3119 488 -3073 500
rect -3119 -488 -3113 488
rect -3079 -488 -3073 488
rect -3119 -500 -3073 -488
rect -2861 488 -2815 500
rect -2861 -488 -2855 488
rect -2821 -488 -2815 488
rect -2861 -500 -2815 -488
rect -2603 488 -2557 500
rect -2603 -488 -2597 488
rect -2563 -488 -2557 488
rect -2603 -500 -2557 -488
rect -2345 488 -2299 500
rect -2345 -488 -2339 488
rect -2305 -488 -2299 488
rect -2345 -500 -2299 -488
rect -2087 488 -2041 500
rect -2087 -488 -2081 488
rect -2047 -488 -2041 488
rect -2087 -500 -2041 -488
rect -1829 488 -1783 500
rect -1829 -488 -1823 488
rect -1789 -488 -1783 488
rect -1829 -500 -1783 -488
rect -1571 488 -1525 500
rect -1571 -488 -1565 488
rect -1531 -488 -1525 488
rect -1571 -500 -1525 -488
rect -1313 488 -1267 500
rect -1313 -488 -1307 488
rect -1273 -488 -1267 488
rect -1313 -500 -1267 -488
rect -1055 488 -1009 500
rect -1055 -488 -1049 488
rect -1015 -488 -1009 488
rect -1055 -500 -1009 -488
rect -797 488 -751 500
rect -797 -488 -791 488
rect -757 -488 -751 488
rect -797 -500 -751 -488
rect -539 488 -493 500
rect -539 -488 -533 488
rect -499 -488 -493 488
rect -539 -500 -493 -488
rect -281 488 -235 500
rect -281 -488 -275 488
rect -241 -488 -235 488
rect -281 -500 -235 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 235 488 281 500
rect 235 -488 241 488
rect 275 -488 281 488
rect 235 -500 281 -488
rect 493 488 539 500
rect 493 -488 499 488
rect 533 -488 539 488
rect 493 -500 539 -488
rect 751 488 797 500
rect 751 -488 757 488
rect 791 -488 797 488
rect 751 -500 797 -488
rect 1009 488 1055 500
rect 1009 -488 1015 488
rect 1049 -488 1055 488
rect 1009 -500 1055 -488
rect 1267 488 1313 500
rect 1267 -488 1273 488
rect 1307 -488 1313 488
rect 1267 -500 1313 -488
rect 1525 488 1571 500
rect 1525 -488 1531 488
rect 1565 -488 1571 488
rect 1525 -500 1571 -488
rect 1783 488 1829 500
rect 1783 -488 1789 488
rect 1823 -488 1829 488
rect 1783 -500 1829 -488
rect 2041 488 2087 500
rect 2041 -488 2047 488
rect 2081 -488 2087 488
rect 2041 -500 2087 -488
rect 2299 488 2345 500
rect 2299 -488 2305 488
rect 2339 -488 2345 488
rect 2299 -500 2345 -488
rect 2557 488 2603 500
rect 2557 -488 2563 488
rect 2597 -488 2603 488
rect 2557 -500 2603 -488
rect 2815 488 2861 500
rect 2815 -488 2821 488
rect 2855 -488 2861 488
rect 2815 -500 2861 -488
rect 3073 488 3119 500
rect 3073 -488 3079 488
rect 3113 -488 3119 488
rect 3073 -500 3119 -488
rect -3063 -538 -2871 -532
rect -3063 -572 -3051 -538
rect -2883 -572 -2871 -538
rect -3063 -578 -2871 -572
rect -2805 -538 -2613 -532
rect -2805 -572 -2793 -538
rect -2625 -572 -2613 -538
rect -2805 -578 -2613 -572
rect -2547 -538 -2355 -532
rect -2547 -572 -2535 -538
rect -2367 -572 -2355 -538
rect -2547 -578 -2355 -572
rect -2289 -538 -2097 -532
rect -2289 -572 -2277 -538
rect -2109 -572 -2097 -538
rect -2289 -578 -2097 -572
rect -2031 -538 -1839 -532
rect -2031 -572 -2019 -538
rect -1851 -572 -1839 -538
rect -2031 -578 -1839 -572
rect -1773 -538 -1581 -532
rect -1773 -572 -1761 -538
rect -1593 -572 -1581 -538
rect -1773 -578 -1581 -572
rect -1515 -538 -1323 -532
rect -1515 -572 -1503 -538
rect -1335 -572 -1323 -538
rect -1515 -578 -1323 -572
rect -1257 -538 -1065 -532
rect -1257 -572 -1245 -538
rect -1077 -572 -1065 -538
rect -1257 -578 -1065 -572
rect -999 -538 -807 -532
rect -999 -572 -987 -538
rect -819 -572 -807 -538
rect -999 -578 -807 -572
rect -741 -538 -549 -532
rect -741 -572 -729 -538
rect -561 -572 -549 -538
rect -741 -578 -549 -572
rect -483 -538 -291 -532
rect -483 -572 -471 -538
rect -303 -572 -291 -538
rect -483 -578 -291 -572
rect -225 -538 -33 -532
rect -225 -572 -213 -538
rect -45 -572 -33 -538
rect -225 -578 -33 -572
rect 33 -538 225 -532
rect 33 -572 45 -538
rect 213 -572 225 -538
rect 33 -578 225 -572
rect 291 -538 483 -532
rect 291 -572 303 -538
rect 471 -572 483 -538
rect 291 -578 483 -572
rect 549 -538 741 -532
rect 549 -572 561 -538
rect 729 -572 741 -538
rect 549 -578 741 -572
rect 807 -538 999 -532
rect 807 -572 819 -538
rect 987 -572 999 -538
rect 807 -578 999 -572
rect 1065 -538 1257 -532
rect 1065 -572 1077 -538
rect 1245 -572 1257 -538
rect 1065 -578 1257 -572
rect 1323 -538 1515 -532
rect 1323 -572 1335 -538
rect 1503 -572 1515 -538
rect 1323 -578 1515 -572
rect 1581 -538 1773 -532
rect 1581 -572 1593 -538
rect 1761 -572 1773 -538
rect 1581 -578 1773 -572
rect 1839 -538 2031 -532
rect 1839 -572 1851 -538
rect 2019 -572 2031 -538
rect 1839 -578 2031 -572
rect 2097 -538 2289 -532
rect 2097 -572 2109 -538
rect 2277 -572 2289 -538
rect 2097 -578 2289 -572
rect 2355 -538 2547 -532
rect 2355 -572 2367 -538
rect 2535 -572 2547 -538
rect 2355 -578 2547 -572
rect 2613 -538 2805 -532
rect 2613 -572 2625 -538
rect 2793 -572 2805 -538
rect 2613 -578 2805 -572
rect 2871 -538 3063 -532
rect 2871 -572 2883 -538
rect 3051 -572 3063 -538
rect 2871 -578 3063 -572
rect -3119 -622 -3073 -610
rect -3119 -1598 -3113 -622
rect -3079 -1598 -3073 -622
rect -3119 -1610 -3073 -1598
rect -2861 -622 -2815 -610
rect -2861 -1598 -2855 -622
rect -2821 -1598 -2815 -622
rect -2861 -1610 -2815 -1598
rect -2603 -622 -2557 -610
rect -2603 -1598 -2597 -622
rect -2563 -1598 -2557 -622
rect -2603 -1610 -2557 -1598
rect -2345 -622 -2299 -610
rect -2345 -1598 -2339 -622
rect -2305 -1598 -2299 -622
rect -2345 -1610 -2299 -1598
rect -2087 -622 -2041 -610
rect -2087 -1598 -2081 -622
rect -2047 -1598 -2041 -622
rect -2087 -1610 -2041 -1598
rect -1829 -622 -1783 -610
rect -1829 -1598 -1823 -622
rect -1789 -1598 -1783 -622
rect -1829 -1610 -1783 -1598
rect -1571 -622 -1525 -610
rect -1571 -1598 -1565 -622
rect -1531 -1598 -1525 -622
rect -1571 -1610 -1525 -1598
rect -1313 -622 -1267 -610
rect -1313 -1598 -1307 -622
rect -1273 -1598 -1267 -622
rect -1313 -1610 -1267 -1598
rect -1055 -622 -1009 -610
rect -1055 -1598 -1049 -622
rect -1015 -1598 -1009 -622
rect -1055 -1610 -1009 -1598
rect -797 -622 -751 -610
rect -797 -1598 -791 -622
rect -757 -1598 -751 -622
rect -797 -1610 -751 -1598
rect -539 -622 -493 -610
rect -539 -1598 -533 -622
rect -499 -1598 -493 -622
rect -539 -1610 -493 -1598
rect -281 -622 -235 -610
rect -281 -1598 -275 -622
rect -241 -1598 -235 -622
rect -281 -1610 -235 -1598
rect -23 -622 23 -610
rect -23 -1598 -17 -622
rect 17 -1598 23 -622
rect -23 -1610 23 -1598
rect 235 -622 281 -610
rect 235 -1598 241 -622
rect 275 -1598 281 -622
rect 235 -1610 281 -1598
rect 493 -622 539 -610
rect 493 -1598 499 -622
rect 533 -1598 539 -622
rect 493 -1610 539 -1598
rect 751 -622 797 -610
rect 751 -1598 757 -622
rect 791 -1598 797 -622
rect 751 -1610 797 -1598
rect 1009 -622 1055 -610
rect 1009 -1598 1015 -622
rect 1049 -1598 1055 -622
rect 1009 -1610 1055 -1598
rect 1267 -622 1313 -610
rect 1267 -1598 1273 -622
rect 1307 -1598 1313 -622
rect 1267 -1610 1313 -1598
rect 1525 -622 1571 -610
rect 1525 -1598 1531 -622
rect 1565 -1598 1571 -622
rect 1525 -1610 1571 -1598
rect 1783 -622 1829 -610
rect 1783 -1598 1789 -622
rect 1823 -1598 1829 -622
rect 1783 -1610 1829 -1598
rect 2041 -622 2087 -610
rect 2041 -1598 2047 -622
rect 2081 -1598 2087 -622
rect 2041 -1610 2087 -1598
rect 2299 -622 2345 -610
rect 2299 -1598 2305 -622
rect 2339 -1598 2345 -622
rect 2299 -1610 2345 -1598
rect 2557 -622 2603 -610
rect 2557 -1598 2563 -622
rect 2597 -1598 2603 -622
rect 2557 -1610 2603 -1598
rect 2815 -622 2861 -610
rect 2815 -1598 2821 -622
rect 2855 -1598 2861 -622
rect 2815 -1610 2861 -1598
rect 3073 -622 3119 -610
rect 3073 -1598 3079 -622
rect 3113 -1598 3119 -622
rect 3073 -1610 3119 -1598
rect -3063 -1648 -2871 -1642
rect -3063 -1682 -3051 -1648
rect -2883 -1682 -2871 -1648
rect -3063 -1688 -2871 -1682
rect -2805 -1648 -2613 -1642
rect -2805 -1682 -2793 -1648
rect -2625 -1682 -2613 -1648
rect -2805 -1688 -2613 -1682
rect -2547 -1648 -2355 -1642
rect -2547 -1682 -2535 -1648
rect -2367 -1682 -2355 -1648
rect -2547 -1688 -2355 -1682
rect -2289 -1648 -2097 -1642
rect -2289 -1682 -2277 -1648
rect -2109 -1682 -2097 -1648
rect -2289 -1688 -2097 -1682
rect -2031 -1648 -1839 -1642
rect -2031 -1682 -2019 -1648
rect -1851 -1682 -1839 -1648
rect -2031 -1688 -1839 -1682
rect -1773 -1648 -1581 -1642
rect -1773 -1682 -1761 -1648
rect -1593 -1682 -1581 -1648
rect -1773 -1688 -1581 -1682
rect -1515 -1648 -1323 -1642
rect -1515 -1682 -1503 -1648
rect -1335 -1682 -1323 -1648
rect -1515 -1688 -1323 -1682
rect -1257 -1648 -1065 -1642
rect -1257 -1682 -1245 -1648
rect -1077 -1682 -1065 -1648
rect -1257 -1688 -1065 -1682
rect -999 -1648 -807 -1642
rect -999 -1682 -987 -1648
rect -819 -1682 -807 -1648
rect -999 -1688 -807 -1682
rect -741 -1648 -549 -1642
rect -741 -1682 -729 -1648
rect -561 -1682 -549 -1648
rect -741 -1688 -549 -1682
rect -483 -1648 -291 -1642
rect -483 -1682 -471 -1648
rect -303 -1682 -291 -1648
rect -483 -1688 -291 -1682
rect -225 -1648 -33 -1642
rect -225 -1682 -213 -1648
rect -45 -1682 -33 -1648
rect -225 -1688 -33 -1682
rect 33 -1648 225 -1642
rect 33 -1682 45 -1648
rect 213 -1682 225 -1648
rect 33 -1688 225 -1682
rect 291 -1648 483 -1642
rect 291 -1682 303 -1648
rect 471 -1682 483 -1648
rect 291 -1688 483 -1682
rect 549 -1648 741 -1642
rect 549 -1682 561 -1648
rect 729 -1682 741 -1648
rect 549 -1688 741 -1682
rect 807 -1648 999 -1642
rect 807 -1682 819 -1648
rect 987 -1682 999 -1648
rect 807 -1688 999 -1682
rect 1065 -1648 1257 -1642
rect 1065 -1682 1077 -1648
rect 1245 -1682 1257 -1648
rect 1065 -1688 1257 -1682
rect 1323 -1648 1515 -1642
rect 1323 -1682 1335 -1648
rect 1503 -1682 1515 -1648
rect 1323 -1688 1515 -1682
rect 1581 -1648 1773 -1642
rect 1581 -1682 1593 -1648
rect 1761 -1682 1773 -1648
rect 1581 -1688 1773 -1682
rect 1839 -1648 2031 -1642
rect 1839 -1682 1851 -1648
rect 2019 -1682 2031 -1648
rect 1839 -1688 2031 -1682
rect 2097 -1648 2289 -1642
rect 2097 -1682 2109 -1648
rect 2277 -1682 2289 -1648
rect 2097 -1688 2289 -1682
rect 2355 -1648 2547 -1642
rect 2355 -1682 2367 -1648
rect 2535 -1682 2547 -1648
rect 2355 -1688 2547 -1682
rect 2613 -1648 2805 -1642
rect 2613 -1682 2625 -1648
rect 2793 -1682 2805 -1648
rect 2613 -1688 2805 -1682
rect 2871 -1648 3063 -1642
rect 2871 -1682 2883 -1648
rect 3051 -1682 3063 -1648
rect 2871 -1688 3063 -1682
rect -3119 -1732 -3073 -1720
rect -3119 -2708 -3113 -1732
rect -3079 -2708 -3073 -1732
rect -3119 -2720 -3073 -2708
rect -2861 -1732 -2815 -1720
rect -2861 -2708 -2855 -1732
rect -2821 -2708 -2815 -1732
rect -2861 -2720 -2815 -2708
rect -2603 -1732 -2557 -1720
rect -2603 -2708 -2597 -1732
rect -2563 -2708 -2557 -1732
rect -2603 -2720 -2557 -2708
rect -2345 -1732 -2299 -1720
rect -2345 -2708 -2339 -1732
rect -2305 -2708 -2299 -1732
rect -2345 -2720 -2299 -2708
rect -2087 -1732 -2041 -1720
rect -2087 -2708 -2081 -1732
rect -2047 -2708 -2041 -1732
rect -2087 -2720 -2041 -2708
rect -1829 -1732 -1783 -1720
rect -1829 -2708 -1823 -1732
rect -1789 -2708 -1783 -1732
rect -1829 -2720 -1783 -2708
rect -1571 -1732 -1525 -1720
rect -1571 -2708 -1565 -1732
rect -1531 -2708 -1525 -1732
rect -1571 -2720 -1525 -2708
rect -1313 -1732 -1267 -1720
rect -1313 -2708 -1307 -1732
rect -1273 -2708 -1267 -1732
rect -1313 -2720 -1267 -2708
rect -1055 -1732 -1009 -1720
rect -1055 -2708 -1049 -1732
rect -1015 -2708 -1009 -1732
rect -1055 -2720 -1009 -2708
rect -797 -1732 -751 -1720
rect -797 -2708 -791 -1732
rect -757 -2708 -751 -1732
rect -797 -2720 -751 -2708
rect -539 -1732 -493 -1720
rect -539 -2708 -533 -1732
rect -499 -2708 -493 -1732
rect -539 -2720 -493 -2708
rect -281 -1732 -235 -1720
rect -281 -2708 -275 -1732
rect -241 -2708 -235 -1732
rect -281 -2720 -235 -2708
rect -23 -1732 23 -1720
rect -23 -2708 -17 -1732
rect 17 -2708 23 -1732
rect -23 -2720 23 -2708
rect 235 -1732 281 -1720
rect 235 -2708 241 -1732
rect 275 -2708 281 -1732
rect 235 -2720 281 -2708
rect 493 -1732 539 -1720
rect 493 -2708 499 -1732
rect 533 -2708 539 -1732
rect 493 -2720 539 -2708
rect 751 -1732 797 -1720
rect 751 -2708 757 -1732
rect 791 -2708 797 -1732
rect 751 -2720 797 -2708
rect 1009 -1732 1055 -1720
rect 1009 -2708 1015 -1732
rect 1049 -2708 1055 -1732
rect 1009 -2720 1055 -2708
rect 1267 -1732 1313 -1720
rect 1267 -2708 1273 -1732
rect 1307 -2708 1313 -1732
rect 1267 -2720 1313 -2708
rect 1525 -1732 1571 -1720
rect 1525 -2708 1531 -1732
rect 1565 -2708 1571 -1732
rect 1525 -2720 1571 -2708
rect 1783 -1732 1829 -1720
rect 1783 -2708 1789 -1732
rect 1823 -2708 1829 -1732
rect 1783 -2720 1829 -2708
rect 2041 -1732 2087 -1720
rect 2041 -2708 2047 -1732
rect 2081 -2708 2087 -1732
rect 2041 -2720 2087 -2708
rect 2299 -1732 2345 -1720
rect 2299 -2708 2305 -1732
rect 2339 -2708 2345 -1732
rect 2299 -2720 2345 -2708
rect 2557 -1732 2603 -1720
rect 2557 -2708 2563 -1732
rect 2597 -2708 2603 -1732
rect 2557 -2720 2603 -2708
rect 2815 -1732 2861 -1720
rect 2815 -2708 2821 -1732
rect 2855 -2708 2861 -1732
rect 2815 -2720 2861 -2708
rect 3073 -1732 3119 -1720
rect 3073 -2708 3079 -1732
rect 3113 -2708 3119 -1732
rect 3073 -2720 3119 -2708
rect -3063 -2758 -2871 -2752
rect -3063 -2792 -3051 -2758
rect -2883 -2792 -2871 -2758
rect -3063 -2798 -2871 -2792
rect -2805 -2758 -2613 -2752
rect -2805 -2792 -2793 -2758
rect -2625 -2792 -2613 -2758
rect -2805 -2798 -2613 -2792
rect -2547 -2758 -2355 -2752
rect -2547 -2792 -2535 -2758
rect -2367 -2792 -2355 -2758
rect -2547 -2798 -2355 -2792
rect -2289 -2758 -2097 -2752
rect -2289 -2792 -2277 -2758
rect -2109 -2792 -2097 -2758
rect -2289 -2798 -2097 -2792
rect -2031 -2758 -1839 -2752
rect -2031 -2792 -2019 -2758
rect -1851 -2792 -1839 -2758
rect -2031 -2798 -1839 -2792
rect -1773 -2758 -1581 -2752
rect -1773 -2792 -1761 -2758
rect -1593 -2792 -1581 -2758
rect -1773 -2798 -1581 -2792
rect -1515 -2758 -1323 -2752
rect -1515 -2792 -1503 -2758
rect -1335 -2792 -1323 -2758
rect -1515 -2798 -1323 -2792
rect -1257 -2758 -1065 -2752
rect -1257 -2792 -1245 -2758
rect -1077 -2792 -1065 -2758
rect -1257 -2798 -1065 -2792
rect -999 -2758 -807 -2752
rect -999 -2792 -987 -2758
rect -819 -2792 -807 -2758
rect -999 -2798 -807 -2792
rect -741 -2758 -549 -2752
rect -741 -2792 -729 -2758
rect -561 -2792 -549 -2758
rect -741 -2798 -549 -2792
rect -483 -2758 -291 -2752
rect -483 -2792 -471 -2758
rect -303 -2792 -291 -2758
rect -483 -2798 -291 -2792
rect -225 -2758 -33 -2752
rect -225 -2792 -213 -2758
rect -45 -2792 -33 -2758
rect -225 -2798 -33 -2792
rect 33 -2758 225 -2752
rect 33 -2792 45 -2758
rect 213 -2792 225 -2758
rect 33 -2798 225 -2792
rect 291 -2758 483 -2752
rect 291 -2792 303 -2758
rect 471 -2792 483 -2758
rect 291 -2798 483 -2792
rect 549 -2758 741 -2752
rect 549 -2792 561 -2758
rect 729 -2792 741 -2758
rect 549 -2798 741 -2792
rect 807 -2758 999 -2752
rect 807 -2792 819 -2758
rect 987 -2792 999 -2758
rect 807 -2798 999 -2792
rect 1065 -2758 1257 -2752
rect 1065 -2792 1077 -2758
rect 1245 -2792 1257 -2758
rect 1065 -2798 1257 -2792
rect 1323 -2758 1515 -2752
rect 1323 -2792 1335 -2758
rect 1503 -2792 1515 -2758
rect 1323 -2798 1515 -2792
rect 1581 -2758 1773 -2752
rect 1581 -2792 1593 -2758
rect 1761 -2792 1773 -2758
rect 1581 -2798 1773 -2792
rect 1839 -2758 2031 -2752
rect 1839 -2792 1851 -2758
rect 2019 -2792 2031 -2758
rect 1839 -2798 2031 -2792
rect 2097 -2758 2289 -2752
rect 2097 -2792 2109 -2758
rect 2277 -2792 2289 -2758
rect 2097 -2798 2289 -2792
rect 2355 -2758 2547 -2752
rect 2355 -2792 2367 -2758
rect 2535 -2792 2547 -2758
rect 2355 -2798 2547 -2792
rect 2613 -2758 2805 -2752
rect 2613 -2792 2625 -2758
rect 2793 -2792 2805 -2758
rect 2613 -2798 2805 -2792
rect 2871 -2758 3063 -2752
rect 2871 -2792 2883 -2758
rect 3051 -2792 3063 -2758
rect 2871 -2798 3063 -2792
<< properties >>
string FIXED_BBOX -3230 -2913 3230 2913
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 1.0 m 5 nf 24 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
