magic
tech sky130A
magscale 1 2
timestamp 1730992408
<< error_s >>
rect 628 -1154 752 -902
rect 14110 -1154 15010 -658
<< dnwell >>
rect 628 -1154 15010 8321
<< nwell >>
rect 3870 1488 12152 1656
rect 3870 -902 4240 1488
rect 7458 -902 7736 1488
rect 8440 -902 8718 1488
rect 11924 -902 12152 1488
rect 3870 -1104 12152 -902
rect 752 -1154 12152 -1104
<< mvnsubdiff >>
rect 4074 1456 4152 1496
rect 12014 1442 12076 1482
rect 4074 -826 4152 -786
rect 7546 1394 7620 1434
rect 8534 1398 8612 1438
rect 7546 -888 7620 -808
rect 8534 -884 8612 -804
rect 12014 -864 12076 -824
rect 4066 -1030 7510 -1018
rect 4066 -1076 4132 -1030
rect 7486 -1076 7510 -1030
rect 4066 -1088 7510 -1076
rect 8654 -1030 12070 -1018
rect 8654 -1074 8678 -1030
rect 12044 -1074 12070 -1030
rect 8654 -1086 12070 -1074
<< mvnsubdiffcont >>
rect 4074 -786 4152 1456
rect 7546 -808 7620 1394
rect 8534 -804 8612 1398
rect 12014 -824 12076 1442
rect 4132 -1076 7486 -1030
rect 8678 -1074 12044 -1030
<< poly >>
rect 7940 1170 8006 1236
rect 8142 1170 8224 1236
rect 7932 -440 8014 -374
rect 8150 -440 8216 -374
<< locali >>
rect 10532 8282 12396 8286
rect 10532 8240 10550 8282
rect 12380 8240 12396 8282
rect 10532 8228 12396 8240
rect 10534 2430 12434 2460
rect 10534 2358 10558 2430
rect 12414 2358 12434 2430
rect 10534 2352 12434 2358
rect 1884 2166 11362 2196
rect 1884 2094 1918 2166
rect 11194 2094 11362 2166
rect 1884 2062 11362 2094
rect 1884 1718 2004 2062
rect 11238 1718 11362 2062
rect 1884 1688 11362 1718
rect 1884 1616 1922 1688
rect 11194 1616 11362 1688
rect 1884 1584 11362 1616
rect 4060 1456 4170 1502
rect 778 1412 866 1426
rect 3750 1412 3838 1424
rect 778 1396 3838 1412
rect 778 1356 866 1396
rect 3746 1356 3838 1396
rect 778 1338 3838 1356
rect 778 1294 866 1338
rect 778 -904 806 1294
rect 852 -904 866 1294
rect 1138 -798 1254 1192
rect 1416 -798 1532 1192
rect 1694 -798 1810 1192
rect 1972 -798 2088 1192
rect 2250 -798 2366 1192
rect 2528 -798 2644 1192
rect 2806 -798 2922 1192
rect 3084 -798 3200 1192
rect 3362 -798 3478 1192
rect 3750 1182 3838 1338
rect 3750 -790 3768 1182
rect 3814 -790 3838 1182
rect 778 -956 866 -904
rect 3750 -956 3838 -790
rect 778 -974 3838 -956
rect 778 -1014 866 -974
rect 3746 -1014 3838 -974
rect 778 -1028 3838 -1014
rect 832 -1030 3838 -1028
rect 4060 -786 4074 1456
rect 4152 -786 4170 1456
rect 4060 -1012 4170 -786
rect 4288 1412 4352 1444
rect 4288 770 4300 1412
rect 4340 770 4352 1412
rect 4288 734 4352 770
rect 7352 1412 7416 1444
rect 7352 770 7364 1412
rect 7404 770 7416 1412
rect 4288 724 4364 734
rect 7352 732 7416 770
rect 4288 528 4308 724
rect 4346 528 4364 724
rect 4288 520 4364 528
rect 7338 726 7416 732
rect 7338 528 7348 726
rect 7388 528 7416 726
rect 7338 520 7416 528
rect 4288 482 4352 520
rect 4288 -856 4302 482
rect 4342 -812 4352 482
rect 7352 482 7416 520
rect 7352 -812 7364 482
rect 4342 -830 7364 -812
rect 4342 -856 4410 -830
rect 4288 -872 4410 -856
rect 7290 -856 7364 -830
rect 7404 -856 7416 482
rect 7290 -872 7416 -856
rect 4288 -884 7416 -872
rect 7534 1394 7644 1510
rect 7534 -808 7542 1394
rect 7620 -808 7644 1394
rect 7798 1404 8358 1432
rect 7798 1334 7834 1404
rect 8322 1334 8358 1404
rect 7798 1282 8358 1334
rect 8522 1398 8632 1490
rect 8142 1186 8156 1220
rect 8210 1186 8224 1220
rect 7778 428 7828 434
rect 7778 228 7794 428
rect 7778 220 7828 228
rect 7932 -424 7944 -390
rect 8002 -424 8014 -390
rect 7796 -540 8356 -488
rect 7796 -610 7830 -540
rect 8318 -610 8356 -540
rect 7796 -638 8356 -610
rect 7534 -944 7644 -808
rect 8522 -804 8534 1398
rect 8612 -804 8632 1398
rect 8522 -944 8632 -804
rect 8754 1420 8824 1446
rect 8754 1086 8768 1420
rect 8812 1086 8824 1420
rect 8754 1028 8824 1086
rect 8754 828 8778 1028
rect 8818 828 8824 1028
rect 8754 778 8824 828
rect 8754 -812 8768 778
rect 8810 -812 8824 778
rect 11810 1402 11880 1452
rect 11810 1068 11822 1402
rect 11866 1068 11880 1402
rect 11810 1028 11880 1068
rect 11810 830 11818 1028
rect 11858 830 11880 1028
rect 11810 776 11880 830
rect 11810 -812 11822 776
rect 8754 -814 11822 -812
rect 11864 -812 11880 776
rect 11974 1442 12076 1522
rect 11974 1416 12014 1442
rect 11864 -814 11884 -812
rect 8754 -828 11884 -814
rect 8754 -856 8872 -828
rect 8758 -866 8872 -856
rect 11768 -866 11884 -828
rect 8758 -880 11884 -866
rect 11974 -826 11984 1416
rect 12062 -826 12076 -824
rect 7534 -994 8632 -944
rect 11974 -994 12076 -826
rect 7534 -1012 12078 -994
rect 4060 -1018 12078 -1012
rect 4060 -1076 4132 -1018
rect 7506 -1022 12078 -1018
rect 7506 -1038 8674 -1022
rect 7506 -1070 7576 -1038
rect 7486 -1076 7576 -1070
rect 4060 -1088 7576 -1076
rect 8602 -1070 8674 -1038
rect 12058 -1070 12078 -1022
rect 8602 -1074 8678 -1070
rect 12044 -1074 12078 -1070
rect 8602 -1088 12078 -1074
<< viali >>
rect 10550 8240 12380 8282
rect 10533 2509 10567 8177
rect 12348 7074 12384 8042
rect 12692 7946 14878 7980
rect 12348 5964 12384 6932
rect 12348 4856 12384 5824
rect 12348 3748 12384 4716
rect 12348 2634 12384 3602
rect 10558 2358 12414 2430
rect 1918 2094 11194 2166
rect 1922 1616 11194 1688
rect 866 1356 3746 1396
rect 806 -904 852 1294
rect 3768 -790 3814 1182
rect 866 -1014 3746 -974
rect 4074 -786 4152 1456
rect 4300 770 4340 1412
rect 7364 770 7404 1412
rect 4308 528 4346 724
rect 7348 528 7388 726
rect 4302 -856 4342 482
rect 4410 -872 7290 -830
rect 7364 -856 7404 482
rect 7542 -808 7546 1394
rect 7546 -808 7620 1394
rect 7834 1334 8322 1404
rect 8156 1186 8210 1220
rect 7794 228 7830 428
rect 8328 222 8362 434
rect 7944 -424 8002 -390
rect 7830 -610 8318 -540
rect 8534 -804 8612 1398
rect 8768 1086 8812 1420
rect 8778 828 8818 1028
rect 8768 -812 8810 778
rect 11822 1068 11866 1402
rect 11818 830 11858 1028
rect 11822 -814 11864 776
rect 8872 -866 11768 -828
rect 11984 -824 12014 1416
rect 12014 -824 12076 1416
rect 12596 -526 12630 7884
rect 14940 -526 14974 7884
rect 12692 -622 14878 -588
rect 11984 -826 12062 -824
rect 4132 -1030 7506 -1018
rect 4132 -1070 7486 -1030
rect 7486 -1070 7506 -1030
rect 8674 -1030 12058 -1022
rect 8674 -1070 8678 -1030
rect 8678 -1070 12044 -1030
rect 12044 -1070 12058 -1030
<< metal1 >>
rect 10518 8282 12398 8288
rect 10518 8240 10550 8282
rect 12380 8240 12398 8282
rect 10518 8220 10564 8240
rect 12314 8220 12398 8240
rect 10518 8210 12398 8220
rect 10518 8177 10582 8210
rect 10518 2509 10533 8177
rect 10567 2509 10582 8177
rect 12482 8140 12682 8308
rect 10704 8108 12682 8140
rect 10704 8094 12548 8108
rect 10644 8058 10722 8064
rect 10644 7590 10650 8058
rect 10716 7590 10722 8058
rect 10644 7584 10722 7590
rect 11160 8058 11238 8064
rect 11160 7590 11166 8058
rect 11232 7590 11238 8058
rect 11160 7584 11238 7590
rect 11676 8058 11754 8064
rect 11676 7590 11682 8058
rect 11748 7590 11754 8058
rect 11676 7584 11754 7590
rect 12192 8058 12270 8064
rect 12192 7590 12198 8058
rect 12264 7590 12270 8058
rect 12192 7584 12270 7590
rect 12332 8042 12398 8054
rect 10904 7406 10982 7412
rect 10904 7072 10910 7406
rect 10976 7072 10982 7406
rect 10904 7066 10982 7072
rect 11420 7406 11498 7412
rect 11420 7072 11426 7406
rect 11492 7072 11498 7406
rect 11420 7066 11498 7072
rect 11936 7406 12014 7412
rect 11936 7072 11942 7406
rect 12008 7072 12014 7406
rect 11936 7066 12014 7072
rect 12332 7074 12348 8042
rect 12384 7074 12398 8042
rect 12332 7058 12398 7074
rect 12482 7030 12548 8094
rect 14424 7988 14916 8218
rect 10710 6984 12548 7030
rect 10904 6942 10982 6948
rect 10904 6608 10910 6942
rect 10976 6608 10982 6942
rect 10904 6602 10982 6608
rect 11420 6942 11498 6948
rect 11420 6608 11426 6942
rect 11492 6608 11498 6942
rect 11420 6602 11498 6608
rect 11936 6942 12014 6948
rect 11936 6608 11942 6942
rect 12008 6608 12014 6942
rect 11936 6602 12014 6608
rect 12330 6932 12396 6946
rect 10646 6326 10724 6332
rect 10646 5960 10652 6326
rect 10718 5960 10724 6326
rect 10646 5954 10724 5960
rect 11162 6326 11240 6332
rect 11162 5960 11168 6326
rect 11234 5960 11240 6326
rect 11162 5954 11240 5960
rect 11678 6326 11756 6332
rect 11678 5960 11684 6326
rect 11750 5960 11756 6326
rect 11678 5954 11756 5960
rect 12194 6326 12272 6332
rect 12194 5960 12200 6326
rect 12266 5960 12272 6326
rect 12194 5954 12272 5960
rect 12330 5964 12348 6932
rect 12384 5964 12396 6932
rect 12330 5950 12396 5964
rect 12482 5920 12548 6984
rect 10710 5874 12548 5920
rect 12334 5824 12400 5832
rect 10646 5818 10724 5824
rect 10646 5452 10652 5818
rect 10718 5452 10724 5818
rect 10646 5446 10724 5452
rect 11162 5818 11240 5824
rect 11162 5452 11168 5818
rect 11234 5452 11240 5818
rect 11162 5446 11240 5452
rect 11678 5818 11756 5824
rect 11678 5452 11684 5818
rect 11750 5452 11756 5818
rect 11678 5446 11756 5452
rect 12194 5818 12272 5824
rect 12194 5452 12200 5818
rect 12266 5452 12272 5818
rect 12194 5446 12272 5452
rect 10904 5186 10982 5192
rect 10904 4852 10910 5186
rect 10976 4852 10982 5186
rect 10904 4846 10982 4852
rect 11420 5186 11498 5192
rect 11420 4852 11426 5186
rect 11492 4852 11498 5186
rect 11420 4846 11498 4852
rect 11936 5186 12014 5192
rect 11936 4852 11942 5186
rect 12008 4852 12014 5186
rect 11936 4846 12014 4852
rect 12334 4856 12348 5824
rect 12384 4856 12400 5824
rect 12334 4842 12400 4856
rect 12482 4810 12548 5874
rect 10710 4764 12548 4810
rect 10904 4722 10982 4728
rect 10904 4388 10910 4722
rect 10976 4388 10982 4722
rect 10904 4382 10982 4388
rect 11420 4722 11498 4728
rect 11420 4388 11426 4722
rect 11492 4388 11498 4722
rect 11420 4382 11498 4388
rect 11936 4722 12014 4728
rect 11936 4388 11942 4722
rect 12008 4388 12014 4722
rect 11936 4382 12014 4388
rect 12334 4716 12400 4726
rect 10646 4122 10724 4128
rect 10646 3756 10652 4122
rect 10718 3756 10724 4122
rect 10646 3750 10724 3756
rect 11162 4122 11240 4128
rect 11162 3756 11168 4122
rect 11234 3756 11240 4122
rect 11162 3750 11240 3756
rect 11678 4122 11756 4128
rect 11678 3756 11684 4122
rect 11750 3756 11756 4122
rect 11678 3750 11756 3756
rect 12194 4122 12272 4128
rect 12194 3756 12200 4122
rect 12266 3756 12272 4122
rect 12194 3750 12272 3756
rect 12334 3748 12348 4716
rect 12384 3748 12400 4716
rect 12334 3730 12400 3748
rect 12482 3700 12548 4764
rect 10710 3654 12548 3700
rect 10646 3614 10724 3620
rect 10646 3248 10652 3614
rect 10718 3248 10724 3614
rect 10646 3242 10724 3248
rect 11162 3614 11240 3620
rect 11162 3248 11168 3614
rect 11234 3248 11240 3614
rect 11162 3242 11240 3248
rect 11678 3614 11756 3620
rect 11678 3248 11684 3614
rect 11750 3248 11756 3614
rect 11678 3242 11756 3248
rect 12194 3614 12272 3620
rect 12194 3248 12200 3614
rect 12266 3248 12272 3614
rect 12194 3242 12272 3248
rect 12332 3602 12398 3614
rect 10904 2966 10982 2972
rect 10904 2632 10910 2966
rect 10976 2632 10982 2966
rect 10904 2626 10982 2632
rect 11420 2966 11498 2972
rect 11420 2632 11426 2966
rect 11492 2632 11498 2966
rect 11420 2626 11498 2632
rect 11936 2966 12014 2972
rect 11936 2632 11942 2966
rect 12008 2632 12014 2966
rect 11936 2626 12014 2632
rect 12332 2634 12348 3602
rect 12384 2634 12398 3602
rect 12332 2618 12398 2634
rect 12482 2590 12548 3654
rect 10704 2544 12548 2590
rect 10518 2460 10582 2509
rect 10518 2430 12434 2460
rect 10518 2358 10558 2430
rect 12414 2358 12434 2430
rect 10518 2352 12434 2358
rect 1876 2166 11228 2200
rect 1876 2094 1918 2166
rect 11194 2094 11228 2166
rect 1876 2064 11228 2094
rect 11436 2064 11454 2200
rect 1876 2058 11454 2064
rect 1876 1726 2010 2058
rect 11184 2056 11454 2058
rect 10706 1944 11138 1960
rect 10706 1838 10723 1944
rect 11120 1838 11138 1944
rect 10706 1822 11138 1838
rect 11234 1726 11368 2056
rect 1876 1722 11420 1726
rect 1876 1688 11230 1722
rect 1876 1616 1922 1688
rect 11194 1616 11230 1688
rect 1876 1614 11230 1616
rect 11398 1614 11420 1722
rect 1876 1584 11420 1614
rect 4058 1456 4170 1504
rect 778 1422 866 1426
rect 3750 1422 3838 1424
rect 778 1396 3838 1422
rect 778 1356 866 1396
rect 3746 1356 3838 1396
rect 778 1332 3838 1356
rect 778 1294 866 1332
rect 778 -904 806 1294
rect 852 -904 866 1294
rect 1010 1234 3994 1280
rect 916 1128 994 1134
rect 916 472 922 1128
rect 988 472 994 1128
rect 916 466 994 472
rect 1138 -124 1254 1192
rect 1416 1132 1532 1192
rect 1406 1126 1548 1132
rect 1406 472 1412 1126
rect 1542 472 1548 1126
rect 1406 466 1548 472
rect 1128 -130 1270 -124
rect 1128 -784 1134 -130
rect 1264 -784 1270 -130
rect 1128 -790 1270 -784
rect 1138 -798 1254 -790
rect 1416 -798 1532 466
rect 1694 -124 1810 1192
rect 1972 1132 2088 1192
rect 1962 1126 2104 1132
rect 1962 472 1968 1126
rect 2098 472 2104 1126
rect 1962 466 2104 472
rect 1684 -130 1826 -124
rect 1684 -784 1690 -130
rect 1820 -784 1826 -130
rect 1684 -790 1826 -784
rect 1694 -798 1810 -790
rect 1972 -798 2088 466
rect 2250 -124 2366 1192
rect 2528 1132 2644 1192
rect 2518 1126 2660 1132
rect 2518 472 2524 1126
rect 2654 472 2660 1126
rect 2518 466 2660 472
rect 2240 -130 2382 -124
rect 2240 -784 2246 -130
rect 2376 -784 2382 -130
rect 2240 -790 2382 -784
rect 2250 -798 2366 -790
rect 2528 -798 2644 466
rect 2806 -124 2922 1192
rect 3084 1132 3200 1192
rect 3362 1132 3478 1192
rect 3750 1182 3838 1202
rect 3618 1134 3696 1140
rect 3074 1126 3216 1132
rect 3074 472 3080 1126
rect 3210 472 3216 1126
rect 3618 478 3624 1134
rect 3690 478 3696 1134
rect 3618 472 3696 478
rect 3074 466 3216 472
rect 2796 -130 2938 -124
rect 2796 -784 2802 -130
rect 2932 -784 2938 -130
rect 2796 -790 2938 -784
rect 2806 -798 2922 -790
rect 3084 -798 3200 466
rect 3362 -124 3478 466
rect 3352 -130 3494 -124
rect 3352 -784 3358 -130
rect 3488 -784 3494 -130
rect 3352 -790 3494 -784
rect 3750 -790 3768 1182
rect 3814 -790 3838 1182
rect 3919 358 3994 1234
rect 3894 348 3994 358
rect 3894 -18 3904 348
rect 3982 -18 3994 348
rect 3894 -30 3994 -18
rect 3362 -798 3478 -790
rect 3750 -810 3838 -790
rect 3919 -848 3994 -30
rect 1010 -894 3994 -848
rect 4058 -786 4074 1456
rect 4152 -786 4170 1456
rect 4674 1498 7750 1554
rect 4290 1412 4356 1440
rect 4290 770 4300 1412
rect 4340 770 4356 1412
rect 4290 734 4356 770
rect 4402 734 4492 1340
rect 4276 728 4360 734
rect 4276 526 4282 728
rect 4356 526 4360 728
rect 4276 520 4360 526
rect 778 -940 866 -904
rect 778 -974 3838 -940
rect 778 -1014 866 -974
rect 3746 -1014 3838 -974
rect 778 -1028 3838 -1014
rect 832 -1030 3838 -1028
rect 4058 -998 4170 -786
rect 4290 482 4356 520
rect 4290 -856 4302 482
rect 4342 -812 4356 482
rect 4402 -766 4492 520
rect 4674 -780 4726 1498
rect 4902 1034 5068 1340
rect 4902 -766 5068 820
rect 5250 -780 5302 1498
rect 5478 734 5644 1340
rect 5478 -766 5644 520
rect 5826 -780 5878 1498
rect 6054 1034 6220 1340
rect 6054 -766 6220 820
rect 6402 -780 6454 1498
rect 6630 734 6796 1340
rect 6630 -766 6796 520
rect 6978 -780 7030 1498
rect 7352 1412 7418 1440
rect 7206 1034 7296 1340
rect 7206 -766 7296 820
rect 7352 770 7364 1412
rect 7404 770 7418 1412
rect 7352 734 7418 770
rect 7528 1394 7638 1422
rect 7336 726 7430 734
rect 7336 530 7344 726
rect 7424 530 7430 726
rect 7336 528 7348 530
rect 7388 528 7430 530
rect 7336 520 7430 528
rect 7352 482 7418 520
rect 7352 -812 7364 482
rect 4342 -830 7364 -812
rect 4342 -856 4410 -830
rect 4292 -872 4410 -856
rect 7290 -856 7364 -830
rect 7404 -856 7418 482
rect 7290 -872 7418 -856
rect 4292 -884 7418 -872
rect 7528 -808 7542 1394
rect 7620 -808 7638 1394
rect 7528 -998 7638 -808
rect 4058 -1018 7638 -998
rect 4058 -1070 4132 -1018
rect 7506 -1036 7638 -1018
rect 7694 1226 7750 1498
rect 8402 1490 11490 1546
rect 7798 1404 8358 1432
rect 7798 1334 7834 1404
rect 8322 1334 8358 1404
rect 7798 1282 8358 1334
rect 8402 1226 8458 1490
rect 7694 1180 8006 1226
rect 8142 1220 8458 1226
rect 8142 1186 8156 1220
rect 8210 1186 8458 1220
rect 8142 1180 8458 1186
rect 7694 -384 7750 1180
rect 8072 1032 8160 1046
rect 8072 820 8080 1032
rect 8150 820 8160 1032
rect 8072 810 8160 820
rect 7862 734 7950 744
rect 7862 522 7872 734
rect 7942 522 7950 734
rect 7862 508 7950 522
rect 7998 434 8082 442
rect 7778 428 7848 434
rect 7778 228 7786 428
rect 7838 228 7848 428
rect 7778 220 7848 228
rect 7998 222 8004 434
rect 8078 222 8082 434
rect 7998 212 8082 222
rect 8208 434 8374 442
rect 8208 222 8214 434
rect 8288 222 8328 434
rect 8362 222 8374 434
rect 8208 212 8374 222
rect 8402 -384 8458 1180
rect 7694 -390 8014 -384
rect 7694 -424 7944 -390
rect 8002 -424 8014 -390
rect 7694 -430 8014 -424
rect 8150 -430 8458 -384
rect 7694 -884 7750 -430
rect 7796 -540 8356 -488
rect 7796 -610 7830 -540
rect 8318 -610 8356 -540
rect 7796 -638 8356 -610
rect 8402 -884 8458 -430
rect 7506 -1070 7576 -1036
rect 4058 -1086 7576 -1070
rect 7694 -1084 7894 -884
rect 8258 -1084 8458 -884
rect 8520 1398 8630 1428
rect 8520 -804 8534 1398
rect 8612 -804 8630 1398
rect 8756 1420 8822 1442
rect 8756 1086 8768 1420
rect 8812 1086 8822 1420
rect 8756 1034 8822 1086
rect 8870 1034 8958 1362
rect 8738 1030 8832 1034
rect 8738 828 8746 1030
rect 8822 828 8832 1030
rect 8738 820 8832 828
rect 8520 -982 8630 -804
rect 8756 778 8822 820
rect 8756 -812 8768 778
rect 8810 -812 8822 778
rect 8870 -744 8958 820
rect 9134 -764 9186 1490
rect 9368 734 9534 1362
rect 9368 -744 9534 520
rect 9710 -764 9762 1490
rect 9944 1034 10110 1362
rect 9944 -744 10110 820
rect 10286 -764 10338 1490
rect 10520 734 10686 1362
rect 10520 -744 10686 520
rect 10862 -764 10914 1490
rect 11096 1034 11262 1362
rect 11096 -744 11262 820
rect 11438 -764 11490 1490
rect 11810 1402 11876 1446
rect 11672 734 11758 1362
rect 11810 1068 11822 1402
rect 11866 1068 11876 1402
rect 11810 1034 11876 1068
rect 11968 1416 12082 1526
rect 11804 1028 11902 1034
rect 11804 830 11814 1028
rect 11894 830 11902 1028
rect 11804 820 11902 830
rect 11672 -744 11758 520
rect 11810 776 11876 820
rect 11810 -812 11822 776
rect 8756 -814 11822 -812
rect 11864 -812 11876 776
rect 11864 -814 11884 -812
rect 8756 -828 11884 -814
rect 8756 -866 8872 -828
rect 11768 -866 11884 -828
rect 8756 -880 11884 -866
rect 11968 -826 11984 1416
rect 12076 -180 12082 1416
rect 12076 -190 12208 -180
rect 12194 -616 12208 -190
rect 12076 -628 12208 -616
rect 12076 -824 12082 -628
rect 12062 -826 12082 -824
rect 11968 -982 12082 -826
rect 8520 -1018 12082 -982
rect 8520 -1038 8674 -1018
rect 8602 -1070 8674 -1038
rect 12058 -1070 12082 -1018
rect 8602 -1088 12082 -1070
rect 12482 -1085 12548 2544
rect 12590 7980 14981 7988
rect 12590 7946 12692 7980
rect 14878 7946 14981 7980
rect 12590 7938 14981 7946
rect 12590 7884 12636 7938
rect 14932 7884 14981 7938
rect 12590 -526 12596 7884
rect 12630 -526 12636 7884
rect 12794 7838 13128 7884
rect 13586 7838 14904 7884
rect 12670 6338 12770 7792
rect 12670 5960 12680 6338
rect 12670 3758 12770 5960
rect 13734 4080 13834 7792
rect 13734 3798 13834 3808
rect 14792 5844 14892 7792
rect 14792 3788 14892 5482
rect 12670 3602 14822 3758
rect 12666 734 12766 3572
rect 12666 -440 12766 518
rect 13738 3564 13838 3574
rect 13738 -128 13838 3292
rect 13738 -438 13838 -428
rect 14782 1560 14882 3568
rect 14782 -444 14882 1364
rect 12796 -526 13110 -480
rect 13618 -526 14886 -480
rect 14932 -526 14940 7884
rect 14974 -526 14981 7884
rect 12590 -581 12636 -526
rect 14932 -581 14981 -526
rect 12590 -588 14981 -581
rect 12590 -622 12692 -588
rect 14878 -622 14981 -588
rect 12590 -628 14981 -622
rect 12592 -629 14981 -628
rect 12664 -660 14888 -629
rect 12664 -724 12692 -660
rect 14868 -724 14888 -660
rect 12664 -742 14888 -724
<< via1 >>
rect 10564 8240 12314 8278
rect 10564 8220 12314 8240
rect 10650 7590 10716 8058
rect 11166 7590 11232 8058
rect 11682 7590 11748 8058
rect 12198 7590 12264 8058
rect 10910 7072 10976 7406
rect 11426 7072 11492 7406
rect 11942 7072 12008 7406
rect 10910 6608 10976 6942
rect 11426 6608 11492 6942
rect 11942 6608 12008 6942
rect 10652 5960 10718 6326
rect 11168 5960 11234 6326
rect 11684 5960 11750 6326
rect 12200 5960 12266 6326
rect 10652 5452 10718 5818
rect 11168 5452 11234 5818
rect 11684 5452 11750 5818
rect 12200 5452 12266 5818
rect 10910 4852 10976 5186
rect 11426 4852 11492 5186
rect 11942 4852 12008 5186
rect 10910 4388 10976 4722
rect 11426 4388 11492 4722
rect 11942 4388 12008 4722
rect 10652 3756 10718 4122
rect 11168 3756 11234 4122
rect 11684 3756 11750 4122
rect 12200 3756 12266 4122
rect 10652 3248 10718 3614
rect 11168 3248 11234 3614
rect 11684 3248 11750 3614
rect 12200 3248 12266 3614
rect 10910 2632 10976 2966
rect 11426 2632 11492 2966
rect 11942 2632 12008 2966
rect 11228 2064 11436 2200
rect 2126 1840 2516 1942
rect 10723 1838 11120 1944
rect 11230 1614 11398 1722
rect 922 472 988 1128
rect 1412 472 1542 1126
rect 1134 -784 1264 -130
rect 1968 472 2098 1126
rect 1690 -784 1820 -130
rect 2524 472 2654 1126
rect 2246 -784 2376 -130
rect 3080 472 3210 1126
rect 3624 478 3690 1134
rect 2802 -784 2932 -130
rect 3358 -784 3488 -130
rect 3904 -18 3982 348
rect 4282 724 4356 728
rect 4282 528 4308 724
rect 4308 528 4346 724
rect 4346 528 4356 724
rect 4282 526 4356 528
rect 4402 520 4492 734
rect 4902 820 5068 1034
rect 5478 520 5644 734
rect 6054 820 6220 1034
rect 6630 520 6796 734
rect 7206 820 7296 1034
rect 7344 530 7348 726
rect 7348 530 7388 726
rect 7388 530 7424 726
rect 4132 -1070 7506 -1018
rect 8080 820 8150 1032
rect 7872 522 7942 734
rect 7786 228 7794 428
rect 7794 228 7830 428
rect 7830 228 7838 428
rect 8004 222 8078 434
rect 8214 222 8288 434
rect 8746 1028 8822 1030
rect 8746 828 8778 1028
rect 8778 828 8818 1028
rect 8818 828 8822 1028
rect 8870 820 8958 1034
rect 9368 520 9534 734
rect 9944 820 10110 1034
rect 10520 520 10686 734
rect 11096 820 11262 1034
rect 11814 830 11818 1028
rect 11818 830 11858 1028
rect 11858 830 11894 1028
rect 11672 520 11758 734
rect 12006 -616 12076 -190
rect 12076 -616 12194 -190
rect 8674 -1022 12058 -1018
rect 8674 -1070 12058 -1022
rect 12680 5960 12770 6338
rect 13734 3808 13834 4080
rect 14792 5482 14892 5844
rect 12666 518 12766 734
rect 13738 3292 13838 3564
rect 13738 -428 13838 -128
rect 14782 1364 14882 1560
rect 12692 -724 14868 -660
<< metal2 >>
rect 10472 8280 14916 8282
rect 10472 8278 12702 8280
rect 10472 8220 10564 8278
rect 12314 8220 12702 8278
rect 10472 8058 12702 8220
rect 10472 7590 10650 8058
rect 10716 7590 11166 8058
rect 11232 7590 11682 8058
rect 11748 7590 12198 8058
rect 12264 7590 12702 8058
rect 10472 7584 12702 7590
rect 12944 7584 14916 8280
rect 10472 7582 14916 7584
rect 628 7406 11682 7414
rect 628 7398 10910 7406
rect 628 6536 644 7398
rect 824 7072 10910 7398
rect 10976 7072 11426 7406
rect 11492 7072 11682 7406
rect 824 6942 11682 7072
rect 824 6608 10910 6942
rect 10976 6608 11426 6942
rect 11492 6608 11682 6942
rect 824 6536 11682 6608
rect 628 6522 11682 6536
rect 11872 7406 14916 7414
rect 11872 7072 11942 7406
rect 12008 7398 14916 7406
rect 12008 7072 13882 7398
rect 11872 6942 13882 7072
rect 11872 6608 11942 6942
rect 12008 6608 13882 6942
rect 11872 6550 13882 6608
rect 14024 6550 14916 7398
rect 11872 6522 14916 6550
rect 10464 6326 12512 6336
rect 10464 5960 10652 6326
rect 10718 5960 11168 6326
rect 11234 5960 11684 6326
rect 11750 5960 12200 6326
rect 12266 5960 12512 6326
rect 12674 5960 12680 6338
rect 12770 5962 14132 6338
rect 14306 5962 14916 6338
rect 12770 5960 14916 5962
rect 10464 5894 12512 5960
rect 10464 5818 12698 5894
rect 10464 5452 10652 5818
rect 10718 5452 11168 5818
rect 11234 5452 11684 5818
rect 11750 5452 12200 5818
rect 12266 5452 12698 5818
rect 10464 5444 12698 5452
rect 12950 5444 12976 5894
rect 13064 5482 13084 5844
rect 13360 5482 14792 5844
rect 14892 5482 14916 5844
rect 628 5238 11678 5254
rect 628 4376 642 5238
rect 822 5186 11678 5238
rect 822 4852 10910 5186
rect 10976 4852 11426 5186
rect 11492 4852 11678 5186
rect 822 4722 11678 4852
rect 822 4388 10910 4722
rect 10976 4388 11426 4722
rect 11492 4388 11678 4722
rect 822 4376 11678 4388
rect 628 4362 11678 4376
rect 11868 5234 14916 5254
rect 11868 5186 13884 5234
rect 11868 4852 11942 5186
rect 12008 4852 13884 5186
rect 11868 4722 13884 4852
rect 11868 4388 11942 4722
rect 12008 4388 13884 4722
rect 11868 4386 13884 4388
rect 14026 4386 14916 5234
rect 11868 4362 14916 4386
rect 10458 4122 12698 4130
rect 10458 3756 10652 4122
rect 10718 3756 11168 4122
rect 11234 3756 11684 4122
rect 11750 3756 12200 4122
rect 12266 3756 12698 4122
rect 10458 3614 12698 3756
rect 10458 3248 10652 3614
rect 10718 3248 11168 3614
rect 11234 3248 11684 3614
rect 11750 3248 12200 3614
rect 12266 3248 12698 3614
rect 10458 3238 12698 3248
rect 12950 3238 12974 4130
rect 13684 4120 14916 4140
rect 13684 4080 14448 4120
rect 13684 3808 13734 4080
rect 13834 3808 14448 4080
rect 13684 3564 14448 3808
rect 13684 3292 13738 3564
rect 13838 3310 14448 3564
rect 14900 3310 14916 4120
rect 13838 3292 14916 3310
rect 13684 3284 14916 3292
rect 628 3046 11686 3060
rect 628 2384 642 3046
rect 822 2966 11686 3046
rect 822 2632 10910 2966
rect 10976 2632 11426 2966
rect 11492 2632 11686 2966
rect 822 2384 11686 2632
rect 628 2368 11686 2384
rect 11882 3044 14916 3060
rect 11882 2966 13884 3044
rect 11882 2632 11942 2966
rect 12008 2632 13884 2966
rect 11882 2390 13884 2632
rect 14024 2390 14916 3044
rect 11882 2368 14916 2390
rect 11214 2200 12702 2206
rect 11214 2064 11228 2200
rect 11436 2064 12702 2200
rect 11214 2062 12702 2064
rect 12946 2062 12956 2206
rect 13472 2114 13772 2138
rect 13472 2006 13498 2114
rect 628 1994 2572 2004
rect 628 1802 638 1994
rect 828 1942 2572 1994
rect 828 1840 2126 1942
rect 2516 1840 2572 1942
rect 828 1802 2572 1840
rect 628 1790 2572 1802
rect 10668 1944 13498 2006
rect 10668 1838 10723 1944
rect 11120 1838 13498 1944
rect 10668 1808 13498 1838
rect 13750 2006 13772 2114
rect 13750 1808 13774 2006
rect 10668 1778 13774 1808
rect 11218 1614 11230 1722
rect 11398 1614 12702 1722
rect 12946 1614 12958 1722
rect 628 1448 3866 1460
rect 628 468 642 1448
rect 822 1134 3866 1448
rect 822 1128 3624 1134
rect 822 472 922 1128
rect 988 1126 3624 1128
rect 988 472 1412 1126
rect 1542 472 1968 1126
rect 2098 472 2524 1126
rect 2654 472 3080 1126
rect 3210 478 3624 1126
rect 3690 478 3866 1134
rect 7348 1364 14126 1560
rect 14316 1364 14782 1560
rect 14882 1364 14926 1560
rect 7348 1034 7544 1364
rect 4276 820 4902 1034
rect 5068 820 6054 1034
rect 6220 820 7206 1034
rect 7296 822 7544 1034
rect 7656 1032 8870 1034
rect 7296 820 7516 822
rect 7656 820 8080 1032
rect 8150 1030 8870 1032
rect 8150 828 8746 1030
rect 8822 828 8870 1030
rect 8150 820 8870 828
rect 8958 820 9944 1034
rect 10110 820 11096 1034
rect 11262 1028 11994 1034
rect 11262 830 11814 1028
rect 11894 830 11994 1028
rect 11262 820 11994 830
rect 4276 728 4402 734
rect 4276 526 4282 728
rect 4356 526 4402 728
rect 4276 520 4402 526
rect 4492 520 5478 734
rect 5644 520 6630 734
rect 6796 726 7872 734
rect 6796 530 7344 726
rect 7424 530 7872 726
rect 6796 522 7872 530
rect 7942 522 8488 734
rect 6796 520 8488 522
rect 8708 520 9368 734
rect 9534 520 10520 734
rect 10686 520 11672 734
rect 11758 520 12666 734
rect 12071 518 12666 520
rect 12766 518 13084 734
rect 13358 518 14926 734
rect 3210 472 3866 478
rect 822 468 3866 472
rect 628 454 3866 468
rect 4276 428 8004 434
rect 3878 348 3994 358
rect 3878 164 3904 348
rect 3982 176 3994 348
rect 4276 228 7786 428
rect 7838 228 8004 428
rect 4276 222 8004 228
rect 8078 222 8214 434
rect 8288 424 14054 434
rect 8288 230 13882 424
rect 14038 230 14054 424
rect 8288 222 14054 230
rect 4276 220 14054 222
rect 3982 164 4082 176
rect 3878 -26 3892 164
rect 4068 -26 4082 164
rect 3878 -38 4082 -26
rect 712 -128 14916 -114
rect 712 -130 13738 -128
rect 712 -784 1134 -130
rect 1264 -784 1690 -130
rect 1820 -784 2246 -130
rect 2376 -784 2802 -130
rect 2932 -784 3358 -130
rect 3488 -190 13738 -130
rect 3488 -616 12006 -190
rect 12194 -428 13738 -190
rect 13838 -132 14916 -128
rect 13838 -428 14438 -132
rect 12194 -616 14438 -428
rect 3488 -660 14438 -616
rect 3488 -724 12692 -660
rect 3488 -784 14438 -724
rect 712 -1018 14438 -784
rect 712 -1070 4132 -1018
rect 7506 -1070 8674 -1018
rect 12058 -1064 14438 -1018
rect 14896 -1064 14916 -132
rect 12058 -1070 14916 -1064
rect 712 -1084 14916 -1070
rect 4016 -1094 7576 -1084
rect 8602 -1094 12094 -1084
<< via2 >>
rect 12702 7584 12944 8280
rect 644 6536 824 7398
rect 13882 6550 14024 7398
rect 14132 5962 14306 6338
rect 12698 5444 12950 5894
rect 13084 5482 13360 5844
rect 642 4376 822 5238
rect 13884 4386 14026 5234
rect 12698 3238 12950 4130
rect 14448 3310 14900 4120
rect 642 2384 822 3046
rect 13884 2390 14024 3044
rect 12702 2062 12946 2206
rect 638 1802 828 1994
rect 13498 1808 13750 2114
rect 12702 1614 12946 1722
rect 642 468 822 1448
rect 14126 1364 14316 1560
rect 13084 518 13358 734
rect 13882 230 14038 424
rect 3892 -18 3904 164
rect 3904 -18 3982 164
rect 3982 -18 4068 164
rect 3892 -26 4068 -18
rect 14438 -660 14896 -132
rect 14438 -724 14868 -660
rect 14868 -724 14896 -660
rect 14438 -1064 14896 -724
<< metal3 >>
rect 12690 8280 12960 8290
rect 12690 7584 12702 8280
rect 12944 7584 12960 8280
rect 13474 8076 13774 8132
rect 13474 7852 13514 8076
rect 13734 7852 13774 8076
rect 628 7398 840 7456
rect 628 6536 644 7398
rect 824 6536 840 7398
rect 628 5238 840 6536
rect 628 4376 642 5238
rect 822 4376 840 5238
rect 628 3046 840 4376
rect 628 2384 642 3046
rect 822 2384 840 3046
rect 628 1994 840 2384
rect 628 1802 638 1994
rect 828 1802 840 1994
rect 628 1448 840 1802
rect 628 468 642 1448
rect 822 468 840 1448
rect 628 374 840 468
rect 12690 5894 12960 7584
rect 12690 5444 12698 5894
rect 12950 5444 12960 5894
rect 12690 4130 12960 5444
rect 12690 3238 12698 4130
rect 12950 3238 12960 4130
rect 12690 2206 12960 3238
rect 12690 2062 12702 2206
rect 12946 2062 12960 2206
rect 12690 1722 12960 2062
rect 12690 1614 12702 1722
rect 12946 1614 12960 1722
rect 4256 176 4586 178
rect 3878 164 4586 176
rect 3878 -26 3892 164
rect 4068 158 4586 164
rect 4068 -26 4284 158
rect 3878 -38 4284 -26
rect 4256 -94 4284 -38
rect 4562 -94 4586 158
rect 12690 124 12960 1614
rect 13074 6794 13374 7750
rect 13074 6570 13114 6794
rect 13334 6570 13374 6794
rect 13074 5844 13374 6570
rect 13074 5482 13084 5844
rect 13360 5482 13374 5844
rect 13074 4188 13374 5482
rect 13074 3964 13114 4188
rect 13334 3964 13374 4188
rect 13074 1572 13374 3964
rect 13074 1348 13114 1572
rect 13334 1348 13374 1572
rect 13074 734 13374 1348
rect 13074 518 13084 734
rect 13358 518 13374 734
rect 13074 340 13374 518
rect 13474 5464 13774 7852
rect 13474 5240 13514 5464
rect 13734 5240 13774 5464
rect 13474 2856 13774 5240
rect 13474 2632 13514 2856
rect 13734 2632 13774 2856
rect 13474 2114 13774 2632
rect 13474 1808 13498 2114
rect 13750 1808 13774 2114
rect 4256 -126 4586 -94
rect 13474 -636 13774 1808
rect 13870 7398 14050 7762
rect 13870 6550 13882 7398
rect 14024 6550 14050 7398
rect 13870 5234 14050 6550
rect 13870 4386 13884 5234
rect 14026 4386 14050 5234
rect 13870 3044 14050 4386
rect 13870 2390 13884 3044
rect 14024 2390 14050 3044
rect 13870 424 14050 2390
rect 13870 230 13882 424
rect 14038 230 14050 424
rect 13870 204 14050 230
rect 14120 6338 14322 8154
rect 14120 5962 14132 6338
rect 14306 5962 14322 6338
rect 14120 1560 14322 5962
rect 14120 1364 14126 1560
rect 14316 1364 14322 1560
rect 14120 -940 14322 1364
rect 14422 4120 14922 8284
rect 14422 3310 14448 4120
rect 14900 3310 14922 4120
rect 14422 -132 14922 3310
rect 14422 -1064 14438 -132
rect 14896 -1064 14922 -132
rect 14422 -1090 14922 -1064
<< via3 >>
rect 13514 7852 13734 8076
rect 4284 -94 4562 158
rect 13114 6570 13334 6794
rect 13114 3964 13334 4188
rect 13114 1348 13334 1572
rect 13514 5240 13734 5464
rect 13514 2632 13734 2856
<< metal4 >>
rect 13474 8076 13774 8116
rect 13474 8012 13514 8076
rect 12458 7908 13514 8012
rect 13474 7852 13514 7908
rect 13734 7852 13774 8076
rect 13474 7814 13774 7852
rect 13074 6794 13374 6834
rect 13074 6732 13114 6794
rect 12466 6628 13114 6732
rect 13074 6570 13114 6628
rect 13334 6570 13374 6794
rect 13074 6530 13374 6570
rect 13474 5464 13774 5504
rect 13474 5400 13514 5464
rect 12466 5296 13514 5400
rect 13474 5240 13514 5296
rect 13734 5240 13774 5464
rect 13474 5200 13774 5240
rect 13074 4188 13374 4228
rect 13074 4120 13114 4188
rect 12466 4016 13114 4120
rect 13074 3964 13114 4016
rect 13334 3964 13374 4188
rect 13074 3924 13374 3964
rect 13474 2856 13774 2896
rect 13474 2788 13514 2856
rect 12466 2684 13514 2788
rect 13474 2632 13514 2684
rect 13734 2632 13774 2856
rect 13474 2592 13774 2632
rect 13074 1572 13374 1612
rect 13074 1508 13114 1572
rect 12466 1404 13114 1508
rect 13074 1348 13114 1404
rect 13334 1348 13374 1572
rect 13074 1308 13374 1348
rect 4366 178 4468 512
rect 4256 158 4586 178
rect 4256 -94 4284 158
rect 4562 -94 4586 158
rect 4256 -126 4586 -94
use sky130_fd_pr__cap_mim_m3_1_BHK9HY  sky130_fd_pr__cap_mim_m3_1_BHK9HY_0 paramcells
timestamp 1730992408
transform 0 1 6770 1 0 4214
box -3798 -5800 3798 5800
use sky130_fd_pr__nfet_05v0_nvt_FEJX3A  sky130_fd_pr__nfet_05v0_nvt_FEJX3A_0 paramcells
timestamp 1730992408
transform -1 0 10317 0 1 293
box -1580 -1194 1580 1194
use sky130_fd_pr__nfet_g5v0d10v5_7WHXCK  sky130_fd_pr__nfet_g5v0d10v5_7WHXCK_0 paramcells
timestamp 1730992408
transform 1 0 11458 0 1 5343
box -973 -2978 973 2978
use sky130_fd_pr__nfet_01v8_lvt_AJ3MPE  XM2 paramcells
timestamp 1730992408
transform -1 0 8078 0 1 398
box -320 -960 320 960
use sky130_fd_pr__pfet_01v8_lvt_UX3DP3  XM6 paramcells
timestamp 1730992408
transform 1 0 13785 0 1 3679
box -1225 -4337 1225 4337
use sky130_fd_pr__pfet_g5v0d10v5_8UL4MK  XM8 paramcells
timestamp 1730992408
transform 1 0 2311 0 1 193
box -1559 -1297 1559 1297
use sky130_fd_pr__nfet_05v0_nvt_FEJX3A  XM10
timestamp 1730992408
transform 1 0 5849 0 1 293
box -1580 -1194 1580 1194
use sky130_fd_pr__res_high_po_0p69_FJD3D2  XR1 paramcells
timestamp 1730992408
transform 0 1 6622 -1 0 1891
box -235 -4682 235 4682
<< labels >>
flabel metal2 13062 -1020 13262 -820 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal2 13052 8032 13252 8232 0 FreeSans 256 0 0 0 VSS
port 5 nsew
flabel metal1 12482 8108 12682 8308 0 FreeSans 256 0 0 0 VBIAS
port 4 nsew
flabel metal3 628 1502 840 1702 0 FreeSans 256 0 0 0 VOUT
port 1 nsew
flabel metal1 8258 -1084 8458 -884 0 FreeSans 256 0 0 0 VINP
port 3 nsew
flabel metal1 7694 -1084 7894 -884 0 FreeSans 256 0 0 0 VINN
port 2 nsew
<< end >>
