magic
tech sky130A
magscale 1 2
timestamp 1730992408
<< pwell >>
rect -973 -2978 973 2978
<< mvnmos >>
rect -745 1720 -545 2720
rect -487 1720 -287 2720
rect -229 1720 -29 2720
rect 29 1720 229 2720
rect 287 1720 487 2720
rect 545 1720 745 2720
rect -745 610 -545 1610
rect -487 610 -287 1610
rect -229 610 -29 1610
rect 29 610 229 1610
rect 287 610 487 1610
rect 545 610 745 1610
rect -745 -500 -545 500
rect -487 -500 -287 500
rect -229 -500 -29 500
rect 29 -500 229 500
rect 287 -500 487 500
rect 545 -500 745 500
rect -745 -1610 -545 -610
rect -487 -1610 -287 -610
rect -229 -1610 -29 -610
rect 29 -1610 229 -610
rect 287 -1610 487 -610
rect 545 -1610 745 -610
rect -745 -2720 -545 -1720
rect -487 -2720 -287 -1720
rect -229 -2720 -29 -1720
rect 29 -2720 229 -1720
rect 287 -2720 487 -1720
rect 545 -2720 745 -1720
<< mvndiff >>
rect -803 2708 -745 2720
rect -803 1732 -791 2708
rect -757 1732 -745 2708
rect -803 1720 -745 1732
rect -545 2708 -487 2720
rect -545 1732 -533 2708
rect -499 1732 -487 2708
rect -545 1720 -487 1732
rect -287 2708 -229 2720
rect -287 1732 -275 2708
rect -241 1732 -229 2708
rect -287 1720 -229 1732
rect -29 2708 29 2720
rect -29 1732 -17 2708
rect 17 1732 29 2708
rect -29 1720 29 1732
rect 229 2708 287 2720
rect 229 1732 241 2708
rect 275 1732 287 2708
rect 229 1720 287 1732
rect 487 2708 545 2720
rect 487 1732 499 2708
rect 533 1732 545 2708
rect 487 1720 545 1732
rect 745 2708 803 2720
rect 745 1732 757 2708
rect 791 1732 803 2708
rect 745 1720 803 1732
rect -803 1598 -745 1610
rect -803 622 -791 1598
rect -757 622 -745 1598
rect -803 610 -745 622
rect -545 1598 -487 1610
rect -545 622 -533 1598
rect -499 622 -487 1598
rect -545 610 -487 622
rect -287 1598 -229 1610
rect -287 622 -275 1598
rect -241 622 -229 1598
rect -287 610 -229 622
rect -29 1598 29 1610
rect -29 622 -17 1598
rect 17 622 29 1598
rect -29 610 29 622
rect 229 1598 287 1610
rect 229 622 241 1598
rect 275 622 287 1598
rect 229 610 287 622
rect 487 1598 545 1610
rect 487 622 499 1598
rect 533 622 545 1598
rect 487 610 545 622
rect 745 1598 803 1610
rect 745 622 757 1598
rect 791 622 803 1598
rect 745 610 803 622
rect -803 488 -745 500
rect -803 -488 -791 488
rect -757 -488 -745 488
rect -803 -500 -745 -488
rect -545 488 -487 500
rect -545 -488 -533 488
rect -499 -488 -487 488
rect -545 -500 -487 -488
rect -287 488 -229 500
rect -287 -488 -275 488
rect -241 -488 -229 488
rect -287 -500 -229 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 229 488 287 500
rect 229 -488 241 488
rect 275 -488 287 488
rect 229 -500 287 -488
rect 487 488 545 500
rect 487 -488 499 488
rect 533 -488 545 488
rect 487 -500 545 -488
rect 745 488 803 500
rect 745 -488 757 488
rect 791 -488 803 488
rect 745 -500 803 -488
rect -803 -622 -745 -610
rect -803 -1598 -791 -622
rect -757 -1598 -745 -622
rect -803 -1610 -745 -1598
rect -545 -622 -487 -610
rect -545 -1598 -533 -622
rect -499 -1598 -487 -622
rect -545 -1610 -487 -1598
rect -287 -622 -229 -610
rect -287 -1598 -275 -622
rect -241 -1598 -229 -622
rect -287 -1610 -229 -1598
rect -29 -622 29 -610
rect -29 -1598 -17 -622
rect 17 -1598 29 -622
rect -29 -1610 29 -1598
rect 229 -622 287 -610
rect 229 -1598 241 -622
rect 275 -1598 287 -622
rect 229 -1610 287 -1598
rect 487 -622 545 -610
rect 487 -1598 499 -622
rect 533 -1598 545 -622
rect 487 -1610 545 -1598
rect 745 -622 803 -610
rect 745 -1598 757 -622
rect 791 -1598 803 -622
rect 745 -1610 803 -1598
rect -803 -1732 -745 -1720
rect -803 -2708 -791 -1732
rect -757 -2708 -745 -1732
rect -803 -2720 -745 -2708
rect -545 -1732 -487 -1720
rect -545 -2708 -533 -1732
rect -499 -2708 -487 -1732
rect -545 -2720 -487 -2708
rect -287 -1732 -229 -1720
rect -287 -2708 -275 -1732
rect -241 -2708 -229 -1732
rect -287 -2720 -229 -2708
rect -29 -1732 29 -1720
rect -29 -2708 -17 -1732
rect 17 -2708 29 -1732
rect -29 -2720 29 -2708
rect 229 -1732 287 -1720
rect 229 -2708 241 -1732
rect 275 -2708 287 -1732
rect 229 -2720 287 -2708
rect 487 -1732 545 -1720
rect 487 -2708 499 -1732
rect 533 -2708 545 -1732
rect 487 -2720 545 -2708
rect 745 -1732 803 -1720
rect 745 -2708 757 -1732
rect 791 -2708 803 -1732
rect 745 -2720 803 -2708
<< mvndiffc >>
rect -791 1732 -757 2708
rect -533 1732 -499 2708
rect -275 1732 -241 2708
rect -17 1732 17 2708
rect 241 1732 275 2708
rect 499 1732 533 2708
rect 757 1732 791 2708
rect -791 622 -757 1598
rect -533 622 -499 1598
rect -275 622 -241 1598
rect -17 622 17 1598
rect 241 622 275 1598
rect 499 622 533 1598
rect 757 622 791 1598
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect -791 -1598 -757 -622
rect -533 -1598 -499 -622
rect -275 -1598 -241 -622
rect -17 -1598 17 -622
rect 241 -1598 275 -622
rect 499 -1598 533 -622
rect 757 -1598 791 -622
rect -791 -2708 -757 -1732
rect -533 -2708 -499 -1732
rect -275 -2708 -241 -1732
rect -17 -2708 17 -1732
rect 241 -2708 275 -1732
rect 499 -2708 533 -1732
rect 757 -2708 791 -1732
<< mvpsubdiff >>
rect -937 2930 937 2942
rect -937 2896 -829 2930
rect 829 2896 937 2930
rect -937 2884 937 2896
rect -937 2834 -879 2884
rect -937 -2834 -925 2834
rect -891 -2834 -879 2834
rect 879 2834 937 2884
rect -937 -2884 -879 -2834
rect 879 -2834 891 2834
rect 925 -2834 937 2834
rect 879 -2884 937 -2834
rect -937 -2896 937 -2884
rect -937 -2930 -829 -2896
rect 829 -2930 937 -2896
rect -937 -2942 937 -2930
<< mvpsubdiffcont >>
rect -829 2896 829 2930
rect -925 -2834 -891 2834
rect 891 -2834 925 2834
rect -829 -2930 829 -2896
<< poly >>
rect -745 2792 -545 2808
rect -745 2758 -729 2792
rect -561 2758 -545 2792
rect -745 2720 -545 2758
rect -487 2792 -287 2808
rect -487 2758 -471 2792
rect -303 2758 -287 2792
rect -487 2720 -287 2758
rect -229 2792 -29 2808
rect -229 2758 -213 2792
rect -45 2758 -29 2792
rect -229 2720 -29 2758
rect 29 2792 229 2808
rect 29 2758 45 2792
rect 213 2758 229 2792
rect 29 2720 229 2758
rect 287 2792 487 2808
rect 287 2758 303 2792
rect 471 2758 487 2792
rect 287 2720 487 2758
rect 545 2792 745 2808
rect 545 2758 561 2792
rect 729 2758 745 2792
rect 545 2720 745 2758
rect -745 1682 -545 1720
rect -745 1648 -729 1682
rect -561 1648 -545 1682
rect -745 1610 -545 1648
rect -487 1682 -287 1720
rect -487 1648 -471 1682
rect -303 1648 -287 1682
rect -487 1610 -287 1648
rect -229 1682 -29 1720
rect -229 1648 -213 1682
rect -45 1648 -29 1682
rect -229 1610 -29 1648
rect 29 1682 229 1720
rect 29 1648 45 1682
rect 213 1648 229 1682
rect 29 1610 229 1648
rect 287 1682 487 1720
rect 287 1648 303 1682
rect 471 1648 487 1682
rect 287 1610 487 1648
rect 545 1682 745 1720
rect 545 1648 561 1682
rect 729 1648 745 1682
rect 545 1610 745 1648
rect -745 572 -545 610
rect -745 538 -729 572
rect -561 538 -545 572
rect -745 500 -545 538
rect -487 572 -287 610
rect -487 538 -471 572
rect -303 538 -287 572
rect -487 500 -287 538
rect -229 572 -29 610
rect -229 538 -213 572
rect -45 538 -29 572
rect -229 500 -29 538
rect 29 572 229 610
rect 29 538 45 572
rect 213 538 229 572
rect 29 500 229 538
rect 287 572 487 610
rect 287 538 303 572
rect 471 538 487 572
rect 287 500 487 538
rect 545 572 745 610
rect 545 538 561 572
rect 729 538 745 572
rect 545 500 745 538
rect -745 -538 -545 -500
rect -745 -572 -729 -538
rect -561 -572 -545 -538
rect -745 -610 -545 -572
rect -487 -538 -287 -500
rect -487 -572 -471 -538
rect -303 -572 -287 -538
rect -487 -610 -287 -572
rect -229 -538 -29 -500
rect -229 -572 -213 -538
rect -45 -572 -29 -538
rect -229 -610 -29 -572
rect 29 -538 229 -500
rect 29 -572 45 -538
rect 213 -572 229 -538
rect 29 -610 229 -572
rect 287 -538 487 -500
rect 287 -572 303 -538
rect 471 -572 487 -538
rect 287 -610 487 -572
rect 545 -538 745 -500
rect 545 -572 561 -538
rect 729 -572 745 -538
rect 545 -610 745 -572
rect -745 -1648 -545 -1610
rect -745 -1682 -729 -1648
rect -561 -1682 -545 -1648
rect -745 -1720 -545 -1682
rect -487 -1648 -287 -1610
rect -487 -1682 -471 -1648
rect -303 -1682 -287 -1648
rect -487 -1720 -287 -1682
rect -229 -1648 -29 -1610
rect -229 -1682 -213 -1648
rect -45 -1682 -29 -1648
rect -229 -1720 -29 -1682
rect 29 -1648 229 -1610
rect 29 -1682 45 -1648
rect 213 -1682 229 -1648
rect 29 -1720 229 -1682
rect 287 -1648 487 -1610
rect 287 -1682 303 -1648
rect 471 -1682 487 -1648
rect 287 -1720 487 -1682
rect 545 -1648 745 -1610
rect 545 -1682 561 -1648
rect 729 -1682 745 -1648
rect 545 -1720 745 -1682
rect -745 -2758 -545 -2720
rect -745 -2792 -729 -2758
rect -561 -2792 -545 -2758
rect -745 -2808 -545 -2792
rect -487 -2758 -287 -2720
rect -487 -2792 -471 -2758
rect -303 -2792 -287 -2758
rect -487 -2808 -287 -2792
rect -229 -2758 -29 -2720
rect -229 -2792 -213 -2758
rect -45 -2792 -29 -2758
rect -229 -2808 -29 -2792
rect 29 -2758 229 -2720
rect 29 -2792 45 -2758
rect 213 -2792 229 -2758
rect 29 -2808 229 -2792
rect 287 -2758 487 -2720
rect 287 -2792 303 -2758
rect 471 -2792 487 -2758
rect 287 -2808 487 -2792
rect 545 -2758 745 -2720
rect 545 -2792 561 -2758
rect 729 -2792 745 -2758
rect 545 -2808 745 -2792
<< polycont >>
rect -729 2758 -561 2792
rect -471 2758 -303 2792
rect -213 2758 -45 2792
rect 45 2758 213 2792
rect 303 2758 471 2792
rect 561 2758 729 2792
rect -729 1648 -561 1682
rect -471 1648 -303 1682
rect -213 1648 -45 1682
rect 45 1648 213 1682
rect 303 1648 471 1682
rect 561 1648 729 1682
rect -729 538 -561 572
rect -471 538 -303 572
rect -213 538 -45 572
rect 45 538 213 572
rect 303 538 471 572
rect 561 538 729 572
rect -729 -572 -561 -538
rect -471 -572 -303 -538
rect -213 -572 -45 -538
rect 45 -572 213 -538
rect 303 -572 471 -538
rect 561 -572 729 -538
rect -729 -1682 -561 -1648
rect -471 -1682 -303 -1648
rect -213 -1682 -45 -1648
rect 45 -1682 213 -1648
rect 303 -1682 471 -1648
rect 561 -1682 729 -1648
rect -729 -2792 -561 -2758
rect -471 -2792 -303 -2758
rect -213 -2792 -45 -2758
rect 45 -2792 213 -2758
rect 303 -2792 471 -2758
rect 561 -2792 729 -2758
<< locali >>
rect -925 2896 -829 2930
rect 829 2896 925 2930
rect -925 2834 -891 2896
rect 891 2834 925 2896
rect -745 2758 -729 2792
rect -561 2758 -545 2792
rect -487 2758 -471 2792
rect -303 2758 -287 2792
rect -229 2758 -213 2792
rect -45 2758 -29 2792
rect 29 2758 45 2792
rect 213 2758 229 2792
rect 287 2758 303 2792
rect 471 2758 487 2792
rect 545 2758 561 2792
rect 729 2758 745 2792
rect -791 2708 -757 2724
rect -791 1716 -757 1732
rect -533 2708 -499 2724
rect -533 1716 -499 1732
rect -275 2708 -241 2724
rect -275 1716 -241 1732
rect -17 2708 17 2724
rect -17 1716 17 1732
rect 241 2708 275 2724
rect 241 1716 275 1732
rect 499 2708 533 2724
rect 499 1716 533 1732
rect 757 2708 791 2724
rect 757 1716 791 1732
rect -745 1648 -729 1682
rect -561 1648 -545 1682
rect -487 1648 -471 1682
rect -303 1648 -287 1682
rect -229 1648 -213 1682
rect -45 1648 -29 1682
rect 29 1648 45 1682
rect 213 1648 229 1682
rect 287 1648 303 1682
rect 471 1648 487 1682
rect 545 1648 561 1682
rect 729 1648 745 1682
rect -791 1598 -757 1614
rect -791 606 -757 622
rect -533 1598 -499 1614
rect -533 606 -499 622
rect -275 1598 -241 1614
rect -275 606 -241 622
rect -17 1598 17 1614
rect -17 606 17 622
rect 241 1598 275 1614
rect 241 606 275 622
rect 499 1598 533 1614
rect 499 606 533 622
rect 757 1598 791 1614
rect 757 606 791 622
rect -745 538 -729 572
rect -561 538 -545 572
rect -487 538 -471 572
rect -303 538 -287 572
rect -229 538 -213 572
rect -45 538 -29 572
rect 29 538 45 572
rect 213 538 229 572
rect 287 538 303 572
rect 471 538 487 572
rect 545 538 561 572
rect 729 538 745 572
rect -791 488 -757 504
rect -791 -504 -757 -488
rect -533 488 -499 504
rect -533 -504 -499 -488
rect -275 488 -241 504
rect -275 -504 -241 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 241 488 275 504
rect 241 -504 275 -488
rect 499 488 533 504
rect 499 -504 533 -488
rect 757 488 791 504
rect 757 -504 791 -488
rect -745 -572 -729 -538
rect -561 -572 -545 -538
rect -487 -572 -471 -538
rect -303 -572 -287 -538
rect -229 -572 -213 -538
rect -45 -572 -29 -538
rect 29 -572 45 -538
rect 213 -572 229 -538
rect 287 -572 303 -538
rect 471 -572 487 -538
rect 545 -572 561 -538
rect 729 -572 745 -538
rect -791 -622 -757 -606
rect -791 -1614 -757 -1598
rect -533 -622 -499 -606
rect -533 -1614 -499 -1598
rect -275 -622 -241 -606
rect -275 -1614 -241 -1598
rect -17 -622 17 -606
rect -17 -1614 17 -1598
rect 241 -622 275 -606
rect 241 -1614 275 -1598
rect 499 -622 533 -606
rect 499 -1614 533 -1598
rect 757 -622 791 -606
rect 757 -1614 791 -1598
rect -745 -1682 -729 -1648
rect -561 -1682 -545 -1648
rect -487 -1682 -471 -1648
rect -303 -1682 -287 -1648
rect -229 -1682 -213 -1648
rect -45 -1682 -29 -1648
rect 29 -1682 45 -1648
rect 213 -1682 229 -1648
rect 287 -1682 303 -1648
rect 471 -1682 487 -1648
rect 545 -1682 561 -1648
rect 729 -1682 745 -1648
rect -791 -1732 -757 -1716
rect -791 -2724 -757 -2708
rect -533 -1732 -499 -1716
rect -533 -2724 -499 -2708
rect -275 -1732 -241 -1716
rect -275 -2724 -241 -2708
rect -17 -1732 17 -1716
rect -17 -2724 17 -2708
rect 241 -1732 275 -1716
rect 241 -2724 275 -2708
rect 499 -1732 533 -1716
rect 499 -2724 533 -2708
rect 757 -1732 791 -1716
rect 757 -2724 791 -2708
rect -745 -2792 -729 -2758
rect -561 -2792 -545 -2758
rect -487 -2792 -471 -2758
rect -303 -2792 -287 -2758
rect -229 -2792 -213 -2758
rect -45 -2792 -29 -2758
rect 29 -2792 45 -2758
rect 213 -2792 229 -2758
rect 287 -2792 303 -2758
rect 471 -2792 487 -2758
rect 545 -2792 561 -2758
rect 729 -2792 745 -2758
rect -925 -2896 -891 -2834
rect 891 -2896 925 -2834
rect -925 -2930 -829 -2896
rect 829 -2930 925 -2896
<< viali >>
rect -729 2758 -561 2792
rect -471 2758 -303 2792
rect -213 2758 -45 2792
rect 45 2758 213 2792
rect 303 2758 471 2792
rect 561 2758 729 2792
rect -791 1732 -757 2708
rect -533 1732 -499 2708
rect -275 1732 -241 2708
rect -17 1732 17 2708
rect 241 1732 275 2708
rect 499 1732 533 2708
rect 757 1732 791 2708
rect -729 1648 -561 1682
rect -471 1648 -303 1682
rect -213 1648 -45 1682
rect 45 1648 213 1682
rect 303 1648 471 1682
rect 561 1648 729 1682
rect -791 622 -757 1598
rect -533 622 -499 1598
rect -275 622 -241 1598
rect -17 622 17 1598
rect 241 622 275 1598
rect 499 622 533 1598
rect 757 622 791 1598
rect -729 538 -561 572
rect -471 538 -303 572
rect -213 538 -45 572
rect 45 538 213 572
rect 303 538 471 572
rect 561 538 729 572
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect -729 -572 -561 -538
rect -471 -572 -303 -538
rect -213 -572 -45 -538
rect 45 -572 213 -538
rect 303 -572 471 -538
rect 561 -572 729 -538
rect -791 -1598 -757 -622
rect -533 -1598 -499 -622
rect -275 -1598 -241 -622
rect -17 -1598 17 -622
rect 241 -1598 275 -622
rect 499 -1598 533 -622
rect 757 -1598 791 -622
rect -729 -1682 -561 -1648
rect -471 -1682 -303 -1648
rect -213 -1682 -45 -1648
rect 45 -1682 213 -1648
rect 303 -1682 471 -1648
rect 561 -1682 729 -1648
rect -791 -2708 -757 -1732
rect -533 -2708 -499 -1732
rect -275 -2708 -241 -1732
rect -17 -2708 17 -1732
rect 241 -2708 275 -1732
rect 499 -2708 533 -1732
rect 757 -2708 791 -1732
rect -729 -2792 -561 -2758
rect -471 -2792 -303 -2758
rect -213 -2792 -45 -2758
rect 45 -2792 213 -2758
rect 303 -2792 471 -2758
rect 561 -2792 729 -2758
<< metal1 >>
rect -741 2792 -549 2798
rect -741 2758 -729 2792
rect -561 2758 -549 2792
rect -741 2752 -549 2758
rect -483 2792 -291 2798
rect -483 2758 -471 2792
rect -303 2758 -291 2792
rect -483 2752 -291 2758
rect -225 2792 -33 2798
rect -225 2758 -213 2792
rect -45 2758 -33 2792
rect -225 2752 -33 2758
rect 33 2792 225 2798
rect 33 2758 45 2792
rect 213 2758 225 2792
rect 33 2752 225 2758
rect 291 2792 483 2798
rect 291 2758 303 2792
rect 471 2758 483 2792
rect 291 2752 483 2758
rect 549 2792 741 2798
rect 549 2758 561 2792
rect 729 2758 741 2792
rect 549 2752 741 2758
rect -797 2708 -751 2720
rect -797 1732 -791 2708
rect -757 1732 -751 2708
rect -797 1720 -751 1732
rect -539 2708 -493 2720
rect -539 1732 -533 2708
rect -499 1732 -493 2708
rect -539 1720 -493 1732
rect -281 2708 -235 2720
rect -281 1732 -275 2708
rect -241 1732 -235 2708
rect -281 1720 -235 1732
rect -23 2708 23 2720
rect -23 1732 -17 2708
rect 17 1732 23 2708
rect -23 1720 23 1732
rect 235 2708 281 2720
rect 235 1732 241 2708
rect 275 1732 281 2708
rect 235 1720 281 1732
rect 493 2708 539 2720
rect 493 1732 499 2708
rect 533 1732 539 2708
rect 493 1720 539 1732
rect 751 2708 797 2720
rect 751 1732 757 2708
rect 791 1732 797 2708
rect 751 1720 797 1732
rect -741 1682 -549 1688
rect -741 1648 -729 1682
rect -561 1648 -549 1682
rect -741 1642 -549 1648
rect -483 1682 -291 1688
rect -483 1648 -471 1682
rect -303 1648 -291 1682
rect -483 1642 -291 1648
rect -225 1682 -33 1688
rect -225 1648 -213 1682
rect -45 1648 -33 1682
rect -225 1642 -33 1648
rect 33 1682 225 1688
rect 33 1648 45 1682
rect 213 1648 225 1682
rect 33 1642 225 1648
rect 291 1682 483 1688
rect 291 1648 303 1682
rect 471 1648 483 1682
rect 291 1642 483 1648
rect 549 1682 741 1688
rect 549 1648 561 1682
rect 729 1648 741 1682
rect 549 1642 741 1648
rect -797 1598 -751 1610
rect -797 622 -791 1598
rect -757 622 -751 1598
rect -797 610 -751 622
rect -539 1598 -493 1610
rect -539 622 -533 1598
rect -499 622 -493 1598
rect -539 610 -493 622
rect -281 1598 -235 1610
rect -281 622 -275 1598
rect -241 622 -235 1598
rect -281 610 -235 622
rect -23 1598 23 1610
rect -23 622 -17 1598
rect 17 622 23 1598
rect -23 610 23 622
rect 235 1598 281 1610
rect 235 622 241 1598
rect 275 622 281 1598
rect 235 610 281 622
rect 493 1598 539 1610
rect 493 622 499 1598
rect 533 622 539 1598
rect 493 610 539 622
rect 751 1598 797 1610
rect 751 622 757 1598
rect 791 622 797 1598
rect 751 610 797 622
rect -741 572 -549 578
rect -741 538 -729 572
rect -561 538 -549 572
rect -741 532 -549 538
rect -483 572 -291 578
rect -483 538 -471 572
rect -303 538 -291 572
rect -483 532 -291 538
rect -225 572 -33 578
rect -225 538 -213 572
rect -45 538 -33 572
rect -225 532 -33 538
rect 33 572 225 578
rect 33 538 45 572
rect 213 538 225 572
rect 33 532 225 538
rect 291 572 483 578
rect 291 538 303 572
rect 471 538 483 572
rect 291 532 483 538
rect 549 572 741 578
rect 549 538 561 572
rect 729 538 741 572
rect 549 532 741 538
rect -797 488 -751 500
rect -797 -488 -791 488
rect -757 -488 -751 488
rect -797 -500 -751 -488
rect -539 488 -493 500
rect -539 -488 -533 488
rect -499 -488 -493 488
rect -539 -500 -493 -488
rect -281 488 -235 500
rect -281 -488 -275 488
rect -241 -488 -235 488
rect -281 -500 -235 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 235 488 281 500
rect 235 -488 241 488
rect 275 -488 281 488
rect 235 -500 281 -488
rect 493 488 539 500
rect 493 -488 499 488
rect 533 -488 539 488
rect 493 -500 539 -488
rect 751 488 797 500
rect 751 -488 757 488
rect 791 -488 797 488
rect 751 -500 797 -488
rect -741 -538 -549 -532
rect -741 -572 -729 -538
rect -561 -572 -549 -538
rect -741 -578 -549 -572
rect -483 -538 -291 -532
rect -483 -572 -471 -538
rect -303 -572 -291 -538
rect -483 -578 -291 -572
rect -225 -538 -33 -532
rect -225 -572 -213 -538
rect -45 -572 -33 -538
rect -225 -578 -33 -572
rect 33 -538 225 -532
rect 33 -572 45 -538
rect 213 -572 225 -538
rect 33 -578 225 -572
rect 291 -538 483 -532
rect 291 -572 303 -538
rect 471 -572 483 -538
rect 291 -578 483 -572
rect 549 -538 741 -532
rect 549 -572 561 -538
rect 729 -572 741 -538
rect 549 -578 741 -572
rect -797 -622 -751 -610
rect -797 -1598 -791 -622
rect -757 -1598 -751 -622
rect -797 -1610 -751 -1598
rect -539 -622 -493 -610
rect -539 -1598 -533 -622
rect -499 -1598 -493 -622
rect -539 -1610 -493 -1598
rect -281 -622 -235 -610
rect -281 -1598 -275 -622
rect -241 -1598 -235 -622
rect -281 -1610 -235 -1598
rect -23 -622 23 -610
rect -23 -1598 -17 -622
rect 17 -1598 23 -622
rect -23 -1610 23 -1598
rect 235 -622 281 -610
rect 235 -1598 241 -622
rect 275 -1598 281 -622
rect 235 -1610 281 -1598
rect 493 -622 539 -610
rect 493 -1598 499 -622
rect 533 -1598 539 -622
rect 493 -1610 539 -1598
rect 751 -622 797 -610
rect 751 -1598 757 -622
rect 791 -1598 797 -622
rect 751 -1610 797 -1598
rect -741 -1648 -549 -1642
rect -741 -1682 -729 -1648
rect -561 -1682 -549 -1648
rect -741 -1688 -549 -1682
rect -483 -1648 -291 -1642
rect -483 -1682 -471 -1648
rect -303 -1682 -291 -1648
rect -483 -1688 -291 -1682
rect -225 -1648 -33 -1642
rect -225 -1682 -213 -1648
rect -45 -1682 -33 -1648
rect -225 -1688 -33 -1682
rect 33 -1648 225 -1642
rect 33 -1682 45 -1648
rect 213 -1682 225 -1648
rect 33 -1688 225 -1682
rect 291 -1648 483 -1642
rect 291 -1682 303 -1648
rect 471 -1682 483 -1648
rect 291 -1688 483 -1682
rect 549 -1648 741 -1642
rect 549 -1682 561 -1648
rect 729 -1682 741 -1648
rect 549 -1688 741 -1682
rect -797 -1732 -751 -1720
rect -797 -2708 -791 -1732
rect -757 -2708 -751 -1732
rect -797 -2720 -751 -2708
rect -539 -1732 -493 -1720
rect -539 -2708 -533 -1732
rect -499 -2708 -493 -1732
rect -539 -2720 -493 -2708
rect -281 -1732 -235 -1720
rect -281 -2708 -275 -1732
rect -241 -2708 -235 -1732
rect -281 -2720 -235 -2708
rect -23 -1732 23 -1720
rect -23 -2708 -17 -1732
rect 17 -2708 23 -1732
rect -23 -2720 23 -2708
rect 235 -1732 281 -1720
rect 235 -2708 241 -1732
rect 275 -2708 281 -1732
rect 235 -2720 281 -2708
rect 493 -1732 539 -1720
rect 493 -2708 499 -1732
rect 533 -2708 539 -1732
rect 493 -2720 539 -2708
rect 751 -1732 797 -1720
rect 751 -2708 757 -1732
rect 791 -2708 797 -1732
rect 751 -2720 797 -2708
rect -741 -2758 -549 -2752
rect -741 -2792 -729 -2758
rect -561 -2792 -549 -2758
rect -741 -2798 -549 -2792
rect -483 -2758 -291 -2752
rect -483 -2792 -471 -2758
rect -303 -2792 -291 -2758
rect -483 -2798 -291 -2792
rect -225 -2758 -33 -2752
rect -225 -2792 -213 -2758
rect -45 -2792 -33 -2758
rect -225 -2798 -33 -2792
rect 33 -2758 225 -2752
rect 33 -2792 45 -2758
rect 213 -2792 225 -2758
rect 33 -2798 225 -2792
rect 291 -2758 483 -2752
rect 291 -2792 303 -2758
rect 471 -2792 483 -2758
rect 291 -2798 483 -2792
rect 549 -2758 741 -2752
rect 549 -2792 561 -2758
rect 729 -2792 741 -2758
rect 549 -2798 741 -2792
<< properties >>
string FIXED_BBOX -908 -2913 908 2913
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 1.0 m 5 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
