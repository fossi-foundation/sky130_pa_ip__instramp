magic
tech sky130A
magscale 1 2
timestamp 1730743893
<< poly >>
rect 8200 970 8484 1036
rect 8192 -640 8476 -574
<< locali >>
rect 766 2264 12420 2436
rect 1880 2062 11362 2196
rect 1880 1718 2004 2062
rect 11238 1718 11362 2062
rect 1880 1584 11362 1718
rect 4532 1202 12066 1358
rect 1138 -798 1254 1192
rect 1416 -798 1532 1192
rect 1694 -798 1810 1192
rect 1972 -798 2088 1192
rect 2250 -798 2366 1192
rect 2528 -798 2644 1192
rect 2806 -798 2922 1192
rect 3084 -798 3200 1192
rect 3362 -798 3478 1192
rect 7592 1102 9024 1202
<< metal1 >>
rect 12482 8140 12682 8308
rect 944 8108 12682 8140
rect 944 8094 12548 8108
rect 12482 7030 12548 8094
rect 13198 7894 13514 7906
rect 13198 7884 13216 7894
rect 12794 7838 13216 7884
rect 13494 7884 13514 7894
rect 13494 7838 14844 7884
rect 944 6984 12548 7030
rect 12482 5920 12548 6984
rect 944 5874 12548 5920
rect 12482 4810 12548 5874
rect 944 4764 12548 4810
rect 12482 3700 12548 4764
rect 944 3654 12548 3700
rect 12482 2590 12548 3654
rect 12806 3750 14848 3754
rect 12806 3608 13212 3750
rect 13500 3608 14848 3750
rect 944 2544 12548 2590
rect 10706 1944 11138 1960
rect 10706 1838 10723 1944
rect 11120 1838 11138 1944
rect 10706 1822 11138 1838
rect 1010 1234 3612 1280
rect 1138 -798 1254 1192
rect 1416 -798 1532 1192
rect 1694 -798 1810 1192
rect 1972 -798 2088 1192
rect 2250 -798 2366 1192
rect 2528 -798 2644 1192
rect 2806 -798 2922 1192
rect 3084 -798 3200 1192
rect 3362 -798 3478 1192
rect 4716 1040 7420 1086
rect 9184 1060 11888 1106
rect 4602 808 4710 1008
rect 5122 808 5286 1008
rect 5698 808 5862 1008
rect 6274 808 6438 1008
rect 6850 808 7014 1008
rect 7426 808 7546 1008
rect 8200 980 8484 1026
rect 9070 828 9178 1028
rect 9590 828 9754 1028
rect 10166 828 10330 1028
rect 10742 828 10906 1028
rect 11318 828 11482 1028
rect 11894 828 12014 1028
rect 4716 730 7420 776
rect 9184 750 11888 796
rect 4716 622 7420 668
rect 9184 642 11888 688
rect 4602 390 4710 590
rect 5122 390 5286 590
rect 5698 390 5862 590
rect 6274 390 6438 590
rect 6850 390 7014 590
rect 7426 390 7546 590
rect 9070 410 9178 610
rect 9590 410 9754 610
rect 10166 410 10330 610
rect 10742 410 10906 610
rect 11318 410 11482 610
rect 11894 410 12014 610
rect 4716 312 7420 358
rect 9184 332 11888 378
rect 4716 204 7420 250
rect 9184 224 11888 270
rect 4602 -28 4710 172
rect 5122 -28 5286 172
rect 5698 -28 5862 172
rect 6274 -28 6438 172
rect 6850 -28 7014 172
rect 7426 -28 7546 172
rect 9070 -8 9178 192
rect 9590 -8 9754 192
rect 10166 -8 10330 192
rect 10742 -8 10906 192
rect 11318 -8 11482 192
rect 11894 -8 12014 192
rect 4716 -106 7420 -60
rect 9184 -86 11888 -40
rect 4716 -214 7420 -168
rect 9184 -194 11888 -148
rect 4602 -446 4710 -246
rect 5122 -446 5286 -246
rect 5698 -446 5862 -246
rect 6274 -446 6438 -246
rect 6850 -446 7014 -246
rect 7426 -446 7546 -246
rect 9070 -426 9178 -226
rect 9590 -426 9754 -226
rect 10166 -426 10330 -226
rect 10742 -426 10906 -226
rect 11318 -426 11482 -226
rect 11894 -426 12014 -226
rect 4716 -524 7420 -478
rect 9184 -504 11888 -458
rect 12796 -486 14846 -480
rect 12796 -526 13218 -486
rect 13198 -542 13218 -526
rect 13496 -526 14846 -486
rect 13496 -542 13514 -526
rect 4716 -632 7420 -586
rect 8192 -630 8476 -584
rect 9184 -612 11888 -566
rect 1010 -894 3612 -848
rect 4602 -864 4710 -664
rect 5122 -864 5286 -664
rect 5698 -864 5862 -664
rect 6274 -864 6438 -664
rect 6850 -864 7014 -664
rect 7426 -864 7546 -664
rect 9070 -844 9178 -644
rect 9590 -844 9754 -644
rect 10166 -844 10330 -644
rect 10742 -844 10906 -644
rect 11318 -844 11482 -644
rect 11894 -844 12014 -644
rect 4716 -942 7420 -896
rect 7846 -1084 8046 -884
rect 8590 -1092 8790 -892
rect 9184 -922 11888 -876
<< via1 >>
rect 13216 7838 13494 7894
rect 13212 3608 13500 3750
rect 2126 1840 2516 1942
rect 10723 1838 11120 1944
rect 13218 -542 13496 -486
<< metal2 >>
rect 724 7936 15018 8282
rect 724 7610 13148 7936
rect 13206 7896 13506 7906
rect 13206 7660 13216 7896
rect 13494 7660 13506 7896
rect 13206 7650 13506 7660
rect 13568 7610 15018 7936
rect 724 7582 15018 7610
rect 628 7398 14916 7414
rect 628 6536 644 7398
rect 824 6536 14916 7398
rect 628 6522 14916 6536
rect 912 5444 12512 6336
rect 12714 5482 15008 6338
rect 628 5238 14900 5254
rect 628 4376 642 5238
rect 822 4376 14900 5238
rect 628 4362 14900 4376
rect 882 3268 12420 4160
rect 12730 3820 15024 4140
rect 12730 3528 13122 3820
rect 13194 3582 13212 3780
rect 13500 3582 13518 3780
rect 13594 3528 15024 3820
rect 12730 3284 15024 3528
rect 628 3046 14906 3060
rect 628 2384 642 3046
rect 822 2384 14906 3046
rect 628 2368 14906 2384
rect 12704 2114 13004 2138
rect 628 2074 2572 2084
rect 628 1894 640 2074
rect 828 1942 2572 2074
rect 12704 2006 12730 2114
rect 828 1894 2126 1942
rect 628 1880 2126 1894
rect 2074 1840 2126 1880
rect 2516 1840 2572 1942
rect 2074 1790 2572 1840
rect 10668 1944 12730 2006
rect 10668 1838 10723 1944
rect 11120 1838 12730 1944
rect 10668 1808 12730 1838
rect 12982 2006 13004 2114
rect 12982 1808 13006 2006
rect 10668 1778 13006 1808
rect 13140 1684 15016 2140
rect 628 1448 3866 1460
rect 628 468 642 1448
rect 822 468 3866 1448
rect 12722 1284 15016 1684
rect 4350 620 12222 834
rect 628 454 3866 468
rect 4350 320 12222 534
rect 4350 20 12222 234
rect 12600 222 14894 1078
rect 12616 -114 15006 -6
rect 712 -248 15006 -114
rect 712 -574 13148 -248
rect 13206 -296 13506 -284
rect 13206 -542 13218 -296
rect 13496 -542 13506 -296
rect 13206 -546 13506 -542
rect 13562 -574 15006 -248
rect 712 -1084 15006 -574
<< via2 >>
rect 13216 7894 13494 7896
rect 13216 7838 13494 7894
rect 13216 7660 13494 7838
rect 644 6536 824 7398
rect 642 4376 822 5238
rect 13212 3750 13500 3780
rect 13212 3608 13500 3750
rect 13212 3582 13500 3608
rect 642 2384 822 3046
rect 640 1894 828 2074
rect 12730 1808 12982 2114
rect 642 468 822 1448
rect 13218 -486 13496 -296
rect 13218 -532 13496 -486
<< metal3 >>
rect 13206 7896 13506 7906
rect 628 7398 840 7456
rect 628 6536 644 7398
rect 824 6536 840 7398
rect 628 5238 840 6536
rect 628 4376 642 5238
rect 822 4376 840 5238
rect 628 3046 840 4376
rect 628 2384 642 3046
rect 822 2384 840 3046
rect 628 2074 840 2384
rect 628 1894 640 2074
rect 828 1894 840 2074
rect 628 1448 840 1894
rect 628 468 642 1448
rect 822 468 840 1448
rect 628 374 840 468
rect 12706 5516 13006 7750
rect 12706 5292 12746 5516
rect 12966 5292 13006 5516
rect 12706 2908 13006 5292
rect 12706 2684 12746 2908
rect 12966 2684 13006 2908
rect 12706 2114 13006 2684
rect 12706 1808 12730 2114
rect 12982 1808 13006 2114
rect 12706 300 13006 1808
rect 12706 76 12746 300
rect 12966 76 13006 300
rect 12706 36 13006 76
rect 13206 7660 13216 7896
rect 13494 7660 13506 7896
rect 13206 6794 13506 7660
rect 13206 6570 13246 6794
rect 13466 6570 13506 6794
rect 13206 4188 13506 6570
rect 13206 3964 13246 4188
rect 13466 3964 13506 4188
rect 13206 3780 13506 3964
rect 13206 3582 13212 3780
rect 13500 3582 13506 3780
rect 13206 1572 13506 3582
rect 13206 1348 13246 1572
rect 13466 1348 13506 1572
rect 13206 -296 13506 1348
rect 13206 -532 13218 -296
rect 13496 -532 13506 -296
rect 13206 -546 13506 -532
rect 13722 -1090 14222 8284
rect 14422 -1090 14922 8284
<< via3 >>
rect 12746 5292 12966 5516
rect 12746 2684 12966 2908
rect 12746 76 12966 300
rect 13246 6570 13466 6794
rect 13246 3964 13466 4188
rect 13246 1348 13466 1572
<< metal4 >>
rect 13206 6794 13506 6834
rect 13206 6732 13246 6794
rect 12466 6628 13246 6732
rect 13206 6570 13246 6628
rect 13466 6570 13506 6794
rect 13206 6530 13506 6570
rect 12706 5516 13006 5556
rect 12706 5452 12746 5516
rect 1040 5348 1074 5452
rect 12466 5348 12746 5452
rect 12706 5292 12746 5348
rect 12966 5292 13006 5516
rect 12706 5252 13006 5292
rect 13206 4188 13506 4228
rect 13206 4120 13246 4188
rect 12466 4016 13246 4120
rect 13206 3964 13246 4016
rect 13466 3964 13506 4188
rect 13206 3924 13506 3964
rect 12706 2908 13006 2948
rect 12706 2840 12746 2908
rect 1040 2736 1074 2840
rect 12466 2736 12746 2840
rect 12706 2684 12746 2736
rect 12966 2684 13006 2908
rect 12706 2644 13006 2684
rect 13206 1572 13506 1612
rect 13206 1508 13246 1572
rect 12466 1404 13246 1508
rect 13206 1348 13246 1404
rect 13466 1348 13506 1572
rect 13206 1308 13506 1348
rect 12706 300 13006 340
rect 12706 228 12746 300
rect 1040 124 1074 228
rect 12464 124 12746 228
rect 12706 76 12746 124
rect 12966 76 13006 300
rect 12706 36 13006 76
use sky130_fd_pr__cap_mim_m3_1_BHK9HY  XC1 paramcells
timestamp 1730739923
transform 0 1 6770 -1 0 3922
box -3798 -5800 3798 5800
use sky130_fd_pr__nfet_01v8_lvt_AJ3MPE  XM2
timestamp 1730739923
transform -1 0 8338 0 1 198
box -320 -960 320 960
use sky130_fd_pr__nfet_g5v0d10v5_3WU84W  XM5
timestamp 1730737834
transform 1 0 6587 0 1 5342
box -5875 -2978 5875 2978
use sky130_fd_pr__pfet_01v8_lvt_UX3DP3  XM6
timestamp 1730737834
transform 1 0 13819 0 1 3679
box -1225 -4337 1225 4337
use sky130_fd_pr__pfet_g5v0d10v5_8UL4MK  XM8 paramcells
timestamp 1729620069
transform 1 0 2311 0 1 193
box -1559 -1297 1559 1297
use sky130_fd_pr__nfet_05v0_nvt_RLJRR9  XM10 paramcells
timestamp 1730739923
transform 1 0 6068 0 1 72
box -1580 -1194 1580 1194
use sky130_fd_pr__nfet_05v0_nvt_RLJRR9  XM12
timestamp 1730739923
transform -1 0 10536 0 1 92
box -1580 -1194 1580 1194
use sky130_fd_pr__res_high_po_0p69_FJD3D2  XR1 paramcells
timestamp 1730739923
transform 0 1 6622 -1 0 1891
box -235 -4682 235 4682
<< labels >>
flabel metal1 7846 -1084 8046 -884 0 FreeSans 256 0 0 0 VINN
port 2 nsew
flabel metal1 8590 -1092 8790 -892 0 FreeSans 256 0 0 0 VINP
port 3 nsew
flabel metal3 628 1602 840 1802 0 FreeSans 256 0 0 0 VOUT
port 1 nsew
flabel metal2 13062 -1020 13262 -820 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal2 13052 8032 13252 8232 0 FreeSans 256 0 0 0 VSS
port 5 nsew
flabel metal1 12482 8108 12682 8308 0 FreeSans 256 0 0 0 VBIAS
port 4 nsew
<< end >>
