magic
tech sky130A
magscale 1 2
timestamp 1730992408
<< pwell >>
rect -1580 -1194 1580 1194
<< mvnnmos >>
rect -1352 736 -952 936
rect -776 736 -376 936
rect -200 736 200 936
rect 376 736 776 936
rect 952 736 1352 936
rect -1352 318 -952 518
rect -776 318 -376 518
rect -200 318 200 518
rect 376 318 776 518
rect 952 318 1352 518
rect -1352 -100 -952 100
rect -776 -100 -376 100
rect -200 -100 200 100
rect 376 -100 776 100
rect 952 -100 1352 100
rect -1352 -518 -952 -318
rect -776 -518 -376 -318
rect -200 -518 200 -318
rect 376 -518 776 -318
rect 952 -518 1352 -318
rect -1352 -936 -952 -736
rect -776 -936 -376 -736
rect -200 -936 200 -736
rect 376 -936 776 -736
rect 952 -936 1352 -736
<< mvndiff >>
rect -1410 924 -1352 936
rect -1410 748 -1398 924
rect -1364 748 -1352 924
rect -1410 736 -1352 748
rect -952 924 -894 936
rect -952 748 -940 924
rect -906 748 -894 924
rect -952 736 -894 748
rect -834 924 -776 936
rect -834 748 -822 924
rect -788 748 -776 924
rect -834 736 -776 748
rect -376 924 -318 936
rect -376 748 -364 924
rect -330 748 -318 924
rect -376 736 -318 748
rect -258 924 -200 936
rect -258 748 -246 924
rect -212 748 -200 924
rect -258 736 -200 748
rect 200 924 258 936
rect 200 748 212 924
rect 246 748 258 924
rect 200 736 258 748
rect 318 924 376 936
rect 318 748 330 924
rect 364 748 376 924
rect 318 736 376 748
rect 776 924 834 936
rect 776 748 788 924
rect 822 748 834 924
rect 776 736 834 748
rect 894 924 952 936
rect 894 748 906 924
rect 940 748 952 924
rect 894 736 952 748
rect 1352 924 1410 936
rect 1352 748 1364 924
rect 1398 748 1410 924
rect 1352 736 1410 748
rect -1410 506 -1352 518
rect -1410 330 -1398 506
rect -1364 330 -1352 506
rect -1410 318 -1352 330
rect -952 506 -894 518
rect -952 330 -940 506
rect -906 330 -894 506
rect -952 318 -894 330
rect -834 506 -776 518
rect -834 330 -822 506
rect -788 330 -776 506
rect -834 318 -776 330
rect -376 506 -318 518
rect -376 330 -364 506
rect -330 330 -318 506
rect -376 318 -318 330
rect -258 506 -200 518
rect -258 330 -246 506
rect -212 330 -200 506
rect -258 318 -200 330
rect 200 506 258 518
rect 200 330 212 506
rect 246 330 258 506
rect 200 318 258 330
rect 318 506 376 518
rect 318 330 330 506
rect 364 330 376 506
rect 318 318 376 330
rect 776 506 834 518
rect 776 330 788 506
rect 822 330 834 506
rect 776 318 834 330
rect 894 506 952 518
rect 894 330 906 506
rect 940 330 952 506
rect 894 318 952 330
rect 1352 506 1410 518
rect 1352 330 1364 506
rect 1398 330 1410 506
rect 1352 318 1410 330
rect -1410 88 -1352 100
rect -1410 -88 -1398 88
rect -1364 -88 -1352 88
rect -1410 -100 -1352 -88
rect -952 88 -894 100
rect -952 -88 -940 88
rect -906 -88 -894 88
rect -952 -100 -894 -88
rect -834 88 -776 100
rect -834 -88 -822 88
rect -788 -88 -776 88
rect -834 -100 -776 -88
rect -376 88 -318 100
rect -376 -88 -364 88
rect -330 -88 -318 88
rect -376 -100 -318 -88
rect -258 88 -200 100
rect -258 -88 -246 88
rect -212 -88 -200 88
rect -258 -100 -200 -88
rect 200 88 258 100
rect 200 -88 212 88
rect 246 -88 258 88
rect 200 -100 258 -88
rect 318 88 376 100
rect 318 -88 330 88
rect 364 -88 376 88
rect 318 -100 376 -88
rect 776 88 834 100
rect 776 -88 788 88
rect 822 -88 834 88
rect 776 -100 834 -88
rect 894 88 952 100
rect 894 -88 906 88
rect 940 -88 952 88
rect 894 -100 952 -88
rect 1352 88 1410 100
rect 1352 -88 1364 88
rect 1398 -88 1410 88
rect 1352 -100 1410 -88
rect -1410 -330 -1352 -318
rect -1410 -506 -1398 -330
rect -1364 -506 -1352 -330
rect -1410 -518 -1352 -506
rect -952 -330 -894 -318
rect -952 -506 -940 -330
rect -906 -506 -894 -330
rect -952 -518 -894 -506
rect -834 -330 -776 -318
rect -834 -506 -822 -330
rect -788 -506 -776 -330
rect -834 -518 -776 -506
rect -376 -330 -318 -318
rect -376 -506 -364 -330
rect -330 -506 -318 -330
rect -376 -518 -318 -506
rect -258 -330 -200 -318
rect -258 -506 -246 -330
rect -212 -506 -200 -330
rect -258 -518 -200 -506
rect 200 -330 258 -318
rect 200 -506 212 -330
rect 246 -506 258 -330
rect 200 -518 258 -506
rect 318 -330 376 -318
rect 318 -506 330 -330
rect 364 -506 376 -330
rect 318 -518 376 -506
rect 776 -330 834 -318
rect 776 -506 788 -330
rect 822 -506 834 -330
rect 776 -518 834 -506
rect 894 -330 952 -318
rect 894 -506 906 -330
rect 940 -506 952 -330
rect 894 -518 952 -506
rect 1352 -330 1410 -318
rect 1352 -506 1364 -330
rect 1398 -506 1410 -330
rect 1352 -518 1410 -506
rect -1410 -748 -1352 -736
rect -1410 -924 -1398 -748
rect -1364 -924 -1352 -748
rect -1410 -936 -1352 -924
rect -952 -748 -894 -736
rect -952 -924 -940 -748
rect -906 -924 -894 -748
rect -952 -936 -894 -924
rect -834 -748 -776 -736
rect -834 -924 -822 -748
rect -788 -924 -776 -748
rect -834 -936 -776 -924
rect -376 -748 -318 -736
rect -376 -924 -364 -748
rect -330 -924 -318 -748
rect -376 -936 -318 -924
rect -258 -748 -200 -736
rect -258 -924 -246 -748
rect -212 -924 -200 -748
rect -258 -936 -200 -924
rect 200 -748 258 -736
rect 200 -924 212 -748
rect 246 -924 258 -748
rect 200 -936 258 -924
rect 318 -748 376 -736
rect 318 -924 330 -748
rect 364 -924 376 -748
rect 318 -936 376 -924
rect 776 -748 834 -736
rect 776 -924 788 -748
rect 822 -924 834 -748
rect 776 -936 834 -924
rect 894 -748 952 -736
rect 894 -924 906 -748
rect 940 -924 952 -748
rect 894 -936 952 -924
rect 1352 -748 1410 -736
rect 1352 -924 1364 -748
rect 1398 -924 1410 -748
rect 1352 -936 1410 -924
<< mvndiffc >>
rect -1398 748 -1364 924
rect -940 748 -906 924
rect -822 748 -788 924
rect -364 748 -330 924
rect -246 748 -212 924
rect 212 748 246 924
rect 330 748 364 924
rect 788 748 822 924
rect 906 748 940 924
rect 1364 748 1398 924
rect -1398 330 -1364 506
rect -940 330 -906 506
rect -822 330 -788 506
rect -364 330 -330 506
rect -246 330 -212 506
rect 212 330 246 506
rect 330 330 364 506
rect 788 330 822 506
rect 906 330 940 506
rect 1364 330 1398 506
rect -1398 -88 -1364 88
rect -940 -88 -906 88
rect -822 -88 -788 88
rect -364 -88 -330 88
rect -246 -88 -212 88
rect 212 -88 246 88
rect 330 -88 364 88
rect 788 -88 822 88
rect 906 -88 940 88
rect 1364 -88 1398 88
rect -1398 -506 -1364 -330
rect -940 -506 -906 -330
rect -822 -506 -788 -330
rect -364 -506 -330 -330
rect -246 -506 -212 -330
rect 212 -506 246 -330
rect 330 -506 364 -330
rect 788 -506 822 -330
rect 906 -506 940 -330
rect 1364 -506 1398 -330
rect -1398 -924 -1364 -748
rect -940 -924 -906 -748
rect -822 -924 -788 -748
rect -364 -924 -330 -748
rect -246 -924 -212 -748
rect 212 -924 246 -748
rect 330 -924 364 -748
rect 788 -924 822 -748
rect 906 -924 940 -748
rect 1364 -924 1398 -748
<< mvpsubdiff >>
rect -1544 1146 1544 1158
rect -1544 1112 -1436 1146
rect 1436 1112 1544 1146
rect -1544 1100 1544 1112
rect -1544 1050 -1486 1100
rect -1544 -1050 -1532 1050
rect -1498 -1050 -1486 1050
rect 1486 1050 1544 1100
rect -1544 -1100 -1486 -1050
rect 1486 -1050 1498 1050
rect 1532 -1050 1544 1050
rect 1486 -1100 1544 -1050
rect -1544 -1112 1544 -1100
rect -1544 -1146 -1436 -1112
rect 1436 -1146 1544 -1112
rect -1544 -1158 1544 -1146
<< mvpsubdiffcont >>
rect -1436 1112 1436 1146
rect -1532 -1050 -1498 1050
rect 1498 -1050 1532 1050
rect -1436 -1146 1436 -1112
<< poly >>
rect -1260 1008 -1044 1024
rect -1260 991 -1244 1008
rect -1352 974 -1244 991
rect -1060 991 -1044 1008
rect -684 1008 -468 1024
rect -684 991 -668 1008
rect -1060 974 -952 991
rect -1352 936 -952 974
rect -776 974 -668 991
rect -484 991 -468 1008
rect -108 1008 108 1024
rect -108 991 -92 1008
rect -484 974 -376 991
rect -776 936 -376 974
rect -200 974 -92 991
rect 92 991 108 1008
rect 468 1008 684 1024
rect 468 991 484 1008
rect 92 974 200 991
rect -200 936 200 974
rect 376 974 484 991
rect 668 991 684 1008
rect 1044 1008 1260 1024
rect 1044 991 1060 1008
rect 668 974 776 991
rect 376 936 776 974
rect 952 974 1060 991
rect 1244 991 1260 1008
rect 1244 974 1352 991
rect 952 936 1352 974
rect -1352 698 -952 736
rect -1352 681 -1244 698
rect -1260 664 -1244 681
rect -1060 681 -952 698
rect -776 698 -376 736
rect -776 681 -668 698
rect -1060 664 -1044 681
rect -1260 648 -1044 664
rect -684 664 -668 681
rect -484 681 -376 698
rect -200 698 200 736
rect -200 681 -92 698
rect -484 664 -468 681
rect -684 648 -468 664
rect -108 664 -92 681
rect 92 681 200 698
rect 376 698 776 736
rect 376 681 484 698
rect 92 664 108 681
rect -108 648 108 664
rect 468 664 484 681
rect 668 681 776 698
rect 952 698 1352 736
rect 952 681 1060 698
rect 668 664 684 681
rect 468 648 684 664
rect 1044 664 1060 681
rect 1244 681 1352 698
rect 1244 664 1260 681
rect 1044 648 1260 664
rect -1260 590 -1044 606
rect -1260 573 -1244 590
rect -1352 556 -1244 573
rect -1060 573 -1044 590
rect -684 590 -468 606
rect -684 573 -668 590
rect -1060 556 -952 573
rect -1352 518 -952 556
rect -776 556 -668 573
rect -484 573 -468 590
rect -108 590 108 606
rect -108 573 -92 590
rect -484 556 -376 573
rect -776 518 -376 556
rect -200 556 -92 573
rect 92 573 108 590
rect 468 590 684 606
rect 468 573 484 590
rect 92 556 200 573
rect -200 518 200 556
rect 376 556 484 573
rect 668 573 684 590
rect 1044 590 1260 606
rect 1044 573 1060 590
rect 668 556 776 573
rect 376 518 776 556
rect 952 556 1060 573
rect 1244 573 1260 590
rect 1244 556 1352 573
rect 952 518 1352 556
rect -1352 280 -952 318
rect -1352 263 -1244 280
rect -1260 246 -1244 263
rect -1060 263 -952 280
rect -776 280 -376 318
rect -776 263 -668 280
rect -1060 246 -1044 263
rect -1260 230 -1044 246
rect -684 246 -668 263
rect -484 263 -376 280
rect -200 280 200 318
rect -200 263 -92 280
rect -484 246 -468 263
rect -684 230 -468 246
rect -108 246 -92 263
rect 92 263 200 280
rect 376 280 776 318
rect 376 263 484 280
rect 92 246 108 263
rect -108 230 108 246
rect 468 246 484 263
rect 668 263 776 280
rect 952 280 1352 318
rect 952 263 1060 280
rect 668 246 684 263
rect 468 230 684 246
rect 1044 246 1060 263
rect 1244 263 1352 280
rect 1244 246 1260 263
rect 1044 230 1260 246
rect -1260 172 -1044 188
rect -1260 155 -1244 172
rect -1352 138 -1244 155
rect -1060 155 -1044 172
rect -684 172 -468 188
rect -684 155 -668 172
rect -1060 138 -952 155
rect -1352 100 -952 138
rect -776 138 -668 155
rect -484 155 -468 172
rect -108 172 108 188
rect -108 155 -92 172
rect -484 138 -376 155
rect -776 100 -376 138
rect -200 138 -92 155
rect 92 155 108 172
rect 468 172 684 188
rect 468 155 484 172
rect 92 138 200 155
rect -200 100 200 138
rect 376 138 484 155
rect 668 155 684 172
rect 1044 172 1260 188
rect 1044 155 1060 172
rect 668 138 776 155
rect 376 100 776 138
rect 952 138 1060 155
rect 1244 155 1260 172
rect 1244 138 1352 155
rect 952 100 1352 138
rect -1352 -138 -952 -100
rect -1352 -155 -1244 -138
rect -1260 -172 -1244 -155
rect -1060 -155 -952 -138
rect -776 -138 -376 -100
rect -776 -155 -668 -138
rect -1060 -172 -1044 -155
rect -1260 -188 -1044 -172
rect -684 -172 -668 -155
rect -484 -155 -376 -138
rect -200 -138 200 -100
rect -200 -155 -92 -138
rect -484 -172 -468 -155
rect -684 -188 -468 -172
rect -108 -172 -92 -155
rect 92 -155 200 -138
rect 376 -138 776 -100
rect 376 -155 484 -138
rect 92 -172 108 -155
rect -108 -188 108 -172
rect 468 -172 484 -155
rect 668 -155 776 -138
rect 952 -138 1352 -100
rect 952 -155 1060 -138
rect 668 -172 684 -155
rect 468 -188 684 -172
rect 1044 -172 1060 -155
rect 1244 -155 1352 -138
rect 1244 -172 1260 -155
rect 1044 -188 1260 -172
rect -1260 -246 -1044 -230
rect -1260 -263 -1244 -246
rect -1352 -280 -1244 -263
rect -1060 -263 -1044 -246
rect -684 -246 -468 -230
rect -684 -263 -668 -246
rect -1060 -280 -952 -263
rect -1352 -318 -952 -280
rect -776 -280 -668 -263
rect -484 -263 -468 -246
rect -108 -246 108 -230
rect -108 -263 -92 -246
rect -484 -280 -376 -263
rect -776 -318 -376 -280
rect -200 -280 -92 -263
rect 92 -263 108 -246
rect 468 -246 684 -230
rect 468 -263 484 -246
rect 92 -280 200 -263
rect -200 -318 200 -280
rect 376 -280 484 -263
rect 668 -263 684 -246
rect 1044 -246 1260 -230
rect 1044 -263 1060 -246
rect 668 -280 776 -263
rect 376 -318 776 -280
rect 952 -280 1060 -263
rect 1244 -263 1260 -246
rect 1244 -280 1352 -263
rect 952 -318 1352 -280
rect -1352 -556 -952 -518
rect -1352 -573 -1244 -556
rect -1260 -590 -1244 -573
rect -1060 -573 -952 -556
rect -776 -556 -376 -518
rect -776 -573 -668 -556
rect -1060 -590 -1044 -573
rect -1260 -606 -1044 -590
rect -684 -590 -668 -573
rect -484 -573 -376 -556
rect -200 -556 200 -518
rect -200 -573 -92 -556
rect -484 -590 -468 -573
rect -684 -606 -468 -590
rect -108 -590 -92 -573
rect 92 -573 200 -556
rect 376 -556 776 -518
rect 376 -573 484 -556
rect 92 -590 108 -573
rect -108 -606 108 -590
rect 468 -590 484 -573
rect 668 -573 776 -556
rect 952 -556 1352 -518
rect 952 -573 1060 -556
rect 668 -590 684 -573
rect 468 -606 684 -590
rect 1044 -590 1060 -573
rect 1244 -573 1352 -556
rect 1244 -590 1260 -573
rect 1044 -606 1260 -590
rect -1260 -664 -1044 -648
rect -1260 -681 -1244 -664
rect -1352 -698 -1244 -681
rect -1060 -681 -1044 -664
rect -684 -664 -468 -648
rect -684 -681 -668 -664
rect -1060 -698 -952 -681
rect -1352 -736 -952 -698
rect -776 -698 -668 -681
rect -484 -681 -468 -664
rect -108 -664 108 -648
rect -108 -681 -92 -664
rect -484 -698 -376 -681
rect -776 -736 -376 -698
rect -200 -698 -92 -681
rect 92 -681 108 -664
rect 468 -664 684 -648
rect 468 -681 484 -664
rect 92 -698 200 -681
rect -200 -736 200 -698
rect 376 -698 484 -681
rect 668 -681 684 -664
rect 1044 -664 1260 -648
rect 1044 -681 1060 -664
rect 668 -698 776 -681
rect 376 -736 776 -698
rect 952 -698 1060 -681
rect 1244 -681 1260 -664
rect 1244 -698 1352 -681
rect 952 -736 1352 -698
rect -1352 -974 -952 -936
rect -1352 -991 -1244 -974
rect -1260 -1008 -1244 -991
rect -1060 -991 -952 -974
rect -776 -974 -376 -936
rect -776 -991 -668 -974
rect -1060 -1008 -1044 -991
rect -1260 -1024 -1044 -1008
rect -684 -1008 -668 -991
rect -484 -991 -376 -974
rect -200 -974 200 -936
rect -200 -991 -92 -974
rect -484 -1008 -468 -991
rect -684 -1024 -468 -1008
rect -108 -1008 -92 -991
rect 92 -991 200 -974
rect 376 -974 776 -936
rect 376 -991 484 -974
rect 92 -1008 108 -991
rect -108 -1024 108 -1008
rect 468 -1008 484 -991
rect 668 -991 776 -974
rect 952 -974 1352 -936
rect 952 -991 1060 -974
rect 668 -1008 684 -991
rect 468 -1024 684 -1008
rect 1044 -1008 1060 -991
rect 1244 -991 1352 -974
rect 1244 -1008 1260 -991
rect 1044 -1024 1260 -1008
<< polycont >>
rect -1244 974 -1060 1008
rect -668 974 -484 1008
rect -92 974 92 1008
rect 484 974 668 1008
rect 1060 974 1244 1008
rect -1244 664 -1060 698
rect -668 664 -484 698
rect -92 664 92 698
rect 484 664 668 698
rect 1060 664 1244 698
rect -1244 556 -1060 590
rect -668 556 -484 590
rect -92 556 92 590
rect 484 556 668 590
rect 1060 556 1244 590
rect -1244 246 -1060 280
rect -668 246 -484 280
rect -92 246 92 280
rect 484 246 668 280
rect 1060 246 1244 280
rect -1244 138 -1060 172
rect -668 138 -484 172
rect -92 138 92 172
rect 484 138 668 172
rect 1060 138 1244 172
rect -1244 -172 -1060 -138
rect -668 -172 -484 -138
rect -92 -172 92 -138
rect 484 -172 668 -138
rect 1060 -172 1244 -138
rect -1244 -280 -1060 -246
rect -668 -280 -484 -246
rect -92 -280 92 -246
rect 484 -280 668 -246
rect 1060 -280 1244 -246
rect -1244 -590 -1060 -556
rect -668 -590 -484 -556
rect -92 -590 92 -556
rect 484 -590 668 -556
rect 1060 -590 1244 -556
rect -1244 -698 -1060 -664
rect -668 -698 -484 -664
rect -92 -698 92 -664
rect 484 -698 668 -664
rect 1060 -698 1244 -664
rect -1244 -1008 -1060 -974
rect -668 -1008 -484 -974
rect -92 -1008 92 -974
rect 484 -1008 668 -974
rect 1060 -1008 1244 -974
<< locali >>
rect -1532 1112 -1436 1146
rect 1436 1112 1532 1146
rect -1532 1050 -1498 1112
rect 1498 1050 1532 1112
rect -1260 974 -1244 1008
rect -1060 974 -1044 1008
rect -684 974 -668 1008
rect -484 974 -468 1008
rect -108 974 -92 1008
rect 92 974 108 1008
rect 468 974 484 1008
rect 668 974 684 1008
rect 1044 974 1060 1008
rect 1244 974 1260 1008
rect -1398 924 -1364 940
rect -1398 732 -1364 748
rect -940 924 -906 940
rect -940 732 -906 748
rect -822 924 -788 940
rect -822 732 -788 748
rect -364 924 -330 940
rect -364 732 -330 748
rect -246 924 -212 940
rect -246 732 -212 748
rect 212 924 246 940
rect 212 732 246 748
rect 330 924 364 940
rect 330 732 364 748
rect 788 924 822 940
rect 788 732 822 748
rect 906 924 940 940
rect 906 732 940 748
rect 1364 924 1398 940
rect 1364 732 1398 748
rect -1260 664 -1244 698
rect -1060 664 -1044 698
rect -684 664 -668 698
rect -484 664 -468 698
rect -108 664 -92 698
rect 92 664 108 698
rect 468 664 484 698
rect 668 664 684 698
rect 1044 664 1060 698
rect 1244 664 1260 698
rect -1260 556 -1244 590
rect -1060 556 -1044 590
rect -684 556 -668 590
rect -484 556 -468 590
rect -108 556 -92 590
rect 92 556 108 590
rect 468 556 484 590
rect 668 556 684 590
rect 1044 556 1060 590
rect 1244 556 1260 590
rect -1398 506 -1364 522
rect -1398 314 -1364 330
rect -940 506 -906 522
rect -940 314 -906 330
rect -822 506 -788 522
rect -822 314 -788 330
rect -364 506 -330 522
rect -364 314 -330 330
rect -246 506 -212 522
rect -246 314 -212 330
rect 212 506 246 522
rect 212 314 246 330
rect 330 506 364 522
rect 330 314 364 330
rect 788 506 822 522
rect 788 314 822 330
rect 906 506 940 522
rect 906 314 940 330
rect 1364 506 1398 522
rect 1364 314 1398 330
rect -1260 246 -1244 280
rect -1060 246 -1044 280
rect -684 246 -668 280
rect -484 246 -468 280
rect -108 246 -92 280
rect 92 246 108 280
rect 468 246 484 280
rect 668 246 684 280
rect 1044 246 1060 280
rect 1244 246 1260 280
rect -1260 138 -1244 172
rect -1060 138 -1044 172
rect -684 138 -668 172
rect -484 138 -468 172
rect -108 138 -92 172
rect 92 138 108 172
rect 468 138 484 172
rect 668 138 684 172
rect 1044 138 1060 172
rect 1244 138 1260 172
rect -1398 88 -1364 104
rect -1398 -104 -1364 -88
rect -940 88 -906 104
rect -940 -104 -906 -88
rect -822 88 -788 104
rect -822 -104 -788 -88
rect -364 88 -330 104
rect -364 -104 -330 -88
rect -246 88 -212 104
rect -246 -104 -212 -88
rect 212 88 246 104
rect 212 -104 246 -88
rect 330 88 364 104
rect 330 -104 364 -88
rect 788 88 822 104
rect 788 -104 822 -88
rect 906 88 940 104
rect 906 -104 940 -88
rect 1364 88 1398 104
rect 1364 -104 1398 -88
rect -1260 -172 -1244 -138
rect -1060 -172 -1044 -138
rect -684 -172 -668 -138
rect -484 -172 -468 -138
rect -108 -172 -92 -138
rect 92 -172 108 -138
rect 468 -172 484 -138
rect 668 -172 684 -138
rect 1044 -172 1060 -138
rect 1244 -172 1260 -138
rect -1260 -280 -1244 -246
rect -1060 -280 -1044 -246
rect -684 -280 -668 -246
rect -484 -280 -468 -246
rect -108 -280 -92 -246
rect 92 -280 108 -246
rect 468 -280 484 -246
rect 668 -280 684 -246
rect 1044 -280 1060 -246
rect 1244 -280 1260 -246
rect -1398 -330 -1364 -314
rect -1398 -522 -1364 -506
rect -940 -330 -906 -314
rect -940 -522 -906 -506
rect -822 -330 -788 -314
rect -822 -522 -788 -506
rect -364 -330 -330 -314
rect -364 -522 -330 -506
rect -246 -330 -212 -314
rect -246 -522 -212 -506
rect 212 -330 246 -314
rect 212 -522 246 -506
rect 330 -330 364 -314
rect 330 -522 364 -506
rect 788 -330 822 -314
rect 788 -522 822 -506
rect 906 -330 940 -314
rect 906 -522 940 -506
rect 1364 -330 1398 -314
rect 1364 -522 1398 -506
rect -1260 -590 -1244 -556
rect -1060 -590 -1044 -556
rect -684 -590 -668 -556
rect -484 -590 -468 -556
rect -108 -590 -92 -556
rect 92 -590 108 -556
rect 468 -590 484 -556
rect 668 -590 684 -556
rect 1044 -590 1060 -556
rect 1244 -590 1260 -556
rect -1260 -698 -1244 -664
rect -1060 -698 -1044 -664
rect -684 -698 -668 -664
rect -484 -698 -468 -664
rect -108 -698 -92 -664
rect 92 -698 108 -664
rect 468 -698 484 -664
rect 668 -698 684 -664
rect 1044 -698 1060 -664
rect 1244 -698 1260 -664
rect -1398 -748 -1364 -732
rect -1398 -940 -1364 -924
rect -940 -748 -906 -732
rect -940 -940 -906 -924
rect -822 -748 -788 -732
rect -822 -940 -788 -924
rect -364 -748 -330 -732
rect -364 -940 -330 -924
rect -246 -748 -212 -732
rect -246 -940 -212 -924
rect 212 -748 246 -732
rect 212 -940 246 -924
rect 330 -748 364 -732
rect 330 -940 364 -924
rect 788 -748 822 -732
rect 788 -940 822 -924
rect 906 -748 940 -732
rect 906 -940 940 -924
rect 1364 -748 1398 -732
rect 1364 -940 1398 -924
rect -1260 -1008 -1244 -974
rect -1060 -1008 -1044 -974
rect -684 -1008 -668 -974
rect -484 -1008 -468 -974
rect -108 -1008 -92 -974
rect 92 -1008 108 -974
rect 468 -1008 484 -974
rect 668 -1008 684 -974
rect 1044 -1008 1060 -974
rect 1244 -1008 1260 -974
rect -1532 -1112 -1498 -1050
rect 1498 -1112 1532 -1050
rect -1532 -1146 -1436 -1112
rect 1436 -1146 1532 -1112
<< viali >>
rect -1244 974 -1060 1008
rect -668 974 -484 1008
rect -92 974 92 1008
rect 484 974 668 1008
rect 1060 974 1244 1008
rect -1398 748 -1364 924
rect -940 748 -906 924
rect -822 748 -788 924
rect -364 748 -330 924
rect -246 748 -212 924
rect 212 748 246 924
rect 330 748 364 924
rect 788 748 822 924
rect 906 748 940 924
rect 1364 748 1398 924
rect -1244 664 -1060 698
rect -668 664 -484 698
rect -92 664 92 698
rect 484 664 668 698
rect 1060 664 1244 698
rect -1244 556 -1060 590
rect -668 556 -484 590
rect -92 556 92 590
rect 484 556 668 590
rect 1060 556 1244 590
rect -1398 330 -1364 506
rect -940 330 -906 506
rect -822 330 -788 506
rect -364 330 -330 506
rect -246 330 -212 506
rect 212 330 246 506
rect 330 330 364 506
rect 788 330 822 506
rect 906 330 940 506
rect 1364 330 1398 506
rect -1244 246 -1060 280
rect -668 246 -484 280
rect -92 246 92 280
rect 484 246 668 280
rect 1060 246 1244 280
rect -1244 138 -1060 172
rect -668 138 -484 172
rect -92 138 92 172
rect 484 138 668 172
rect 1060 138 1244 172
rect -1398 -88 -1364 88
rect -940 -88 -906 88
rect -822 -88 -788 88
rect -364 -88 -330 88
rect -246 -88 -212 88
rect 212 -88 246 88
rect 330 -88 364 88
rect 788 -88 822 88
rect 906 -88 940 88
rect 1364 -88 1398 88
rect -1244 -172 -1060 -138
rect -668 -172 -484 -138
rect -92 -172 92 -138
rect 484 -172 668 -138
rect 1060 -172 1244 -138
rect -1244 -280 -1060 -246
rect -668 -280 -484 -246
rect -92 -280 92 -246
rect 484 -280 668 -246
rect 1060 -280 1244 -246
rect -1398 -506 -1364 -330
rect -940 -506 -906 -330
rect -822 -506 -788 -330
rect -364 -506 -330 -330
rect -246 -506 -212 -330
rect 212 -506 246 -330
rect 330 -506 364 -330
rect 788 -506 822 -330
rect 906 -506 940 -330
rect 1364 -506 1398 -330
rect -1244 -590 -1060 -556
rect -668 -590 -484 -556
rect -92 -590 92 -556
rect 484 -590 668 -556
rect 1060 -590 1244 -556
rect -1244 -698 -1060 -664
rect -668 -698 -484 -664
rect -92 -698 92 -664
rect 484 -698 668 -664
rect 1060 -698 1244 -664
rect -1398 -924 -1364 -748
rect -940 -924 -906 -748
rect -822 -924 -788 -748
rect -364 -924 -330 -748
rect -246 -924 -212 -748
rect 212 -924 246 -748
rect 330 -924 364 -748
rect 788 -924 822 -748
rect 906 -924 940 -748
rect 1364 -924 1398 -748
rect -1244 -1008 -1060 -974
rect -668 -1008 -484 -974
rect -92 -1008 92 -974
rect 484 -1008 668 -974
rect 1060 -1008 1244 -974
<< metal1 >>
rect -1256 1008 -1048 1014
rect -1256 974 -1244 1008
rect -1060 974 -1048 1008
rect -1256 968 -1048 974
rect -680 1008 -472 1014
rect -680 974 -668 1008
rect -484 974 -472 1008
rect -680 968 -472 974
rect -104 1008 104 1014
rect -104 974 -92 1008
rect 92 974 104 1008
rect -104 968 104 974
rect 472 1008 680 1014
rect 472 974 484 1008
rect 668 974 680 1008
rect 472 968 680 974
rect 1048 1008 1256 1014
rect 1048 974 1060 1008
rect 1244 974 1256 1008
rect 1048 968 1256 974
rect -1404 924 -1358 936
rect -1404 748 -1398 924
rect -1364 748 -1358 924
rect -1404 736 -1358 748
rect -946 924 -900 936
rect -946 748 -940 924
rect -906 748 -900 924
rect -946 736 -900 748
rect -828 924 -782 936
rect -828 748 -822 924
rect -788 748 -782 924
rect -828 736 -782 748
rect -370 924 -324 936
rect -370 748 -364 924
rect -330 748 -324 924
rect -370 736 -324 748
rect -252 924 -206 936
rect -252 748 -246 924
rect -212 748 -206 924
rect -252 736 -206 748
rect 206 924 252 936
rect 206 748 212 924
rect 246 748 252 924
rect 206 736 252 748
rect 324 924 370 936
rect 324 748 330 924
rect 364 748 370 924
rect 324 736 370 748
rect 782 924 828 936
rect 782 748 788 924
rect 822 748 828 924
rect 782 736 828 748
rect 900 924 946 936
rect 900 748 906 924
rect 940 748 946 924
rect 900 736 946 748
rect 1358 924 1404 936
rect 1358 748 1364 924
rect 1398 748 1404 924
rect 1358 736 1404 748
rect -1256 698 -1048 704
rect -1256 664 -1244 698
rect -1060 664 -1048 698
rect -1256 658 -1048 664
rect -680 698 -472 704
rect -680 664 -668 698
rect -484 664 -472 698
rect -680 658 -472 664
rect -104 698 104 704
rect -104 664 -92 698
rect 92 664 104 698
rect -104 658 104 664
rect 472 698 680 704
rect 472 664 484 698
rect 668 664 680 698
rect 472 658 680 664
rect 1048 698 1256 704
rect 1048 664 1060 698
rect 1244 664 1256 698
rect 1048 658 1256 664
rect -1256 590 -1048 596
rect -1256 556 -1244 590
rect -1060 556 -1048 590
rect -1256 550 -1048 556
rect -680 590 -472 596
rect -680 556 -668 590
rect -484 556 -472 590
rect -680 550 -472 556
rect -104 590 104 596
rect -104 556 -92 590
rect 92 556 104 590
rect -104 550 104 556
rect 472 590 680 596
rect 472 556 484 590
rect 668 556 680 590
rect 472 550 680 556
rect 1048 590 1256 596
rect 1048 556 1060 590
rect 1244 556 1256 590
rect 1048 550 1256 556
rect -1404 506 -1358 518
rect -1404 330 -1398 506
rect -1364 330 -1358 506
rect -1404 318 -1358 330
rect -946 506 -900 518
rect -946 330 -940 506
rect -906 330 -900 506
rect -946 318 -900 330
rect -828 506 -782 518
rect -828 330 -822 506
rect -788 330 -782 506
rect -828 318 -782 330
rect -370 506 -324 518
rect -370 330 -364 506
rect -330 330 -324 506
rect -370 318 -324 330
rect -252 506 -206 518
rect -252 330 -246 506
rect -212 330 -206 506
rect -252 318 -206 330
rect 206 506 252 518
rect 206 330 212 506
rect 246 330 252 506
rect 206 318 252 330
rect 324 506 370 518
rect 324 330 330 506
rect 364 330 370 506
rect 324 318 370 330
rect 782 506 828 518
rect 782 330 788 506
rect 822 330 828 506
rect 782 318 828 330
rect 900 506 946 518
rect 900 330 906 506
rect 940 330 946 506
rect 900 318 946 330
rect 1358 506 1404 518
rect 1358 330 1364 506
rect 1398 330 1404 506
rect 1358 318 1404 330
rect -1256 280 -1048 286
rect -1256 246 -1244 280
rect -1060 246 -1048 280
rect -1256 240 -1048 246
rect -680 280 -472 286
rect -680 246 -668 280
rect -484 246 -472 280
rect -680 240 -472 246
rect -104 280 104 286
rect -104 246 -92 280
rect 92 246 104 280
rect -104 240 104 246
rect 472 280 680 286
rect 472 246 484 280
rect 668 246 680 280
rect 472 240 680 246
rect 1048 280 1256 286
rect 1048 246 1060 280
rect 1244 246 1256 280
rect 1048 240 1256 246
rect -1256 172 -1048 178
rect -1256 138 -1244 172
rect -1060 138 -1048 172
rect -1256 132 -1048 138
rect -680 172 -472 178
rect -680 138 -668 172
rect -484 138 -472 172
rect -680 132 -472 138
rect -104 172 104 178
rect -104 138 -92 172
rect 92 138 104 172
rect -104 132 104 138
rect 472 172 680 178
rect 472 138 484 172
rect 668 138 680 172
rect 472 132 680 138
rect 1048 172 1256 178
rect 1048 138 1060 172
rect 1244 138 1256 172
rect 1048 132 1256 138
rect -1404 88 -1358 100
rect -1404 -88 -1398 88
rect -1364 -88 -1358 88
rect -1404 -100 -1358 -88
rect -946 88 -900 100
rect -946 -88 -940 88
rect -906 -88 -900 88
rect -946 -100 -900 -88
rect -828 88 -782 100
rect -828 -88 -822 88
rect -788 -88 -782 88
rect -828 -100 -782 -88
rect -370 88 -324 100
rect -370 -88 -364 88
rect -330 -88 -324 88
rect -370 -100 -324 -88
rect -252 88 -206 100
rect -252 -88 -246 88
rect -212 -88 -206 88
rect -252 -100 -206 -88
rect 206 88 252 100
rect 206 -88 212 88
rect 246 -88 252 88
rect 206 -100 252 -88
rect 324 88 370 100
rect 324 -88 330 88
rect 364 -88 370 88
rect 324 -100 370 -88
rect 782 88 828 100
rect 782 -88 788 88
rect 822 -88 828 88
rect 782 -100 828 -88
rect 900 88 946 100
rect 900 -88 906 88
rect 940 -88 946 88
rect 900 -100 946 -88
rect 1358 88 1404 100
rect 1358 -88 1364 88
rect 1398 -88 1404 88
rect 1358 -100 1404 -88
rect -1256 -138 -1048 -132
rect -1256 -172 -1244 -138
rect -1060 -172 -1048 -138
rect -1256 -178 -1048 -172
rect -680 -138 -472 -132
rect -680 -172 -668 -138
rect -484 -172 -472 -138
rect -680 -178 -472 -172
rect -104 -138 104 -132
rect -104 -172 -92 -138
rect 92 -172 104 -138
rect -104 -178 104 -172
rect 472 -138 680 -132
rect 472 -172 484 -138
rect 668 -172 680 -138
rect 472 -178 680 -172
rect 1048 -138 1256 -132
rect 1048 -172 1060 -138
rect 1244 -172 1256 -138
rect 1048 -178 1256 -172
rect -1256 -246 -1048 -240
rect -1256 -280 -1244 -246
rect -1060 -280 -1048 -246
rect -1256 -286 -1048 -280
rect -680 -246 -472 -240
rect -680 -280 -668 -246
rect -484 -280 -472 -246
rect -680 -286 -472 -280
rect -104 -246 104 -240
rect -104 -280 -92 -246
rect 92 -280 104 -246
rect -104 -286 104 -280
rect 472 -246 680 -240
rect 472 -280 484 -246
rect 668 -280 680 -246
rect 472 -286 680 -280
rect 1048 -246 1256 -240
rect 1048 -280 1060 -246
rect 1244 -280 1256 -246
rect 1048 -286 1256 -280
rect -1404 -330 -1358 -318
rect -1404 -506 -1398 -330
rect -1364 -506 -1358 -330
rect -1404 -518 -1358 -506
rect -946 -330 -900 -318
rect -946 -506 -940 -330
rect -906 -506 -900 -330
rect -946 -518 -900 -506
rect -828 -330 -782 -318
rect -828 -506 -822 -330
rect -788 -506 -782 -330
rect -828 -518 -782 -506
rect -370 -330 -324 -318
rect -370 -506 -364 -330
rect -330 -506 -324 -330
rect -370 -518 -324 -506
rect -252 -330 -206 -318
rect -252 -506 -246 -330
rect -212 -506 -206 -330
rect -252 -518 -206 -506
rect 206 -330 252 -318
rect 206 -506 212 -330
rect 246 -506 252 -330
rect 206 -518 252 -506
rect 324 -330 370 -318
rect 324 -506 330 -330
rect 364 -506 370 -330
rect 324 -518 370 -506
rect 782 -330 828 -318
rect 782 -506 788 -330
rect 822 -506 828 -330
rect 782 -518 828 -506
rect 900 -330 946 -318
rect 900 -506 906 -330
rect 940 -506 946 -330
rect 900 -518 946 -506
rect 1358 -330 1404 -318
rect 1358 -506 1364 -330
rect 1398 -506 1404 -330
rect 1358 -518 1404 -506
rect -1256 -556 -1048 -550
rect -1256 -590 -1244 -556
rect -1060 -590 -1048 -556
rect -1256 -596 -1048 -590
rect -680 -556 -472 -550
rect -680 -590 -668 -556
rect -484 -590 -472 -556
rect -680 -596 -472 -590
rect -104 -556 104 -550
rect -104 -590 -92 -556
rect 92 -590 104 -556
rect -104 -596 104 -590
rect 472 -556 680 -550
rect 472 -590 484 -556
rect 668 -590 680 -556
rect 472 -596 680 -590
rect 1048 -556 1256 -550
rect 1048 -590 1060 -556
rect 1244 -590 1256 -556
rect 1048 -596 1256 -590
rect -1256 -664 -1048 -658
rect -1256 -698 -1244 -664
rect -1060 -698 -1048 -664
rect -1256 -704 -1048 -698
rect -680 -664 -472 -658
rect -680 -698 -668 -664
rect -484 -698 -472 -664
rect -680 -704 -472 -698
rect -104 -664 104 -658
rect -104 -698 -92 -664
rect 92 -698 104 -664
rect -104 -704 104 -698
rect 472 -664 680 -658
rect 472 -698 484 -664
rect 668 -698 680 -664
rect 472 -704 680 -698
rect 1048 -664 1256 -658
rect 1048 -698 1060 -664
rect 1244 -698 1256 -664
rect 1048 -704 1256 -698
rect -1404 -748 -1358 -736
rect -1404 -924 -1398 -748
rect -1364 -924 -1358 -748
rect -1404 -936 -1358 -924
rect -946 -748 -900 -736
rect -946 -924 -940 -748
rect -906 -924 -900 -748
rect -946 -936 -900 -924
rect -828 -748 -782 -736
rect -828 -924 -822 -748
rect -788 -924 -782 -748
rect -828 -936 -782 -924
rect -370 -748 -324 -736
rect -370 -924 -364 -748
rect -330 -924 -324 -748
rect -370 -936 -324 -924
rect -252 -748 -206 -736
rect -252 -924 -246 -748
rect -212 -924 -206 -748
rect -252 -936 -206 -924
rect 206 -748 252 -736
rect 206 -924 212 -748
rect 246 -924 252 -748
rect 206 -936 252 -924
rect 324 -748 370 -736
rect 324 -924 330 -748
rect 364 -924 370 -748
rect 324 -936 370 -924
rect 782 -748 828 -736
rect 782 -924 788 -748
rect 822 -924 828 -748
rect 782 -936 828 -924
rect 900 -748 946 -736
rect 900 -924 906 -748
rect 940 -924 946 -748
rect 900 -936 946 -924
rect 1358 -748 1404 -736
rect 1358 -924 1364 -748
rect 1398 -924 1404 -748
rect 1358 -936 1404 -924
rect -1256 -974 -1048 -968
rect -1256 -1008 -1244 -974
rect -1060 -1008 -1048 -974
rect -1256 -1014 -1048 -1008
rect -680 -974 -472 -968
rect -680 -1008 -668 -974
rect -484 -1008 -472 -974
rect -680 -1014 -472 -1008
rect -104 -974 104 -968
rect -104 -1008 -92 -974
rect 92 -1008 104 -974
rect -104 -1014 104 -1008
rect 472 -974 680 -968
rect 472 -1008 484 -974
rect 668 -1008 680 -974
rect 472 -1014 680 -1008
rect 1048 -974 1256 -968
rect 1048 -1008 1060 -974
rect 1244 -1008 1256 -974
rect 1048 -1014 1256 -1008
<< properties >>
string FIXED_BBOX -1515 -1129 1515 1129
string gencell sky130_fd_pr__nfet_05v0_nvt
string library sky130
string parameters w 1.0 l 2.0 m 5 nf 5 diffcov 100 polycov 50 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.90 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
