magic
tech sky130A
magscale 1 2
timestamp 1730743893
<< error_p >>
rect 4428 21898 4478 26336
rect 7554 21948 10540 21962
rect 2118 20164 2176 20170
rect 2118 20130 2130 20164
rect 2118 20124 2176 20130
rect 2118 18554 2176 18560
rect 2118 18520 2130 18554
rect 2118 18514 2176 18520
rect 2184 17950 2242 17956
rect 2184 17916 2196 17950
rect 2184 17910 2242 17916
<< error_s >>
rect 2184 16340 2242 16346
rect 2184 16306 2196 16340
rect 2184 16300 2242 16306
rect 4468 10634 4518 15072
rect 7594 10684 10580 10698
rect 2158 8900 2216 8906
rect 2158 8866 2170 8900
rect 2158 8860 2216 8866
rect 2158 7290 2216 7296
rect 2158 7256 2170 7290
rect 2158 7250 2216 7256
rect 2224 6686 2282 6692
rect 2224 6652 2236 6686
rect 2224 6646 2282 6652
rect 2224 5076 2282 5082
rect 2224 5042 2236 5076
rect 2224 5036 2282 5042
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
rect 0 -6400 200 -6200
rect 0 -6800 200 -6600
use sky130_fd_pr__res_xhigh_po_0p35_FDV9Y5  sky130_fd_pr__res_xhigh_po_0p35_FDV9Y5_0 paramcells
timestamp 1729623223
transform 1 0 17765 0 1 12596
box -201 -2582 201 2582
use sky130_fd_pr__res_xhigh_po_0p35_FDV9Y5  sky130_fd_pr__res_xhigh_po_0p35_FDV9Y5_1
timestamp 1729623223
transform 1 0 21547 0 1 12792
box -201 -2582 201 2582
use sky130_fd_pr__res_xhigh_po_0p35_FDV9Y5  sky130_fd_pr__res_xhigh_po_0p35_FDV9Y5_2
timestamp 1729623223
transform 1 0 20601 0 1 12714
box -201 -2582 201 2582
use sky130_fd_pr__res_xhigh_po_0p35_FDV9Y5  sky130_fd_pr__res_xhigh_po_0p35_FDV9Y5_3
timestamp 1729623223
transform 1 0 19537 0 1 12714
box -201 -2582 201 2582
use sky130_fd_pr__res_xhigh_po_0p35_FDV9Y5  sky130_fd_pr__res_xhigh_po_0p35_FDV9Y5_4
timestamp 1729623223
transform 1 0 18553 0 1 12674
box -201 -2582 201 2582
use sky130_fd_pr__res_xhigh_po_0p35_FDVHJ6  sky130_fd_pr__res_xhigh_po_0p35_FDVHJ6_0 paramcells
timestamp 1729623223
transform 1 0 22614 0 1 12792
box -284 -2582 284 2582
use sky130_fd_pr__res_xhigh_po_0p35_FDVHJ6  sky130_fd_pr__res_xhigh_po_0p35_FDVHJ6_1
timestamp 1729623223
transform 1 0 23678 0 1 12792
box -284 -2582 284 2582
use sky130_fd_pr__res_xhigh_po_0p35_HGNRCC  sky130_fd_pr__res_xhigh_po_0p35_HGNRCC_0 paramcells
timestamp 1729623223
transform 1 0 22640 0 1 19212
box -5430 -2582 5430 2582
use sky130_fd_pr__res_xhigh_po_0p35_S4N9LQ  sky130_fd_pr__res_xhigh_po_0p35_S4N9LQ_0 paramcells
timestamp 1729623223
transform 1 0 20732 0 1 6964
box -2774 -2582 2774 2582
use Universal_R_2R_Block2  x1
timestamp 1730737834
transform 1 0 31152 0 1 10818
box 0 -2814 6306 376
use Universal_R_2R_Block2  x2
timestamp 1730737834
transform 1 0 24102 0 1 4044
box 0 -2814 6306 376
use Universal_R_2R_Block2  x3
timestamp 1730737834
transform 1 0 24338 0 1 224
box 0 -2814 6306 376
use Universal_R_2R_Block2  x4
timestamp 1730737834
transform 1 0 24456 0 1 -3518
box 0 -2814 6306 376
use Universal_R_2R_Block2  x5
timestamp 1730737834
transform 1 0 31072 0 1 7078
box 0 -2814 6306 376
use x1_x32_OA  x6
timestamp 1730739923
transform 1 0 1416 0 1 18718
box 0 -2600 14514 7642
use Output_OA  x7
timestamp 1730743893
transform 1 0 656 0 1 -3962
box 628 -1122 15044 8320
use x1_x32_OA  x8
timestamp 1730739923
transform 1 0 1456 0 1 7454
box 0 -2600 14514 7642
use Universal_R_2R_Block2  x9
timestamp 1730737834
transform 1 0 30718 0 1 3690
box 0 -2814 6306 376
use Universal_R_2R_Block2  x10
timestamp 1730737834
transform 1 0 31072 0 1 -130
box 0 -2814 6306 376
use Universal_R_2R_Block2  x11
timestamp 1730737834
transform 1 0 31466 0 1 -3674
box 0 -2814 6306 376
use Universal_R_2R_Block2  x12
timestamp 1730737834
transform 1 0 24140 0 1 7708
box 0 -2814 6306 376
use Universal_R_2R_Block2  x13
timestamp 1730737834
transform 1 0 24534 0 1 11804
box 0 -2814 6306 376
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 V6
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 V5
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 V8
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 V9
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 V7
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 VO1
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 DVDD
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 AVDD
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 VOUT
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 V4
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 V3
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 V2
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 V1
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 V0
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 VCM
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 256 0 0 0 DVSS
port 15 nsew
flabel metal1 0 -6400 200 -6200 0 FreeSans 256 0 0 0 AVSS
port 16 nsew
flabel metal1 0 -6800 200 -6600 0 FreeSans 256 0 0 0 VBIAS
port 17 nsew
<< end >>
