magic
tech sky130A
magscale 1 2
timestamp 1730992657
<< dnwell >>
rect 4136 -18138 33538 19422
<< nwell >>
rect 4056 19214 33618 19502
rect 4056 15034 4342 19214
rect 33332 15034 33618 19214
rect 4056 6360 4400 15034
rect 4056 5286 4342 6360
rect 18658 5864 19012 8508
rect 33270 6360 33618 15034
rect 33332 5314 33618 6360
rect 4056 -3388 4408 5286
rect 4056 -4434 4342 -3388
rect 18666 -3834 19014 -1212
rect 33272 -3360 33618 5314
rect 33330 -3784 33618 -3360
rect 18664 -3884 19014 -3834
rect 33332 -4434 33618 -3784
rect 4056 -13108 4408 -4434
rect 4056 -17910 4342 -13108
rect 18666 -13604 19016 -10960
rect 33274 -13108 33618 -4434
rect 33330 -13532 33618 -13108
rect 33332 -17910 33618 -13532
rect 4056 -18218 33618 -17910
<< nsubdiff >>
rect 4188 19362 33498 19374
rect 4188 19308 4320 19362
rect 33374 19308 33498 19362
rect 4188 19296 33498 19308
rect 4188 19254 4266 19296
rect 4188 -17956 4198 19254
rect 4254 -17956 4266 19254
rect 4188 -18037 4266 -17956
rect 33419 19270 33498 19296
rect 33419 -17940 33430 19270
rect 33486 -17940 33498 19270
rect 33419 -18037 33498 -17940
rect 4188 -18048 33498 -18037
rect 4188 -18102 4342 -18048
rect 33396 -18102 33498 -18048
rect 4188 -18116 33498 -18102
<< nsubdiffcont >>
rect 4320 19308 33374 19362
rect 4198 -17956 4254 19254
rect 33430 -17940 33486 19270
rect 4342 -18102 33396 -18048
<< locali >>
rect 4188 19344 4320 19362
rect 4188 -18098 4196 19344
rect 4256 19308 4320 19344
rect 33374 19342 33498 19362
rect 33374 19308 33426 19342
rect 4256 19250 4398 19308
rect 9028 19250 33426 19308
rect 4256 19224 33426 19250
rect 4256 -18037 4266 19224
rect 18516 8602 20154 9214
rect 17524 -1142 20148 -502
rect 17518 -10860 20156 -10256
rect 33419 -18037 33426 19224
rect 4256 -18044 33426 -18037
rect 4256 -18098 4342 -18044
rect 33368 -18048 33426 -18044
rect 4188 -18108 4342 -18098
rect 33396 -18102 33426 -18048
rect 33368 -18104 33426 -18102
rect 33488 -18104 33498 19342
rect 33368 -18108 33498 -18104
rect 4188 -18116 33498 -18108
<< viali >>
rect 4196 19254 4256 19344
rect 4398 19308 9028 19318
rect 4196 -17956 4198 19254
rect 4198 -17956 4254 19254
rect 4254 -17956 4256 19254
rect 4398 19250 9028 19308
rect 33426 19270 33488 19342
rect 4196 -18098 4256 -17956
rect 33426 -17940 33430 19270
rect 33430 -17940 33486 19270
rect 33486 -17940 33488 19270
rect 4342 -18048 33368 -18044
rect 4342 -18102 33368 -18048
rect 4342 -18108 33368 -18102
rect 33426 -18104 33488 -17940
<< metal1 >>
rect 7288 20969 7488 21596
rect 8176 21396 9078 21596
rect 4488 20894 4988 20916
rect 7288 20912 9615 20969
rect 4488 20628 4506 20894
rect 4968 20884 4988 20894
rect 4968 20634 9082 20884
rect 4968 20628 4988 20634
rect 4488 20610 4988 20628
rect 6038 19636 6720 19652
rect 6038 19434 6074 19636
rect 6706 19564 6720 19636
rect 6706 19434 9174 19564
rect 6038 19420 9174 19434
rect 4188 19354 4266 19362
rect 4188 19344 9084 19354
rect 4188 6898 4196 19344
rect 4256 19318 9084 19344
rect 4256 19250 4398 19318
rect 9028 19250 9084 19318
rect 4256 19224 9084 19250
rect 33418 19342 33498 19362
rect 4188 5940 4194 6898
rect 4188 -2854 4196 5940
rect 4256 1398 4266 19224
rect 6862 14517 6928 16823
rect 33418 11150 33426 19342
rect 33488 11150 33498 19342
rect 33418 10310 33424 11150
rect 33490 10310 33498 11150
rect 4258 564 4266 1398
rect 4256 -2854 4266 564
rect 6864 -2624 7218 -2610
rect 6864 -2716 6882 -2624
rect 7200 -2716 7218 -2624
rect 6864 -2728 7218 -2716
rect 4188 -3804 4194 -2854
rect 4258 -3804 4266 -2854
rect 4188 -18098 4196 -3804
rect 4256 -12574 4266 -3804
rect 33418 -2828 33426 10310
rect 33488 1428 33498 10310
rect 33492 594 33498 1428
rect 33488 -2828 33498 594
rect 33418 -3772 33424 -2828
rect 33490 -3772 33498 -2828
rect 30422 -3938 30814 -3928
rect 30422 -4030 30442 -3938
rect 30800 -4030 30814 -3938
rect 30422 -4044 30814 -4030
rect 17512 -10862 18648 -10252
rect 19006 -10862 20158 -10252
rect 4258 -13522 4266 -12574
rect 4256 -18036 4266 -13522
rect 18333 -13624 18806 -13546
rect 17956 -13640 18412 -13624
rect 17956 -13734 17970 -13640
rect 18394 -13734 18412 -13640
rect 17956 -13746 18412 -13734
rect 33418 -18036 33426 -3772
rect 33488 -8322 33498 -3772
rect 33490 -9154 33498 -8322
rect 4256 -18044 33426 -18036
rect 4256 -18098 4342 -18044
rect 4188 -18108 4342 -18098
rect 33368 -18104 33426 -18044
rect 33488 -18104 33498 -9154
rect 33368 -18108 33498 -18104
rect 4188 -18116 33498 -18108
<< via1 >>
rect 4506 20628 4968 20894
rect 6074 19434 6706 19636
rect 4198 10312 4256 11144
rect 4194 5940 4196 6898
rect 4196 5940 4256 6898
rect 6728 17108 6928 17244
rect 33424 10310 33426 11150
rect 33426 10310 33488 11150
rect 33488 10310 33490 11150
rect 19308 5128 23984 5180
rect 4198 564 4256 1398
rect 4256 564 4258 1398
rect 6882 -2716 7200 -2624
rect 4194 -3804 4196 -2854
rect 4196 -3804 4256 -2854
rect 4256 -3804 4258 -2854
rect 4198 -9160 4256 -8320
rect 33432 5950 33488 6890
rect 33426 594 33488 1428
rect 33488 594 33492 1428
rect 33424 -3772 33426 -2828
rect 33426 -3772 33488 -2828
rect 33488 -3772 33490 -2828
rect 30442 -4030 30800 -3938
rect 4196 -13522 4256 -12574
rect 4256 -13522 4258 -12574
rect 4196 -15736 4254 -14594
rect 17970 -13734 18394 -13640
rect 33426 -9154 33488 -8322
rect 33488 -9154 33490 -8322
rect 33432 -13522 33484 -12578
rect 33428 -15736 33486 -14596
<< metal2 >>
rect 10930 21624 11130 21824
rect 13330 21624 13530 21824
rect 15730 21624 15930 21824
rect 18130 21624 18330 21824
rect 20530 21624 20730 21824
rect 22930 21624 23130 21824
rect 25330 21624 25530 21824
rect 27730 21624 27930 21824
rect 30130 21624 30330 21824
rect 32530 21624 32730 21824
rect 4488 20894 4988 20916
rect 4488 20628 4506 20894
rect 4968 20628 4988 20894
rect 4488 20610 4988 20628
rect 6038 19636 6720 19652
rect 6038 19434 6074 19636
rect 6706 19434 6720 19636
rect 6038 19420 6720 19434
rect 4052 17244 4252 17272
rect 4052 17108 6728 17244
rect 6928 17108 6940 17244
rect 4052 17072 4252 17108
rect 6432 16264 6830 16280
rect 6432 15492 6460 16264
rect 6708 15492 6830 16264
rect 6432 15478 6830 15492
rect 4184 11144 4496 11158
rect 4184 10312 4198 11144
rect 4256 10312 4496 11144
rect 4184 10302 4496 10312
rect 33174 11150 33500 11158
rect 33174 10310 33424 11150
rect 33490 10310 33500 11150
rect 33174 10302 33500 10310
rect 4186 6898 4494 6904
rect 4186 5940 4194 6898
rect 4256 5940 4494 6898
rect 4186 5934 4494 5940
rect 33170 6890 33498 6904
rect 33170 5950 33432 6890
rect 33488 5950 33498 6890
rect 33170 5934 33498 5950
rect 4054 5624 4368 5824
rect 33174 1428 33502 1438
rect 4174 1398 4502 1410
rect 4174 564 4198 1398
rect 4258 564 4502 1398
rect 33174 594 33426 1428
rect 33492 594 33502 1428
rect 33174 582 33502 594
rect 4174 554 4502 564
rect 6864 -2624 7218 -2610
rect 6864 -2716 6882 -2624
rect 7200 -2716 7218 -2624
rect 6864 -2728 7218 -2716
rect 33168 -2828 33510 -2816
rect 4178 -2854 4502 -2844
rect 4178 -3804 4194 -2854
rect 4258 -3804 4502 -2854
rect 33168 -3772 33424 -2828
rect 33490 -3772 33510 -2828
rect 33168 -3786 33510 -3772
rect 4178 -3814 4502 -3804
rect 4056 -4100 4364 -3900
rect 30422 -3938 30814 -3928
rect 30422 -4030 30442 -3938
rect 30800 -4030 30814 -3938
rect 30422 -4044 30814 -4030
rect 4180 -8320 4502 -8310
rect 4180 -9160 4198 -8320
rect 4256 -9160 4502 -8320
rect 4180 -9166 4502 -9160
rect 33174 -8322 33502 -8310
rect 33174 -9154 33426 -8322
rect 33490 -9154 33502 -8322
rect 33174 -9166 33502 -9154
rect 4182 -12574 4502 -12564
rect 4182 -13522 4196 -12574
rect 4258 -13522 4502 -12574
rect 4182 -13534 4502 -13522
rect 33180 -12578 33504 -12564
rect 33180 -13522 33432 -12578
rect 33484 -13522 33504 -12578
rect 33180 -13534 33504 -13522
rect 11160 -13640 18408 -13626
rect 11160 -13734 17970 -13640
rect 18394 -13734 18408 -13640
rect 11160 -13754 18408 -13734
rect 4072 -14594 33582 -14582
rect 4072 -15736 4196 -14594
rect 4254 -14596 33582 -14594
rect 4254 -14620 33428 -14596
rect 4254 -15722 4528 -14620
rect 4958 -14622 33428 -14620
rect 4958 -15722 32730 -14622
rect 4254 -15724 32730 -15722
rect 33160 -15724 33428 -14622
rect 4254 -15736 33428 -15724
rect 33486 -15736 33582 -14596
rect 4072 -15746 33582 -15736
rect 4074 -16008 33584 -15980
rect 4074 -16014 30978 -16008
rect 4074 -17122 6480 -16014
rect 6698 -17116 30978 -16014
rect 31196 -17116 33584 -16008
rect 6698 -17122 33584 -17116
rect 4074 -17144 33584 -17122
<< via2 >>
rect 4506 20628 4968 20894
rect 6074 19434 6706 19636
rect 6460 15492 6708 16264
rect 6882 -2716 7200 -2624
rect 30442 -4030 30800 -3938
rect 4528 -15722 4958 -14620
rect 32730 -15724 33160 -14622
rect 6480 -17122 6698 -16014
rect 30978 -17116 31196 -16008
<< metal3 >>
rect 4488 20894 4988 21604
rect 4488 20628 4506 20894
rect 4968 20628 4988 20894
rect 4488 15290 4988 20628
rect 6062 19636 6720 21604
rect 6062 19434 6074 19636
rect 6706 19434 6720 19636
rect 6062 16264 6720 19434
rect 6062 15492 6460 16264
rect 6708 15492 6720 16264
rect 6062 15304 6720 15492
rect 6062 14956 6452 15304
rect 6864 -2624 7218 -2610
rect 6864 -2716 6882 -2624
rect 7200 -2716 7218 -2624
rect 6864 -2728 7218 -2716
rect 6874 -3938 6974 -2728
rect 30422 -3938 30814 -3928
rect 6868 -4030 30442 -3938
rect 30800 -4030 30814 -3938
rect 6868 -4038 30814 -4030
rect 30422 -4044 30814 -4038
rect 4496 -14620 4996 -13524
rect 4496 -15722 4528 -14620
rect 4958 -15722 4996 -14620
rect 4496 -17914 4996 -15722
rect 6458 -16014 6728 -12304
rect 6458 -17122 6480 -16014
rect 6698 -17122 6728 -16014
rect 6458 -17898 6728 -17122
rect 18892 -18218 19104 -18018
use Parallel_10B_Block2  x1
timestamp 1730992657
transform -1 0 33758 0 1 -6634
box 364 -11384 29434 28258
use Input_Stage_v1  x2
timestamp 1730992408
transform -1 0 33454 0 1 23250
box 14128 -37044 29148 -7862
use vbias_gen_pga  x3
timestamp 1730992408
transform 1 0 7039 0 1 16343
box -311 -865 845 909
<< labels >>
flabel metal2 4052 17072 4252 17272 0 FreeSans 256 0 0 0 IBIAS
port 11 nsew
flabel metal2 32530 21624 32730 21824 0 FreeSans 256 90 0 0 V[0]
port 9 nsew
flabel metal2 30130 21624 30330 21824 0 FreeSans 256 90 0 0 V[1]
port 8 nsew
flabel metal2 27730 21624 27930 21824 0 FreeSans 256 90 0 0 V[2]
port 7 nsew
flabel metal2 25330 21624 25530 21824 0 FreeSans 256 90 0 0 V[3]
port 6 nsew
flabel metal2 22930 21624 23130 21824 0 FreeSans 256 90 0 0 V[4]
port 5 nsew
flabel metal2 20530 21624 20730 21824 0 FreeSans 256 90 0 0 V[5]
port 4 nsew
flabel metal2 18130 21624 18330 21824 0 FreeSans 256 90 0 0 V[6]
port 3 nsew
flabel metal2 15730 21624 15930 21824 0 FreeSans 256 90 0 0 V[7]
port 2 nsew
flabel metal2 13330 21624 13530 21824 0 FreeSans 256 90 0 0 V[8]
port 1 nsew
flabel metal2 10930 21624 11130 21824 0 FreeSans 256 90 0 0 V[9]
port 0 nsew
flabel metal2 4056 -4100 4256 -3900 0 FreeSans 256 0 0 0 VIN
port 13 nsew
flabel metal2 4054 5624 4254 5824 0 FreeSans 256 0 0 0 VCM
port 10 nsew
flabel metal3 18900 -18218 19100 -18018 0 FreeSans 256 0 0 0 VOUT
port 15 nsew
flabel metal3 4616 21394 4816 21594 0 FreeSans 256 0 0 0 AVDD
port 12 nsew
flabel metal3 6308 21396 6508 21596 0 FreeSans 256 0 0 0 AVSS
port 16 nsew
flabel metal1 8176 21396 8376 21596 0 FreeSans 256 0 0 0 DVSS
port 17 nsew
flabel metal1 7288 21396 7488 21596 0 FreeSans 256 0 0 0 DVDD
port 14 nsew
<< end >>
