magic
tech sky130A
magscale 1 2
timestamp 1730948043
<< nwell >>
rect -1559 -1297 1559 1297
<< mvpmos >>
rect -1301 -1000 -1201 1000
rect -1023 -1000 -923 1000
rect -745 -1000 -645 1000
rect -467 -1000 -367 1000
rect -189 -1000 -89 1000
rect 89 -1000 189 1000
rect 367 -1000 467 1000
rect 645 -1000 745 1000
rect 923 -1000 1023 1000
rect 1201 -1000 1301 1000
<< mvpdiff >>
rect -1359 988 -1301 1000
rect -1359 -988 -1347 988
rect -1313 -988 -1301 988
rect -1359 -1000 -1301 -988
rect -1201 988 -1143 1000
rect -1201 -988 -1189 988
rect -1155 -988 -1143 988
rect -1201 -1000 -1143 -988
rect -1081 988 -1023 1000
rect -1081 -988 -1069 988
rect -1035 -988 -1023 988
rect -1081 -1000 -1023 -988
rect -923 988 -865 1000
rect -923 -988 -911 988
rect -877 -988 -865 988
rect -923 -1000 -865 -988
rect -803 988 -745 1000
rect -803 -988 -791 988
rect -757 -988 -745 988
rect -803 -1000 -745 -988
rect -645 988 -587 1000
rect -645 -988 -633 988
rect -599 -988 -587 988
rect -645 -1000 -587 -988
rect -525 988 -467 1000
rect -525 -988 -513 988
rect -479 -988 -467 988
rect -525 -1000 -467 -988
rect -367 988 -309 1000
rect -367 -988 -355 988
rect -321 -988 -309 988
rect -367 -1000 -309 -988
rect -247 988 -189 1000
rect -247 -988 -235 988
rect -201 -988 -189 988
rect -247 -1000 -189 -988
rect -89 988 -31 1000
rect -89 -988 -77 988
rect -43 -988 -31 988
rect -89 -1000 -31 -988
rect 31 988 89 1000
rect 31 -988 43 988
rect 77 -988 89 988
rect 31 -1000 89 -988
rect 189 988 247 1000
rect 189 -988 201 988
rect 235 -988 247 988
rect 189 -1000 247 -988
rect 309 988 367 1000
rect 309 -988 321 988
rect 355 -988 367 988
rect 309 -1000 367 -988
rect 467 988 525 1000
rect 467 -988 479 988
rect 513 -988 525 988
rect 467 -1000 525 -988
rect 587 988 645 1000
rect 587 -988 599 988
rect 633 -988 645 988
rect 587 -1000 645 -988
rect 745 988 803 1000
rect 745 -988 757 988
rect 791 -988 803 988
rect 745 -1000 803 -988
rect 865 988 923 1000
rect 865 -988 877 988
rect 911 -988 923 988
rect 865 -1000 923 -988
rect 1023 988 1081 1000
rect 1023 -988 1035 988
rect 1069 -988 1081 988
rect 1023 -1000 1081 -988
rect 1143 988 1201 1000
rect 1143 -988 1155 988
rect 1189 -988 1201 988
rect 1143 -1000 1201 -988
rect 1301 988 1359 1000
rect 1301 -988 1313 988
rect 1347 -988 1359 988
rect 1301 -1000 1359 -988
<< mvpdiffc >>
rect -1347 -988 -1313 988
rect -1189 -988 -1155 988
rect -1069 -988 -1035 988
rect -911 -988 -877 988
rect -791 -988 -757 988
rect -633 -988 -599 988
rect -513 -988 -479 988
rect -355 -988 -321 988
rect -235 -988 -201 988
rect -77 -988 -43 988
rect 43 -988 77 988
rect 201 -988 235 988
rect 321 -988 355 988
rect 479 -988 513 988
rect 599 -988 633 988
rect 757 -988 791 988
rect 877 -988 911 988
rect 1035 -988 1069 988
rect 1155 -988 1189 988
rect 1313 -988 1347 988
<< mvnsubdiff >>
rect -1493 1219 1493 1231
rect -1493 1185 -1385 1219
rect 1385 1185 1493 1219
rect -1493 1173 1493 1185
rect -1493 1123 -1435 1173
rect -1493 -1123 -1481 1123
rect -1447 -1123 -1435 1123
rect 1435 1123 1493 1173
rect -1493 -1173 -1435 -1123
rect 1435 -1123 1447 1123
rect 1481 -1123 1493 1123
rect 1435 -1173 1493 -1123
rect -1493 -1185 1493 -1173
rect -1493 -1219 -1385 -1185
rect 1385 -1219 1493 -1185
rect -1493 -1231 1493 -1219
<< mvnsubdiffcont >>
rect -1385 1185 1385 1219
rect -1481 -1123 -1447 1123
rect 1447 -1123 1481 1123
rect -1385 -1219 1385 -1185
<< poly >>
rect -1301 1081 -1201 1097
rect -1301 1047 -1285 1081
rect -1217 1047 -1201 1081
rect -1301 1000 -1201 1047
rect -1023 1081 -923 1097
rect -1023 1047 -1007 1081
rect -939 1047 -923 1081
rect -1023 1000 -923 1047
rect -745 1081 -645 1097
rect -745 1047 -729 1081
rect -661 1047 -645 1081
rect -745 1000 -645 1047
rect -467 1081 -367 1097
rect -467 1047 -451 1081
rect -383 1047 -367 1081
rect -467 1000 -367 1047
rect -189 1081 -89 1097
rect -189 1047 -173 1081
rect -105 1047 -89 1081
rect -189 1000 -89 1047
rect 89 1081 189 1097
rect 89 1047 105 1081
rect 173 1047 189 1081
rect 89 1000 189 1047
rect 367 1081 467 1097
rect 367 1047 383 1081
rect 451 1047 467 1081
rect 367 1000 467 1047
rect 645 1081 745 1097
rect 645 1047 661 1081
rect 729 1047 745 1081
rect 645 1000 745 1047
rect 923 1081 1023 1097
rect 923 1047 939 1081
rect 1007 1047 1023 1081
rect 923 1000 1023 1047
rect 1201 1081 1301 1097
rect 1201 1047 1217 1081
rect 1285 1047 1301 1081
rect 1201 1000 1301 1047
rect -1301 -1047 -1201 -1000
rect -1301 -1081 -1285 -1047
rect -1217 -1081 -1201 -1047
rect -1301 -1097 -1201 -1081
rect -1023 -1047 -923 -1000
rect -1023 -1081 -1007 -1047
rect -939 -1081 -923 -1047
rect -1023 -1097 -923 -1081
rect -745 -1047 -645 -1000
rect -745 -1081 -729 -1047
rect -661 -1081 -645 -1047
rect -745 -1097 -645 -1081
rect -467 -1047 -367 -1000
rect -467 -1081 -451 -1047
rect -383 -1081 -367 -1047
rect -467 -1097 -367 -1081
rect -189 -1047 -89 -1000
rect -189 -1081 -173 -1047
rect -105 -1081 -89 -1047
rect -189 -1097 -89 -1081
rect 89 -1047 189 -1000
rect 89 -1081 105 -1047
rect 173 -1081 189 -1047
rect 89 -1097 189 -1081
rect 367 -1047 467 -1000
rect 367 -1081 383 -1047
rect 451 -1081 467 -1047
rect 367 -1097 467 -1081
rect 645 -1047 745 -1000
rect 645 -1081 661 -1047
rect 729 -1081 745 -1047
rect 645 -1097 745 -1081
rect 923 -1047 1023 -1000
rect 923 -1081 939 -1047
rect 1007 -1081 1023 -1047
rect 923 -1097 1023 -1081
rect 1201 -1047 1301 -1000
rect 1201 -1081 1217 -1047
rect 1285 -1081 1301 -1047
rect 1201 -1097 1301 -1081
<< polycont >>
rect -1285 1047 -1217 1081
rect -1007 1047 -939 1081
rect -729 1047 -661 1081
rect -451 1047 -383 1081
rect -173 1047 -105 1081
rect 105 1047 173 1081
rect 383 1047 451 1081
rect 661 1047 729 1081
rect 939 1047 1007 1081
rect 1217 1047 1285 1081
rect -1285 -1081 -1217 -1047
rect -1007 -1081 -939 -1047
rect -729 -1081 -661 -1047
rect -451 -1081 -383 -1047
rect -173 -1081 -105 -1047
rect 105 -1081 173 -1047
rect 383 -1081 451 -1047
rect 661 -1081 729 -1047
rect 939 -1081 1007 -1047
rect 1217 -1081 1285 -1047
<< locali >>
rect -1481 1185 -1385 1219
rect 1385 1185 1481 1219
rect -1481 1123 -1447 1185
rect 1447 1123 1481 1185
rect -1301 1047 -1285 1081
rect -1217 1047 -1201 1081
rect -1023 1047 -1007 1081
rect -939 1047 -923 1081
rect -745 1047 -729 1081
rect -661 1047 -645 1081
rect -467 1047 -451 1081
rect -383 1047 -367 1081
rect -189 1047 -173 1081
rect -105 1047 -89 1081
rect 89 1047 105 1081
rect 173 1047 189 1081
rect 367 1047 383 1081
rect 451 1047 467 1081
rect 645 1047 661 1081
rect 729 1047 745 1081
rect 923 1047 939 1081
rect 1007 1047 1023 1081
rect 1201 1047 1217 1081
rect 1285 1047 1301 1081
rect -1347 988 -1313 1004
rect -1347 -1004 -1313 -988
rect -1189 988 -1155 1004
rect -1189 -1004 -1155 -988
rect -1069 988 -1035 1004
rect -1069 -1004 -1035 -988
rect -911 988 -877 1004
rect -911 -1004 -877 -988
rect -791 988 -757 1004
rect -791 -1004 -757 -988
rect -633 988 -599 1004
rect -633 -1004 -599 -988
rect -513 988 -479 1004
rect -513 -1004 -479 -988
rect -355 988 -321 1004
rect -355 -1004 -321 -988
rect -235 988 -201 1004
rect -235 -1004 -201 -988
rect -77 988 -43 1004
rect -77 -1004 -43 -988
rect 43 988 77 1004
rect 43 -1004 77 -988
rect 201 988 235 1004
rect 201 -1004 235 -988
rect 321 988 355 1004
rect 321 -1004 355 -988
rect 479 988 513 1004
rect 479 -1004 513 -988
rect 599 988 633 1004
rect 599 -1004 633 -988
rect 757 988 791 1004
rect 757 -1004 791 -988
rect 877 988 911 1004
rect 877 -1004 911 -988
rect 1035 988 1069 1004
rect 1035 -1004 1069 -988
rect 1155 988 1189 1004
rect 1155 -1004 1189 -988
rect 1313 988 1347 1004
rect 1313 -1004 1347 -988
rect -1301 -1081 -1285 -1047
rect -1217 -1081 -1201 -1047
rect -1023 -1081 -1007 -1047
rect -939 -1081 -923 -1047
rect -745 -1081 -729 -1047
rect -661 -1081 -645 -1047
rect -467 -1081 -451 -1047
rect -383 -1081 -367 -1047
rect -189 -1081 -173 -1047
rect -105 -1081 -89 -1047
rect 89 -1081 105 -1047
rect 173 -1081 189 -1047
rect 367 -1081 383 -1047
rect 451 -1081 467 -1047
rect 645 -1081 661 -1047
rect 729 -1081 745 -1047
rect 923 -1081 939 -1047
rect 1007 -1081 1023 -1047
rect 1201 -1081 1217 -1047
rect 1285 -1081 1301 -1047
rect -1481 -1185 -1447 -1123
rect 1447 -1185 1481 -1123
rect -1481 -1219 -1385 -1185
rect 1385 -1219 1481 -1185
<< viali >>
rect -1285 1047 -1217 1081
rect -1007 1047 -939 1081
rect -729 1047 -661 1081
rect -451 1047 -383 1081
rect -173 1047 -105 1081
rect 105 1047 173 1081
rect 383 1047 451 1081
rect 661 1047 729 1081
rect 939 1047 1007 1081
rect 1217 1047 1285 1081
rect -1347 -988 -1313 988
rect -1189 -988 -1155 988
rect -1069 -988 -1035 988
rect -911 -988 -877 988
rect -791 -988 -757 988
rect -633 -988 -599 988
rect -513 -988 -479 988
rect -355 -988 -321 988
rect -235 -988 -201 988
rect -77 -988 -43 988
rect 43 -988 77 988
rect 201 -988 235 988
rect 321 -988 355 988
rect 479 -988 513 988
rect 599 -988 633 988
rect 757 -988 791 988
rect 877 -988 911 988
rect 1035 -988 1069 988
rect 1155 -988 1189 988
rect 1313 -988 1347 988
rect -1285 -1081 -1217 -1047
rect -1007 -1081 -939 -1047
rect -729 -1081 -661 -1047
rect -451 -1081 -383 -1047
rect -173 -1081 -105 -1047
rect 105 -1081 173 -1047
rect 383 -1081 451 -1047
rect 661 -1081 729 -1047
rect 939 -1081 1007 -1047
rect 1217 -1081 1285 -1047
<< metal1 >>
rect -1297 1081 -1205 1087
rect -1297 1047 -1285 1081
rect -1217 1047 -1205 1081
rect -1297 1041 -1205 1047
rect -1019 1081 -927 1087
rect -1019 1047 -1007 1081
rect -939 1047 -927 1081
rect -1019 1041 -927 1047
rect -741 1081 -649 1087
rect -741 1047 -729 1081
rect -661 1047 -649 1081
rect -741 1041 -649 1047
rect -463 1081 -371 1087
rect -463 1047 -451 1081
rect -383 1047 -371 1081
rect -463 1041 -371 1047
rect -185 1081 -93 1087
rect -185 1047 -173 1081
rect -105 1047 -93 1081
rect -185 1041 -93 1047
rect 93 1081 185 1087
rect 93 1047 105 1081
rect 173 1047 185 1081
rect 93 1041 185 1047
rect 371 1081 463 1087
rect 371 1047 383 1081
rect 451 1047 463 1081
rect 371 1041 463 1047
rect 649 1081 741 1087
rect 649 1047 661 1081
rect 729 1047 741 1081
rect 649 1041 741 1047
rect 927 1081 1019 1087
rect 927 1047 939 1081
rect 1007 1047 1019 1081
rect 927 1041 1019 1047
rect 1205 1081 1297 1087
rect 1205 1047 1217 1081
rect 1285 1047 1297 1081
rect 1205 1041 1297 1047
rect -1353 988 -1307 1000
rect -1353 -988 -1347 988
rect -1313 -988 -1307 988
rect -1353 -1000 -1307 -988
rect -1195 988 -1149 1000
rect -1195 -988 -1189 988
rect -1155 -988 -1149 988
rect -1195 -1000 -1149 -988
rect -1075 988 -1029 1000
rect -1075 -988 -1069 988
rect -1035 -988 -1029 988
rect -1075 -1000 -1029 -988
rect -917 988 -871 1000
rect -917 -988 -911 988
rect -877 -988 -871 988
rect -917 -1000 -871 -988
rect -797 988 -751 1000
rect -797 -988 -791 988
rect -757 -988 -751 988
rect -797 -1000 -751 -988
rect -639 988 -593 1000
rect -639 -988 -633 988
rect -599 -988 -593 988
rect -639 -1000 -593 -988
rect -519 988 -473 1000
rect -519 -988 -513 988
rect -479 -988 -473 988
rect -519 -1000 -473 -988
rect -361 988 -315 1000
rect -361 -988 -355 988
rect -321 -988 -315 988
rect -361 -1000 -315 -988
rect -241 988 -195 1000
rect -241 -988 -235 988
rect -201 -988 -195 988
rect -241 -1000 -195 -988
rect -83 988 -37 1000
rect -83 -988 -77 988
rect -43 -988 -37 988
rect -83 -1000 -37 -988
rect 37 988 83 1000
rect 37 -988 43 988
rect 77 -988 83 988
rect 37 -1000 83 -988
rect 195 988 241 1000
rect 195 -988 201 988
rect 235 -988 241 988
rect 195 -1000 241 -988
rect 315 988 361 1000
rect 315 -988 321 988
rect 355 -988 361 988
rect 315 -1000 361 -988
rect 473 988 519 1000
rect 473 -988 479 988
rect 513 -988 519 988
rect 473 -1000 519 -988
rect 593 988 639 1000
rect 593 -988 599 988
rect 633 -988 639 988
rect 593 -1000 639 -988
rect 751 988 797 1000
rect 751 -988 757 988
rect 791 -988 797 988
rect 751 -1000 797 -988
rect 871 988 917 1000
rect 871 -988 877 988
rect 911 -988 917 988
rect 871 -1000 917 -988
rect 1029 988 1075 1000
rect 1029 -988 1035 988
rect 1069 -988 1075 988
rect 1029 -1000 1075 -988
rect 1149 988 1195 1000
rect 1149 -988 1155 988
rect 1189 -988 1195 988
rect 1149 -1000 1195 -988
rect 1307 988 1353 1000
rect 1307 -988 1313 988
rect 1347 -988 1353 988
rect 1307 -1000 1353 -988
rect -1297 -1047 -1205 -1041
rect -1297 -1081 -1285 -1047
rect -1217 -1081 -1205 -1047
rect -1297 -1087 -1205 -1081
rect -1019 -1047 -927 -1041
rect -1019 -1081 -1007 -1047
rect -939 -1081 -927 -1047
rect -1019 -1087 -927 -1081
rect -741 -1047 -649 -1041
rect -741 -1081 -729 -1047
rect -661 -1081 -649 -1047
rect -741 -1087 -649 -1081
rect -463 -1047 -371 -1041
rect -463 -1081 -451 -1047
rect -383 -1081 -371 -1047
rect -463 -1087 -371 -1081
rect -185 -1047 -93 -1041
rect -185 -1081 -173 -1047
rect -105 -1081 -93 -1047
rect -185 -1087 -93 -1081
rect 93 -1047 185 -1041
rect 93 -1081 105 -1047
rect 173 -1081 185 -1047
rect 93 -1087 185 -1081
rect 371 -1047 463 -1041
rect 371 -1081 383 -1047
rect 451 -1081 463 -1047
rect 371 -1087 463 -1081
rect 649 -1047 741 -1041
rect 649 -1081 661 -1047
rect 729 -1081 741 -1047
rect 649 -1087 741 -1081
rect 927 -1047 1019 -1041
rect 927 -1081 939 -1047
rect 1007 -1081 1019 -1047
rect 927 -1087 1019 -1081
rect 1205 -1047 1297 -1041
rect 1205 -1081 1217 -1047
rect 1285 -1081 1297 -1047
rect 1205 -1087 1297 -1081
<< properties >>
string FIXED_BBOX -1464 -1202 1464 1202
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 10.0 l 0.5 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
