magic
tech sky130A
magscale 1 2
timestamp 1729623223
<< pwell >>
rect -5430 -2582 5430 2582
<< psubdiff >>
rect -5394 2512 -5298 2546
rect 5298 2512 5394 2546
rect -5394 2450 -5360 2512
rect 5360 2450 5394 2512
rect -5394 -2512 -5360 -2450
rect 5360 -2512 5394 -2450
rect -5394 -2546 -5298 -2512
rect 5298 -2546 5394 -2512
<< psubdiffcont >>
rect -5298 2512 5298 2546
rect -5394 -2450 -5360 2450
rect 5360 -2450 5394 2450
rect -5298 -2546 5298 -2512
<< xpolycontact >>
rect -5264 1984 -5194 2416
rect -5264 -2416 -5194 -1984
rect -5098 1984 -5028 2416
rect -5098 -2416 -5028 -1984
rect -4932 1984 -4862 2416
rect -4932 -2416 -4862 -1984
rect -4766 1984 -4696 2416
rect -4766 -2416 -4696 -1984
rect -4600 1984 -4530 2416
rect -4600 -2416 -4530 -1984
rect -4434 1984 -4364 2416
rect -4434 -2416 -4364 -1984
rect -4268 1984 -4198 2416
rect -4268 -2416 -4198 -1984
rect -4102 1984 -4032 2416
rect -4102 -2416 -4032 -1984
rect -3936 1984 -3866 2416
rect -3936 -2416 -3866 -1984
rect -3770 1984 -3700 2416
rect -3770 -2416 -3700 -1984
rect -3604 1984 -3534 2416
rect -3604 -2416 -3534 -1984
rect -3438 1984 -3368 2416
rect -3438 -2416 -3368 -1984
rect -3272 1984 -3202 2416
rect -3272 -2416 -3202 -1984
rect -3106 1984 -3036 2416
rect -3106 -2416 -3036 -1984
rect -2940 1984 -2870 2416
rect -2940 -2416 -2870 -1984
rect -2774 1984 -2704 2416
rect -2774 -2416 -2704 -1984
rect -2608 1984 -2538 2416
rect -2608 -2416 -2538 -1984
rect -2442 1984 -2372 2416
rect -2442 -2416 -2372 -1984
rect -2276 1984 -2206 2416
rect -2276 -2416 -2206 -1984
rect -2110 1984 -2040 2416
rect -2110 -2416 -2040 -1984
rect -1944 1984 -1874 2416
rect -1944 -2416 -1874 -1984
rect -1778 1984 -1708 2416
rect -1778 -2416 -1708 -1984
rect -1612 1984 -1542 2416
rect -1612 -2416 -1542 -1984
rect -1446 1984 -1376 2416
rect -1446 -2416 -1376 -1984
rect -1280 1984 -1210 2416
rect -1280 -2416 -1210 -1984
rect -1114 1984 -1044 2416
rect -1114 -2416 -1044 -1984
rect -948 1984 -878 2416
rect -948 -2416 -878 -1984
rect -782 1984 -712 2416
rect -782 -2416 -712 -1984
rect -616 1984 -546 2416
rect -616 -2416 -546 -1984
rect -450 1984 -380 2416
rect -450 -2416 -380 -1984
rect -284 1984 -214 2416
rect -284 -2416 -214 -1984
rect -118 1984 -48 2416
rect -118 -2416 -48 -1984
rect 48 1984 118 2416
rect 48 -2416 118 -1984
rect 214 1984 284 2416
rect 214 -2416 284 -1984
rect 380 1984 450 2416
rect 380 -2416 450 -1984
rect 546 1984 616 2416
rect 546 -2416 616 -1984
rect 712 1984 782 2416
rect 712 -2416 782 -1984
rect 878 1984 948 2416
rect 878 -2416 948 -1984
rect 1044 1984 1114 2416
rect 1044 -2416 1114 -1984
rect 1210 1984 1280 2416
rect 1210 -2416 1280 -1984
rect 1376 1984 1446 2416
rect 1376 -2416 1446 -1984
rect 1542 1984 1612 2416
rect 1542 -2416 1612 -1984
rect 1708 1984 1778 2416
rect 1708 -2416 1778 -1984
rect 1874 1984 1944 2416
rect 1874 -2416 1944 -1984
rect 2040 1984 2110 2416
rect 2040 -2416 2110 -1984
rect 2206 1984 2276 2416
rect 2206 -2416 2276 -1984
rect 2372 1984 2442 2416
rect 2372 -2416 2442 -1984
rect 2538 1984 2608 2416
rect 2538 -2416 2608 -1984
rect 2704 1984 2774 2416
rect 2704 -2416 2774 -1984
rect 2870 1984 2940 2416
rect 2870 -2416 2940 -1984
rect 3036 1984 3106 2416
rect 3036 -2416 3106 -1984
rect 3202 1984 3272 2416
rect 3202 -2416 3272 -1984
rect 3368 1984 3438 2416
rect 3368 -2416 3438 -1984
rect 3534 1984 3604 2416
rect 3534 -2416 3604 -1984
rect 3700 1984 3770 2416
rect 3700 -2416 3770 -1984
rect 3866 1984 3936 2416
rect 3866 -2416 3936 -1984
rect 4032 1984 4102 2416
rect 4032 -2416 4102 -1984
rect 4198 1984 4268 2416
rect 4198 -2416 4268 -1984
rect 4364 1984 4434 2416
rect 4364 -2416 4434 -1984
rect 4530 1984 4600 2416
rect 4530 -2416 4600 -1984
rect 4696 1984 4766 2416
rect 4696 -2416 4766 -1984
rect 4862 1984 4932 2416
rect 4862 -2416 4932 -1984
rect 5028 1984 5098 2416
rect 5028 -2416 5098 -1984
rect 5194 1984 5264 2416
rect 5194 -2416 5264 -1984
<< xpolyres >>
rect -5264 -1984 -5194 1984
rect -5098 -1984 -5028 1984
rect -4932 -1984 -4862 1984
rect -4766 -1984 -4696 1984
rect -4600 -1984 -4530 1984
rect -4434 -1984 -4364 1984
rect -4268 -1984 -4198 1984
rect -4102 -1984 -4032 1984
rect -3936 -1984 -3866 1984
rect -3770 -1984 -3700 1984
rect -3604 -1984 -3534 1984
rect -3438 -1984 -3368 1984
rect -3272 -1984 -3202 1984
rect -3106 -1984 -3036 1984
rect -2940 -1984 -2870 1984
rect -2774 -1984 -2704 1984
rect -2608 -1984 -2538 1984
rect -2442 -1984 -2372 1984
rect -2276 -1984 -2206 1984
rect -2110 -1984 -2040 1984
rect -1944 -1984 -1874 1984
rect -1778 -1984 -1708 1984
rect -1612 -1984 -1542 1984
rect -1446 -1984 -1376 1984
rect -1280 -1984 -1210 1984
rect -1114 -1984 -1044 1984
rect -948 -1984 -878 1984
rect -782 -1984 -712 1984
rect -616 -1984 -546 1984
rect -450 -1984 -380 1984
rect -284 -1984 -214 1984
rect -118 -1984 -48 1984
rect 48 -1984 118 1984
rect 214 -1984 284 1984
rect 380 -1984 450 1984
rect 546 -1984 616 1984
rect 712 -1984 782 1984
rect 878 -1984 948 1984
rect 1044 -1984 1114 1984
rect 1210 -1984 1280 1984
rect 1376 -1984 1446 1984
rect 1542 -1984 1612 1984
rect 1708 -1984 1778 1984
rect 1874 -1984 1944 1984
rect 2040 -1984 2110 1984
rect 2206 -1984 2276 1984
rect 2372 -1984 2442 1984
rect 2538 -1984 2608 1984
rect 2704 -1984 2774 1984
rect 2870 -1984 2940 1984
rect 3036 -1984 3106 1984
rect 3202 -1984 3272 1984
rect 3368 -1984 3438 1984
rect 3534 -1984 3604 1984
rect 3700 -1984 3770 1984
rect 3866 -1984 3936 1984
rect 4032 -1984 4102 1984
rect 4198 -1984 4268 1984
rect 4364 -1984 4434 1984
rect 4530 -1984 4600 1984
rect 4696 -1984 4766 1984
rect 4862 -1984 4932 1984
rect 5028 -1984 5098 1984
rect 5194 -1984 5264 1984
<< locali >>
rect -5394 2512 -5298 2546
rect 5298 2512 5394 2546
rect -5394 2450 -5360 2512
rect 5360 2450 5394 2512
rect -5394 -2512 -5360 -2450
rect 5360 -2512 5394 -2450
rect -5394 -2546 -5298 -2512
rect 5298 -2546 5394 -2512
<< viali >>
rect -5248 2001 -5210 2398
rect -5082 2001 -5044 2398
rect -4916 2001 -4878 2398
rect -4750 2001 -4712 2398
rect -4584 2001 -4546 2398
rect -4418 2001 -4380 2398
rect -4252 2001 -4214 2398
rect -4086 2001 -4048 2398
rect -3920 2001 -3882 2398
rect -3754 2001 -3716 2398
rect -3588 2001 -3550 2398
rect -3422 2001 -3384 2398
rect -3256 2001 -3218 2398
rect -3090 2001 -3052 2398
rect -2924 2001 -2886 2398
rect -2758 2001 -2720 2398
rect -2592 2001 -2554 2398
rect -2426 2001 -2388 2398
rect -2260 2001 -2222 2398
rect -2094 2001 -2056 2398
rect -1928 2001 -1890 2398
rect -1762 2001 -1724 2398
rect -1596 2001 -1558 2398
rect -1430 2001 -1392 2398
rect -1264 2001 -1226 2398
rect -1098 2001 -1060 2398
rect -932 2001 -894 2398
rect -766 2001 -728 2398
rect -600 2001 -562 2398
rect -434 2001 -396 2398
rect -268 2001 -230 2398
rect -102 2001 -64 2398
rect 64 2001 102 2398
rect 230 2001 268 2398
rect 396 2001 434 2398
rect 562 2001 600 2398
rect 728 2001 766 2398
rect 894 2001 932 2398
rect 1060 2001 1098 2398
rect 1226 2001 1264 2398
rect 1392 2001 1430 2398
rect 1558 2001 1596 2398
rect 1724 2001 1762 2398
rect 1890 2001 1928 2398
rect 2056 2001 2094 2398
rect 2222 2001 2260 2398
rect 2388 2001 2426 2398
rect 2554 2001 2592 2398
rect 2720 2001 2758 2398
rect 2886 2001 2924 2398
rect 3052 2001 3090 2398
rect 3218 2001 3256 2398
rect 3384 2001 3422 2398
rect 3550 2001 3588 2398
rect 3716 2001 3754 2398
rect 3882 2001 3920 2398
rect 4048 2001 4086 2398
rect 4214 2001 4252 2398
rect 4380 2001 4418 2398
rect 4546 2001 4584 2398
rect 4712 2001 4750 2398
rect 4878 2001 4916 2398
rect 5044 2001 5082 2398
rect 5210 2001 5248 2398
rect -5248 -2398 -5210 -2001
rect -5082 -2398 -5044 -2001
rect -4916 -2398 -4878 -2001
rect -4750 -2398 -4712 -2001
rect -4584 -2398 -4546 -2001
rect -4418 -2398 -4380 -2001
rect -4252 -2398 -4214 -2001
rect -4086 -2398 -4048 -2001
rect -3920 -2398 -3882 -2001
rect -3754 -2398 -3716 -2001
rect -3588 -2398 -3550 -2001
rect -3422 -2398 -3384 -2001
rect -3256 -2398 -3218 -2001
rect -3090 -2398 -3052 -2001
rect -2924 -2398 -2886 -2001
rect -2758 -2398 -2720 -2001
rect -2592 -2398 -2554 -2001
rect -2426 -2398 -2388 -2001
rect -2260 -2398 -2222 -2001
rect -2094 -2398 -2056 -2001
rect -1928 -2398 -1890 -2001
rect -1762 -2398 -1724 -2001
rect -1596 -2398 -1558 -2001
rect -1430 -2398 -1392 -2001
rect -1264 -2398 -1226 -2001
rect -1098 -2398 -1060 -2001
rect -932 -2398 -894 -2001
rect -766 -2398 -728 -2001
rect -600 -2398 -562 -2001
rect -434 -2398 -396 -2001
rect -268 -2398 -230 -2001
rect -102 -2398 -64 -2001
rect 64 -2398 102 -2001
rect 230 -2398 268 -2001
rect 396 -2398 434 -2001
rect 562 -2398 600 -2001
rect 728 -2398 766 -2001
rect 894 -2398 932 -2001
rect 1060 -2398 1098 -2001
rect 1226 -2398 1264 -2001
rect 1392 -2398 1430 -2001
rect 1558 -2398 1596 -2001
rect 1724 -2398 1762 -2001
rect 1890 -2398 1928 -2001
rect 2056 -2398 2094 -2001
rect 2222 -2398 2260 -2001
rect 2388 -2398 2426 -2001
rect 2554 -2398 2592 -2001
rect 2720 -2398 2758 -2001
rect 2886 -2398 2924 -2001
rect 3052 -2398 3090 -2001
rect 3218 -2398 3256 -2001
rect 3384 -2398 3422 -2001
rect 3550 -2398 3588 -2001
rect 3716 -2398 3754 -2001
rect 3882 -2398 3920 -2001
rect 4048 -2398 4086 -2001
rect 4214 -2398 4252 -2001
rect 4380 -2398 4418 -2001
rect 4546 -2398 4584 -2001
rect 4712 -2398 4750 -2001
rect 4878 -2398 4916 -2001
rect 5044 -2398 5082 -2001
rect 5210 -2398 5248 -2001
<< metal1 >>
rect -5254 2398 -5204 2410
rect -5254 2001 -5248 2398
rect -5210 2001 -5204 2398
rect -5254 1989 -5204 2001
rect -5088 2398 -5038 2410
rect -5088 2001 -5082 2398
rect -5044 2001 -5038 2398
rect -5088 1989 -5038 2001
rect -4922 2398 -4872 2410
rect -4922 2001 -4916 2398
rect -4878 2001 -4872 2398
rect -4922 1989 -4872 2001
rect -4756 2398 -4706 2410
rect -4756 2001 -4750 2398
rect -4712 2001 -4706 2398
rect -4756 1989 -4706 2001
rect -4590 2398 -4540 2410
rect -4590 2001 -4584 2398
rect -4546 2001 -4540 2398
rect -4590 1989 -4540 2001
rect -4424 2398 -4374 2410
rect -4424 2001 -4418 2398
rect -4380 2001 -4374 2398
rect -4424 1989 -4374 2001
rect -4258 2398 -4208 2410
rect -4258 2001 -4252 2398
rect -4214 2001 -4208 2398
rect -4258 1989 -4208 2001
rect -4092 2398 -4042 2410
rect -4092 2001 -4086 2398
rect -4048 2001 -4042 2398
rect -4092 1989 -4042 2001
rect -3926 2398 -3876 2410
rect -3926 2001 -3920 2398
rect -3882 2001 -3876 2398
rect -3926 1989 -3876 2001
rect -3760 2398 -3710 2410
rect -3760 2001 -3754 2398
rect -3716 2001 -3710 2398
rect -3760 1989 -3710 2001
rect -3594 2398 -3544 2410
rect -3594 2001 -3588 2398
rect -3550 2001 -3544 2398
rect -3594 1989 -3544 2001
rect -3428 2398 -3378 2410
rect -3428 2001 -3422 2398
rect -3384 2001 -3378 2398
rect -3428 1989 -3378 2001
rect -3262 2398 -3212 2410
rect -3262 2001 -3256 2398
rect -3218 2001 -3212 2398
rect -3262 1989 -3212 2001
rect -3096 2398 -3046 2410
rect -3096 2001 -3090 2398
rect -3052 2001 -3046 2398
rect -3096 1989 -3046 2001
rect -2930 2398 -2880 2410
rect -2930 2001 -2924 2398
rect -2886 2001 -2880 2398
rect -2930 1989 -2880 2001
rect -2764 2398 -2714 2410
rect -2764 2001 -2758 2398
rect -2720 2001 -2714 2398
rect -2764 1989 -2714 2001
rect -2598 2398 -2548 2410
rect -2598 2001 -2592 2398
rect -2554 2001 -2548 2398
rect -2598 1989 -2548 2001
rect -2432 2398 -2382 2410
rect -2432 2001 -2426 2398
rect -2388 2001 -2382 2398
rect -2432 1989 -2382 2001
rect -2266 2398 -2216 2410
rect -2266 2001 -2260 2398
rect -2222 2001 -2216 2398
rect -2266 1989 -2216 2001
rect -2100 2398 -2050 2410
rect -2100 2001 -2094 2398
rect -2056 2001 -2050 2398
rect -2100 1989 -2050 2001
rect -1934 2398 -1884 2410
rect -1934 2001 -1928 2398
rect -1890 2001 -1884 2398
rect -1934 1989 -1884 2001
rect -1768 2398 -1718 2410
rect -1768 2001 -1762 2398
rect -1724 2001 -1718 2398
rect -1768 1989 -1718 2001
rect -1602 2398 -1552 2410
rect -1602 2001 -1596 2398
rect -1558 2001 -1552 2398
rect -1602 1989 -1552 2001
rect -1436 2398 -1386 2410
rect -1436 2001 -1430 2398
rect -1392 2001 -1386 2398
rect -1436 1989 -1386 2001
rect -1270 2398 -1220 2410
rect -1270 2001 -1264 2398
rect -1226 2001 -1220 2398
rect -1270 1989 -1220 2001
rect -1104 2398 -1054 2410
rect -1104 2001 -1098 2398
rect -1060 2001 -1054 2398
rect -1104 1989 -1054 2001
rect -938 2398 -888 2410
rect -938 2001 -932 2398
rect -894 2001 -888 2398
rect -938 1989 -888 2001
rect -772 2398 -722 2410
rect -772 2001 -766 2398
rect -728 2001 -722 2398
rect -772 1989 -722 2001
rect -606 2398 -556 2410
rect -606 2001 -600 2398
rect -562 2001 -556 2398
rect -606 1989 -556 2001
rect -440 2398 -390 2410
rect -440 2001 -434 2398
rect -396 2001 -390 2398
rect -440 1989 -390 2001
rect -274 2398 -224 2410
rect -274 2001 -268 2398
rect -230 2001 -224 2398
rect -274 1989 -224 2001
rect -108 2398 -58 2410
rect -108 2001 -102 2398
rect -64 2001 -58 2398
rect -108 1989 -58 2001
rect 58 2398 108 2410
rect 58 2001 64 2398
rect 102 2001 108 2398
rect 58 1989 108 2001
rect 224 2398 274 2410
rect 224 2001 230 2398
rect 268 2001 274 2398
rect 224 1989 274 2001
rect 390 2398 440 2410
rect 390 2001 396 2398
rect 434 2001 440 2398
rect 390 1989 440 2001
rect 556 2398 606 2410
rect 556 2001 562 2398
rect 600 2001 606 2398
rect 556 1989 606 2001
rect 722 2398 772 2410
rect 722 2001 728 2398
rect 766 2001 772 2398
rect 722 1989 772 2001
rect 888 2398 938 2410
rect 888 2001 894 2398
rect 932 2001 938 2398
rect 888 1989 938 2001
rect 1054 2398 1104 2410
rect 1054 2001 1060 2398
rect 1098 2001 1104 2398
rect 1054 1989 1104 2001
rect 1220 2398 1270 2410
rect 1220 2001 1226 2398
rect 1264 2001 1270 2398
rect 1220 1989 1270 2001
rect 1386 2398 1436 2410
rect 1386 2001 1392 2398
rect 1430 2001 1436 2398
rect 1386 1989 1436 2001
rect 1552 2398 1602 2410
rect 1552 2001 1558 2398
rect 1596 2001 1602 2398
rect 1552 1989 1602 2001
rect 1718 2398 1768 2410
rect 1718 2001 1724 2398
rect 1762 2001 1768 2398
rect 1718 1989 1768 2001
rect 1884 2398 1934 2410
rect 1884 2001 1890 2398
rect 1928 2001 1934 2398
rect 1884 1989 1934 2001
rect 2050 2398 2100 2410
rect 2050 2001 2056 2398
rect 2094 2001 2100 2398
rect 2050 1989 2100 2001
rect 2216 2398 2266 2410
rect 2216 2001 2222 2398
rect 2260 2001 2266 2398
rect 2216 1989 2266 2001
rect 2382 2398 2432 2410
rect 2382 2001 2388 2398
rect 2426 2001 2432 2398
rect 2382 1989 2432 2001
rect 2548 2398 2598 2410
rect 2548 2001 2554 2398
rect 2592 2001 2598 2398
rect 2548 1989 2598 2001
rect 2714 2398 2764 2410
rect 2714 2001 2720 2398
rect 2758 2001 2764 2398
rect 2714 1989 2764 2001
rect 2880 2398 2930 2410
rect 2880 2001 2886 2398
rect 2924 2001 2930 2398
rect 2880 1989 2930 2001
rect 3046 2398 3096 2410
rect 3046 2001 3052 2398
rect 3090 2001 3096 2398
rect 3046 1989 3096 2001
rect 3212 2398 3262 2410
rect 3212 2001 3218 2398
rect 3256 2001 3262 2398
rect 3212 1989 3262 2001
rect 3378 2398 3428 2410
rect 3378 2001 3384 2398
rect 3422 2001 3428 2398
rect 3378 1989 3428 2001
rect 3544 2398 3594 2410
rect 3544 2001 3550 2398
rect 3588 2001 3594 2398
rect 3544 1989 3594 2001
rect 3710 2398 3760 2410
rect 3710 2001 3716 2398
rect 3754 2001 3760 2398
rect 3710 1989 3760 2001
rect 3876 2398 3926 2410
rect 3876 2001 3882 2398
rect 3920 2001 3926 2398
rect 3876 1989 3926 2001
rect 4042 2398 4092 2410
rect 4042 2001 4048 2398
rect 4086 2001 4092 2398
rect 4042 1989 4092 2001
rect 4208 2398 4258 2410
rect 4208 2001 4214 2398
rect 4252 2001 4258 2398
rect 4208 1989 4258 2001
rect 4374 2398 4424 2410
rect 4374 2001 4380 2398
rect 4418 2001 4424 2398
rect 4374 1989 4424 2001
rect 4540 2398 4590 2410
rect 4540 2001 4546 2398
rect 4584 2001 4590 2398
rect 4540 1989 4590 2001
rect 4706 2398 4756 2410
rect 4706 2001 4712 2398
rect 4750 2001 4756 2398
rect 4706 1989 4756 2001
rect 4872 2398 4922 2410
rect 4872 2001 4878 2398
rect 4916 2001 4922 2398
rect 4872 1989 4922 2001
rect 5038 2398 5088 2410
rect 5038 2001 5044 2398
rect 5082 2001 5088 2398
rect 5038 1989 5088 2001
rect 5204 2398 5254 2410
rect 5204 2001 5210 2398
rect 5248 2001 5254 2398
rect 5204 1989 5254 2001
rect -5254 -2001 -5204 -1989
rect -5254 -2398 -5248 -2001
rect -5210 -2398 -5204 -2001
rect -5254 -2410 -5204 -2398
rect -5088 -2001 -5038 -1989
rect -5088 -2398 -5082 -2001
rect -5044 -2398 -5038 -2001
rect -5088 -2410 -5038 -2398
rect -4922 -2001 -4872 -1989
rect -4922 -2398 -4916 -2001
rect -4878 -2398 -4872 -2001
rect -4922 -2410 -4872 -2398
rect -4756 -2001 -4706 -1989
rect -4756 -2398 -4750 -2001
rect -4712 -2398 -4706 -2001
rect -4756 -2410 -4706 -2398
rect -4590 -2001 -4540 -1989
rect -4590 -2398 -4584 -2001
rect -4546 -2398 -4540 -2001
rect -4590 -2410 -4540 -2398
rect -4424 -2001 -4374 -1989
rect -4424 -2398 -4418 -2001
rect -4380 -2398 -4374 -2001
rect -4424 -2410 -4374 -2398
rect -4258 -2001 -4208 -1989
rect -4258 -2398 -4252 -2001
rect -4214 -2398 -4208 -2001
rect -4258 -2410 -4208 -2398
rect -4092 -2001 -4042 -1989
rect -4092 -2398 -4086 -2001
rect -4048 -2398 -4042 -2001
rect -4092 -2410 -4042 -2398
rect -3926 -2001 -3876 -1989
rect -3926 -2398 -3920 -2001
rect -3882 -2398 -3876 -2001
rect -3926 -2410 -3876 -2398
rect -3760 -2001 -3710 -1989
rect -3760 -2398 -3754 -2001
rect -3716 -2398 -3710 -2001
rect -3760 -2410 -3710 -2398
rect -3594 -2001 -3544 -1989
rect -3594 -2398 -3588 -2001
rect -3550 -2398 -3544 -2001
rect -3594 -2410 -3544 -2398
rect -3428 -2001 -3378 -1989
rect -3428 -2398 -3422 -2001
rect -3384 -2398 -3378 -2001
rect -3428 -2410 -3378 -2398
rect -3262 -2001 -3212 -1989
rect -3262 -2398 -3256 -2001
rect -3218 -2398 -3212 -2001
rect -3262 -2410 -3212 -2398
rect -3096 -2001 -3046 -1989
rect -3096 -2398 -3090 -2001
rect -3052 -2398 -3046 -2001
rect -3096 -2410 -3046 -2398
rect -2930 -2001 -2880 -1989
rect -2930 -2398 -2924 -2001
rect -2886 -2398 -2880 -2001
rect -2930 -2410 -2880 -2398
rect -2764 -2001 -2714 -1989
rect -2764 -2398 -2758 -2001
rect -2720 -2398 -2714 -2001
rect -2764 -2410 -2714 -2398
rect -2598 -2001 -2548 -1989
rect -2598 -2398 -2592 -2001
rect -2554 -2398 -2548 -2001
rect -2598 -2410 -2548 -2398
rect -2432 -2001 -2382 -1989
rect -2432 -2398 -2426 -2001
rect -2388 -2398 -2382 -2001
rect -2432 -2410 -2382 -2398
rect -2266 -2001 -2216 -1989
rect -2266 -2398 -2260 -2001
rect -2222 -2398 -2216 -2001
rect -2266 -2410 -2216 -2398
rect -2100 -2001 -2050 -1989
rect -2100 -2398 -2094 -2001
rect -2056 -2398 -2050 -2001
rect -2100 -2410 -2050 -2398
rect -1934 -2001 -1884 -1989
rect -1934 -2398 -1928 -2001
rect -1890 -2398 -1884 -2001
rect -1934 -2410 -1884 -2398
rect -1768 -2001 -1718 -1989
rect -1768 -2398 -1762 -2001
rect -1724 -2398 -1718 -2001
rect -1768 -2410 -1718 -2398
rect -1602 -2001 -1552 -1989
rect -1602 -2398 -1596 -2001
rect -1558 -2398 -1552 -2001
rect -1602 -2410 -1552 -2398
rect -1436 -2001 -1386 -1989
rect -1436 -2398 -1430 -2001
rect -1392 -2398 -1386 -2001
rect -1436 -2410 -1386 -2398
rect -1270 -2001 -1220 -1989
rect -1270 -2398 -1264 -2001
rect -1226 -2398 -1220 -2001
rect -1270 -2410 -1220 -2398
rect -1104 -2001 -1054 -1989
rect -1104 -2398 -1098 -2001
rect -1060 -2398 -1054 -2001
rect -1104 -2410 -1054 -2398
rect -938 -2001 -888 -1989
rect -938 -2398 -932 -2001
rect -894 -2398 -888 -2001
rect -938 -2410 -888 -2398
rect -772 -2001 -722 -1989
rect -772 -2398 -766 -2001
rect -728 -2398 -722 -2001
rect -772 -2410 -722 -2398
rect -606 -2001 -556 -1989
rect -606 -2398 -600 -2001
rect -562 -2398 -556 -2001
rect -606 -2410 -556 -2398
rect -440 -2001 -390 -1989
rect -440 -2398 -434 -2001
rect -396 -2398 -390 -2001
rect -440 -2410 -390 -2398
rect -274 -2001 -224 -1989
rect -274 -2398 -268 -2001
rect -230 -2398 -224 -2001
rect -274 -2410 -224 -2398
rect -108 -2001 -58 -1989
rect -108 -2398 -102 -2001
rect -64 -2398 -58 -2001
rect -108 -2410 -58 -2398
rect 58 -2001 108 -1989
rect 58 -2398 64 -2001
rect 102 -2398 108 -2001
rect 58 -2410 108 -2398
rect 224 -2001 274 -1989
rect 224 -2398 230 -2001
rect 268 -2398 274 -2001
rect 224 -2410 274 -2398
rect 390 -2001 440 -1989
rect 390 -2398 396 -2001
rect 434 -2398 440 -2001
rect 390 -2410 440 -2398
rect 556 -2001 606 -1989
rect 556 -2398 562 -2001
rect 600 -2398 606 -2001
rect 556 -2410 606 -2398
rect 722 -2001 772 -1989
rect 722 -2398 728 -2001
rect 766 -2398 772 -2001
rect 722 -2410 772 -2398
rect 888 -2001 938 -1989
rect 888 -2398 894 -2001
rect 932 -2398 938 -2001
rect 888 -2410 938 -2398
rect 1054 -2001 1104 -1989
rect 1054 -2398 1060 -2001
rect 1098 -2398 1104 -2001
rect 1054 -2410 1104 -2398
rect 1220 -2001 1270 -1989
rect 1220 -2398 1226 -2001
rect 1264 -2398 1270 -2001
rect 1220 -2410 1270 -2398
rect 1386 -2001 1436 -1989
rect 1386 -2398 1392 -2001
rect 1430 -2398 1436 -2001
rect 1386 -2410 1436 -2398
rect 1552 -2001 1602 -1989
rect 1552 -2398 1558 -2001
rect 1596 -2398 1602 -2001
rect 1552 -2410 1602 -2398
rect 1718 -2001 1768 -1989
rect 1718 -2398 1724 -2001
rect 1762 -2398 1768 -2001
rect 1718 -2410 1768 -2398
rect 1884 -2001 1934 -1989
rect 1884 -2398 1890 -2001
rect 1928 -2398 1934 -2001
rect 1884 -2410 1934 -2398
rect 2050 -2001 2100 -1989
rect 2050 -2398 2056 -2001
rect 2094 -2398 2100 -2001
rect 2050 -2410 2100 -2398
rect 2216 -2001 2266 -1989
rect 2216 -2398 2222 -2001
rect 2260 -2398 2266 -2001
rect 2216 -2410 2266 -2398
rect 2382 -2001 2432 -1989
rect 2382 -2398 2388 -2001
rect 2426 -2398 2432 -2001
rect 2382 -2410 2432 -2398
rect 2548 -2001 2598 -1989
rect 2548 -2398 2554 -2001
rect 2592 -2398 2598 -2001
rect 2548 -2410 2598 -2398
rect 2714 -2001 2764 -1989
rect 2714 -2398 2720 -2001
rect 2758 -2398 2764 -2001
rect 2714 -2410 2764 -2398
rect 2880 -2001 2930 -1989
rect 2880 -2398 2886 -2001
rect 2924 -2398 2930 -2001
rect 2880 -2410 2930 -2398
rect 3046 -2001 3096 -1989
rect 3046 -2398 3052 -2001
rect 3090 -2398 3096 -2001
rect 3046 -2410 3096 -2398
rect 3212 -2001 3262 -1989
rect 3212 -2398 3218 -2001
rect 3256 -2398 3262 -2001
rect 3212 -2410 3262 -2398
rect 3378 -2001 3428 -1989
rect 3378 -2398 3384 -2001
rect 3422 -2398 3428 -2001
rect 3378 -2410 3428 -2398
rect 3544 -2001 3594 -1989
rect 3544 -2398 3550 -2001
rect 3588 -2398 3594 -2001
rect 3544 -2410 3594 -2398
rect 3710 -2001 3760 -1989
rect 3710 -2398 3716 -2001
rect 3754 -2398 3760 -2001
rect 3710 -2410 3760 -2398
rect 3876 -2001 3926 -1989
rect 3876 -2398 3882 -2001
rect 3920 -2398 3926 -2001
rect 3876 -2410 3926 -2398
rect 4042 -2001 4092 -1989
rect 4042 -2398 4048 -2001
rect 4086 -2398 4092 -2001
rect 4042 -2410 4092 -2398
rect 4208 -2001 4258 -1989
rect 4208 -2398 4214 -2001
rect 4252 -2398 4258 -2001
rect 4208 -2410 4258 -2398
rect 4374 -2001 4424 -1989
rect 4374 -2398 4380 -2001
rect 4418 -2398 4424 -2001
rect 4374 -2410 4424 -2398
rect 4540 -2001 4590 -1989
rect 4540 -2398 4546 -2001
rect 4584 -2398 4590 -2001
rect 4540 -2410 4590 -2398
rect 4706 -2001 4756 -1989
rect 4706 -2398 4712 -2001
rect 4750 -2398 4756 -2001
rect 4706 -2410 4756 -2398
rect 4872 -2001 4922 -1989
rect 4872 -2398 4878 -2001
rect 4916 -2398 4922 -2001
rect 4872 -2410 4922 -2398
rect 5038 -2001 5088 -1989
rect 5038 -2398 5044 -2001
rect 5082 -2398 5088 -2001
rect 5038 -2410 5088 -2398
rect 5204 -2001 5254 -1989
rect 5204 -2398 5210 -2001
rect 5248 -2398 5254 -2001
rect 5204 -2410 5254 -2398
<< properties >>
string FIXED_BBOX -5377 -2529 5377 2529
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 20 m 1 nx 64 wmin 0.350 lmin 0.50 class resistor rho 2000 val 115.361k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
