magic
tech sky130A
magscale 1 2
timestamp 1730992408
<< nwell >>
rect -1225 -4337 1225 4337
<< pmoslvt >>
rect -1029 118 -29 4118
rect 29 118 1029 4118
rect -1029 -4118 -29 -118
rect 29 -4118 1029 -118
<< pdiff >>
rect -1087 4106 -1029 4118
rect -1087 130 -1075 4106
rect -1041 130 -1029 4106
rect -1087 118 -1029 130
rect -29 4106 29 4118
rect -29 130 -17 4106
rect 17 130 29 4106
rect -29 118 29 130
rect 1029 4106 1087 4118
rect 1029 130 1041 4106
rect 1075 130 1087 4106
rect 1029 118 1087 130
rect -1087 -130 -1029 -118
rect -1087 -4106 -1075 -130
rect -1041 -4106 -1029 -130
rect -1087 -4118 -1029 -4106
rect -29 -130 29 -118
rect -29 -4106 -17 -130
rect 17 -4106 29 -130
rect -29 -4118 29 -4106
rect 1029 -130 1087 -118
rect 1029 -4106 1041 -130
rect 1075 -4106 1087 -130
rect 1029 -4118 1087 -4106
<< pdiffc >>
rect -1075 130 -1041 4106
rect -17 130 17 4106
rect 1041 130 1075 4106
rect -1075 -4106 -1041 -130
rect -17 -4106 17 -130
rect 1041 -4106 1075 -130
<< nsubdiff >>
rect -1189 4267 -1093 4301
rect 1093 4267 1189 4301
rect -1189 4205 -1155 4267
rect 1155 4205 1189 4267
rect -1189 -4267 -1155 -4205
rect 1155 -4267 1189 -4205
rect -1189 -4301 -1093 -4267
rect 1093 -4301 1189 -4267
<< nsubdiffcont >>
rect -1093 4267 1093 4301
rect -1189 -4205 -1155 4205
rect 1155 -4205 1189 4205
rect -1093 -4301 1093 -4267
<< poly >>
rect -1029 4199 -29 4215
rect -1029 4165 -1013 4199
rect -45 4165 -29 4199
rect -1029 4118 -29 4165
rect 29 4199 1029 4215
rect 29 4165 45 4199
rect 1013 4165 1029 4199
rect 29 4118 1029 4165
rect -1029 71 -29 118
rect -1029 37 -1013 71
rect -45 37 -29 71
rect -1029 21 -29 37
rect 29 71 1029 118
rect 29 37 45 71
rect 1013 37 1029 71
rect 29 21 1029 37
rect -1029 -37 -29 -21
rect -1029 -71 -1013 -37
rect -45 -71 -29 -37
rect -1029 -118 -29 -71
rect 29 -37 1029 -21
rect 29 -71 45 -37
rect 1013 -71 1029 -37
rect 29 -118 1029 -71
rect -1029 -4165 -29 -4118
rect -1029 -4199 -1013 -4165
rect -45 -4199 -29 -4165
rect -1029 -4215 -29 -4199
rect 29 -4165 1029 -4118
rect 29 -4199 45 -4165
rect 1013 -4199 1029 -4165
rect 29 -4215 1029 -4199
<< polycont >>
rect -1013 4165 -45 4199
rect 45 4165 1013 4199
rect -1013 37 -45 71
rect 45 37 1013 71
rect -1013 -71 -45 -37
rect 45 -71 1013 -37
rect -1013 -4199 -45 -4165
rect 45 -4199 1013 -4165
<< locali >>
rect -1189 4267 -1093 4301
rect 1093 4267 1189 4301
rect -1189 4205 -1155 4267
rect 1155 4205 1189 4267
rect -1029 4165 -1013 4199
rect -45 4165 -29 4199
rect 29 4165 45 4199
rect 1013 4165 1029 4199
rect -1075 4106 -1041 4122
rect -1075 114 -1041 130
rect -17 4106 17 4122
rect -17 114 17 130
rect 1041 4106 1075 4122
rect 1041 114 1075 130
rect -1029 37 -1013 71
rect -45 37 -29 71
rect 29 37 45 71
rect 1013 37 1029 71
rect -1029 -71 -1013 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 1013 -71 1029 -37
rect -1075 -130 -1041 -114
rect -1075 -4122 -1041 -4106
rect -17 -130 17 -114
rect -17 -4122 17 -4106
rect 1041 -130 1075 -114
rect 1041 -4122 1075 -4106
rect -1029 -4199 -1013 -4165
rect -45 -4199 -29 -4165
rect 29 -4199 45 -4165
rect 1013 -4199 1029 -4165
rect -1189 -4267 -1155 -4205
rect 1155 -4267 1189 -4205
rect -1189 -4301 -1093 -4267
rect 1093 -4301 1189 -4267
<< viali >>
rect -1013 4165 -45 4199
rect 45 4165 1013 4199
rect -1075 130 -1041 4106
rect -17 130 17 4106
rect 1041 130 1075 4106
rect -1013 37 -45 71
rect 45 37 1013 71
rect -1013 -71 -45 -37
rect 45 -71 1013 -37
rect -1075 -4106 -1041 -130
rect -17 -4106 17 -130
rect 1041 -4106 1075 -130
rect -1013 -4199 -45 -4165
rect 45 -4199 1013 -4165
<< metal1 >>
rect -1025 4199 -33 4205
rect -1025 4165 -1013 4199
rect -45 4165 -33 4199
rect -1025 4159 -33 4165
rect 33 4199 1025 4205
rect 33 4165 45 4199
rect 1013 4165 1025 4199
rect 33 4159 1025 4165
rect -1081 4106 -1035 4118
rect -1081 130 -1075 4106
rect -1041 130 -1035 4106
rect -1081 118 -1035 130
rect -23 4106 23 4118
rect -23 130 -17 4106
rect 17 130 23 4106
rect -23 118 23 130
rect 1035 4106 1081 4118
rect 1035 130 1041 4106
rect 1075 130 1081 4106
rect 1035 118 1081 130
rect -1025 71 -33 77
rect -1025 37 -1013 71
rect -45 37 -33 71
rect -1025 31 -33 37
rect 33 71 1025 77
rect 33 37 45 71
rect 1013 37 1025 71
rect 33 31 1025 37
rect -1025 -37 -33 -31
rect -1025 -71 -1013 -37
rect -45 -71 -33 -37
rect -1025 -77 -33 -71
rect 33 -37 1025 -31
rect 33 -71 45 -37
rect 1013 -71 1025 -37
rect 33 -77 1025 -71
rect -1081 -130 -1035 -118
rect -1081 -4106 -1075 -130
rect -1041 -4106 -1035 -130
rect -1081 -4118 -1035 -4106
rect -23 -130 23 -118
rect -23 -4106 -17 -130
rect 17 -4106 23 -130
rect -23 -4118 23 -4106
rect 1035 -130 1081 -118
rect 1035 -4106 1041 -130
rect 1075 -4106 1081 -130
rect 1035 -4118 1081 -4106
rect -1025 -4165 -33 -4159
rect -1025 -4199 -1013 -4165
rect -45 -4199 -33 -4165
rect -1025 -4205 -33 -4199
rect 33 -4165 1025 -4159
rect 33 -4199 45 -4165
rect 1013 -4199 1025 -4165
rect 33 -4205 1025 -4199
<< properties >>
string FIXED_BBOX -1172 -4284 1172 4284
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 20.0 l 5.0 m 2 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
