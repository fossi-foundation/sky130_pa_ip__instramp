magic
tech sky130A
magscale 1 2
timestamp 1748311075
<< error_s >>
rect 548 8115 15090 8401
rect 548 1490 834 8115
rect 14804 8016 15090 8115
rect 548 -1152 752 1490
rect 15010 -658 15090 8016
rect 14110 -946 15090 -658
rect 4218 -952 7480 -946
rect 8686 -952 11948 -946
rect 12142 -1152 15090 -946
rect 548 -1232 15090 -1152
<< dnwell >>
rect 628 -1152 15010 8321
<< nwell >>
rect 3870 1538 12142 1706
rect 3870 -952 4218 1538
rect 7480 1488 8686 1538
rect 7480 -902 7708 1488
rect 8448 -902 8686 1488
rect 7480 -952 8686 -902
rect 11948 -952 12142 1538
rect 3870 -1104 12142 -952
rect 752 -1152 12142 -1104
<< mvnsubdiff >>
rect 12014 1442 12056 1466
rect 4074 1356 4152 1396
rect 4074 -826 4152 -786
rect 7546 1394 7620 1434
rect 8534 1398 8612 1438
rect 7546 -888 7620 -808
rect 8534 -884 8612 -804
rect 12014 -864 12056 -824
rect 4066 -1028 7510 -1018
rect 4066 -1074 4100 -1028
rect 7486 -1074 7510 -1028
rect 4066 -1086 7510 -1074
rect 8654 -1028 12074 -1018
rect 8654 -1074 8678 -1028
rect 12050 -1074 12074 -1028
rect 8654 -1086 12074 -1074
<< mvnsubdiffcont >>
rect 4074 -786 4152 1356
rect 7546 -808 7620 1394
rect 8534 -804 8612 1398
rect 12014 -824 12056 1442
rect 4100 -1074 7486 -1028
rect 8678 -1074 12050 -1028
<< poly >>
rect 7940 1170 8006 1236
rect 8142 1170 8224 1236
rect 7932 -440 8014 -374
rect 8150 -440 8216 -374
<< locali >>
rect 6146 8282 12396 8286
rect 6146 8240 6164 8282
rect 12380 8240 12396 8282
rect 6146 8228 12396 8240
rect 6148 2444 12434 2460
rect 6148 2386 6184 2444
rect 12402 2386 12434 2444
rect 6148 2338 12434 2386
rect 1878 2266 11362 2296
rect 1878 2194 1918 2266
rect 11306 2194 11362 2266
rect 1878 2162 11362 2194
rect 1878 1818 2004 2162
rect 11238 1818 11362 2162
rect 1878 1788 11362 1818
rect 1878 1716 1922 1788
rect 11310 1716 11362 1788
rect 1878 1684 11362 1716
rect 778 1412 866 1426
rect 3750 1412 3838 1424
rect 778 1396 3838 1412
rect 4288 1412 4352 1444
rect 778 1356 866 1396
rect 3746 1356 3838 1396
rect 778 1338 3838 1356
rect 778 1294 866 1338
rect 778 -904 806 1294
rect 852 -904 866 1294
rect 1138 -798 1254 1192
rect 1416 -798 1532 1192
rect 1694 -798 1810 1192
rect 1972 -798 2088 1192
rect 2250 -798 2366 1192
rect 2528 -798 2644 1192
rect 2806 -798 2922 1192
rect 3084 -798 3200 1192
rect 3362 -798 3478 1192
rect 3750 1182 3838 1338
rect 3750 -790 3768 1182
rect 3814 -790 3838 1182
rect 778 -956 866 -904
rect 3750 -956 3838 -790
rect 778 -974 3838 -956
rect 778 -1014 866 -974
rect 3746 -1014 3838 -974
rect 778 -1028 3838 -1014
rect 832 -1030 3838 -1028
rect 4060 1356 4170 1402
rect 4060 -786 4074 1356
rect 4152 -786 4170 1356
rect 4060 -1012 4170 -786
rect 4288 770 4300 1412
rect 4340 770 4352 1412
rect 4288 734 4352 770
rect 7352 1412 7416 1444
rect 7352 770 7364 1412
rect 7404 770 7416 1412
rect 4288 724 4364 734
rect 7352 732 7416 770
rect 4288 528 4308 724
rect 4346 528 4364 724
rect 4288 520 4364 528
rect 7338 726 7416 732
rect 7338 528 7348 726
rect 7388 528 7416 726
rect 7338 520 7416 528
rect 4288 482 4352 520
rect 4288 -856 4302 482
rect 4342 -812 4352 482
rect 7352 482 7416 520
rect 7352 -812 7364 482
rect 4342 -830 7364 -812
rect 4342 -856 4410 -830
rect 4288 -872 4410 -856
rect 7290 -856 7364 -830
rect 7404 -856 7416 482
rect 7290 -872 7416 -856
rect 4288 -884 7416 -872
rect 7534 1394 7644 1510
rect 7534 -808 7542 1394
rect 7620 -808 7644 1394
rect 7798 1404 8358 1432
rect 7798 1334 7834 1404
rect 8322 1334 8358 1404
rect 7798 1282 8358 1334
rect 8522 1398 8632 1490
rect 8142 1186 8156 1220
rect 8210 1186 8224 1220
rect 7778 428 7828 434
rect 7778 228 7794 428
rect 7778 220 7828 228
rect 7932 -424 7944 -390
rect 8002 -424 8014 -390
rect 7796 -540 8356 -488
rect 7796 -610 7830 -540
rect 8318 -610 8356 -540
rect 7796 -638 8356 -610
rect 7534 -944 7644 -808
rect 8522 -804 8534 1398
rect 8612 -804 8632 1398
rect 8522 -944 8632 -804
rect 8754 1420 8824 1446
rect 8754 1086 8768 1420
rect 8812 1086 8824 1420
rect 8754 1028 8824 1086
rect 8754 828 8778 1028
rect 8818 828 8824 1028
rect 8754 778 8824 828
rect 8754 -812 8768 778
rect 8810 -812 8824 778
rect 11810 1402 11880 1452
rect 11810 1068 11822 1402
rect 11866 1068 11880 1402
rect 11810 1028 11880 1068
rect 11810 830 11818 1028
rect 11858 830 11880 1028
rect 11810 776 11880 830
rect 11810 -812 11822 776
rect 8754 -814 11822 -812
rect 11864 -814 11880 776
rect 8754 -828 11880 -814
rect 8754 -866 8872 -828
rect 11768 -866 11880 -828
rect 8754 -880 11880 -866
rect 11974 1442 12074 1522
rect 11974 1416 12014 1442
rect 12056 1416 12074 1442
rect 11974 -826 11984 1416
rect 12062 -826 12074 1416
rect 7534 -1012 8632 -944
rect 4060 -1014 8632 -1012
rect 11974 -1014 12074 -826
rect 4060 -1018 12074 -1014
rect 4060 -1028 4102 -1018
rect 7506 -1020 12074 -1018
rect 4060 -1074 4100 -1028
rect 7506 -1038 8674 -1020
rect 7506 -1068 7644 -1038
rect 7486 -1074 7644 -1068
rect 4060 -1086 7644 -1074
rect 8518 -1070 8674 -1038
rect 8518 -1074 8678 -1070
rect 12050 -1074 12074 -1020
rect 8518 -1088 12074 -1074
<< viali >>
rect 6164 8240 12380 8282
rect 6147 2509 6181 8177
rect 12348 7074 12384 8042
rect 12692 7946 14878 7980
rect 12348 5964 12384 6932
rect 12348 4856 12384 5824
rect 12348 3748 12384 4716
rect 12348 2634 12384 3602
rect 6184 2386 12402 2444
rect 1918 2194 11306 2266
rect 1922 1716 11310 1788
rect 866 1356 3746 1396
rect 806 -904 852 1294
rect 3768 -790 3814 1182
rect 866 -1014 3746 -974
rect 4074 -786 4152 1356
rect 4300 770 4340 1412
rect 7364 770 7404 1412
rect 4308 528 4346 724
rect 7348 528 7388 726
rect 4302 -856 4342 482
rect 4410 -872 7290 -830
rect 7364 -856 7404 482
rect 7542 -808 7546 1394
rect 7546 -808 7620 1394
rect 7834 1334 8322 1404
rect 8156 1186 8210 1220
rect 7794 228 7830 428
rect 8328 222 8362 434
rect 7944 -424 8002 -390
rect 7830 -610 8318 -540
rect 8534 -804 8612 1398
rect 8768 1086 8812 1420
rect 8778 828 8818 1028
rect 8768 -812 8810 778
rect 11822 1068 11866 1402
rect 11818 830 11858 1028
rect 11822 -814 11864 776
rect 8872 -866 11768 -828
rect 11984 -824 12014 1416
rect 12014 -824 12056 1416
rect 12056 -824 12062 1416
rect 11984 -826 12062 -824
rect 12596 -526 12630 7884
rect 14940 -526 14974 7884
rect 12692 -622 14878 -588
rect 4102 -1028 7506 -1018
rect 4102 -1068 7486 -1028
rect 7486 -1068 7506 -1028
rect 8674 -1028 12050 -1020
rect 8674 -1070 8678 -1028
rect 8678 -1070 12050 -1028
<< metal1 >>
rect 6132 8282 12398 8288
rect 6132 8240 6164 8282
rect 12380 8240 12398 8282
rect 6132 8220 6178 8240
rect 12314 8220 12398 8240
rect 6132 8210 12398 8220
rect 6132 8177 6196 8210
rect 6132 2509 6147 8177
rect 6181 2509 6196 8177
rect 12482 8140 12682 8308
rect 6330 8108 12682 8140
rect 6330 8094 12548 8108
rect 6258 8058 6336 8064
rect 6258 7590 6264 8058
rect 6330 7590 6336 8058
rect 6258 7584 6336 7590
rect 6774 8058 6852 8064
rect 6774 7590 6780 8058
rect 6846 7590 6852 8058
rect 6774 7584 6852 7590
rect 7290 8058 7368 8064
rect 7290 7590 7296 8058
rect 7362 7590 7368 8058
rect 7290 7584 7368 7590
rect 7806 8058 7884 8064
rect 7806 7590 7812 8058
rect 7878 7590 7884 8058
rect 7806 7584 7884 7590
rect 8322 8058 8400 8064
rect 8322 7590 8328 8058
rect 8394 7590 8400 8058
rect 8322 7584 8400 7590
rect 8838 8058 8916 8064
rect 8838 7590 8844 8058
rect 8910 7590 8916 8058
rect 8838 7584 8916 7590
rect 9354 8058 9432 8064
rect 9354 7590 9360 8058
rect 9426 7590 9432 8058
rect 9354 7584 9432 7590
rect 9870 8058 9948 8064
rect 9870 7590 9876 8058
rect 9942 7590 9948 8058
rect 9870 7584 9948 7590
rect 10386 8058 10464 8064
rect 10386 7590 10392 8058
rect 10458 7590 10464 8058
rect 10386 7584 10464 7590
rect 10902 8058 10980 8064
rect 10902 7590 10908 8058
rect 10974 7590 10980 8058
rect 10902 7584 10980 7590
rect 11418 8058 11496 8064
rect 11418 7590 11424 8058
rect 11490 7590 11496 8058
rect 11418 7584 11496 7590
rect 11934 8058 12012 8064
rect 11934 7590 11940 8058
rect 12006 7590 12012 8058
rect 11934 7584 12012 7590
rect 12332 8042 12398 8054
rect 6518 7406 6596 7412
rect 6518 7072 6524 7406
rect 6590 7072 6596 7406
rect 6518 7066 6596 7072
rect 7034 7406 7112 7412
rect 7034 7072 7040 7406
rect 7106 7072 7112 7406
rect 7034 7066 7112 7072
rect 7550 7406 7628 7412
rect 7550 7072 7556 7406
rect 7622 7072 7628 7406
rect 7550 7066 7628 7072
rect 8066 7406 8144 7412
rect 8066 7072 8072 7406
rect 8138 7072 8144 7406
rect 8066 7066 8144 7072
rect 8582 7406 8660 7412
rect 8582 7072 8588 7406
rect 8654 7072 8660 7406
rect 8582 7066 8660 7072
rect 9098 7406 9176 7412
rect 9098 7072 9104 7406
rect 9170 7072 9176 7406
rect 9098 7066 9176 7072
rect 9614 7406 9692 7412
rect 9614 7072 9620 7406
rect 9686 7072 9692 7406
rect 9614 7066 9692 7072
rect 10130 7406 10208 7412
rect 10130 7072 10136 7406
rect 10202 7072 10208 7406
rect 10130 7066 10208 7072
rect 10646 7406 10724 7412
rect 10646 7072 10652 7406
rect 10718 7072 10724 7406
rect 10646 7066 10724 7072
rect 11162 7406 11240 7412
rect 11162 7072 11168 7406
rect 11234 7072 11240 7406
rect 11162 7066 11240 7072
rect 11678 7406 11756 7412
rect 11678 7072 11684 7406
rect 11750 7072 11756 7406
rect 11678 7066 11756 7072
rect 12194 7406 12272 7412
rect 12194 7072 12200 7406
rect 12266 7072 12272 7406
rect 12194 7066 12272 7072
rect 12332 7074 12348 8042
rect 12384 7074 12398 8042
rect 12332 7058 12398 7074
rect 12482 7030 12548 8094
rect 14424 7988 14916 8218
rect 6330 6984 12548 7030
rect 6518 6942 6596 6948
rect 6518 6608 6524 6942
rect 6590 6608 6596 6942
rect 6518 6602 6596 6608
rect 7034 6942 7112 6948
rect 7034 6608 7040 6942
rect 7106 6608 7112 6942
rect 7034 6602 7112 6608
rect 7550 6942 7628 6948
rect 7550 6608 7556 6942
rect 7622 6608 7628 6942
rect 7550 6602 7628 6608
rect 8066 6942 8144 6948
rect 8066 6608 8072 6942
rect 8138 6608 8144 6942
rect 8066 6602 8144 6608
rect 8582 6942 8660 6948
rect 8582 6608 8588 6942
rect 8654 6608 8660 6942
rect 8582 6602 8660 6608
rect 9098 6942 9176 6948
rect 9098 6608 9104 6942
rect 9170 6608 9176 6942
rect 9098 6602 9176 6608
rect 9614 6942 9692 6948
rect 9614 6608 9620 6942
rect 9686 6608 9692 6942
rect 9614 6602 9692 6608
rect 10130 6942 10208 6948
rect 10130 6608 10136 6942
rect 10202 6608 10208 6942
rect 10130 6602 10208 6608
rect 10646 6942 10724 6948
rect 10646 6608 10652 6942
rect 10718 6608 10724 6942
rect 10646 6602 10724 6608
rect 11162 6942 11240 6948
rect 11162 6608 11168 6942
rect 11234 6608 11240 6942
rect 11162 6602 11240 6608
rect 11678 6942 11756 6948
rect 11678 6608 11684 6942
rect 11750 6608 11756 6942
rect 11678 6602 11756 6608
rect 12194 6942 12272 6948
rect 12194 6608 12200 6942
rect 12266 6608 12272 6942
rect 12194 6602 12272 6608
rect 12330 6932 12396 6946
rect 6260 6326 6338 6332
rect 6260 5960 6266 6326
rect 6332 5960 6338 6326
rect 6260 5954 6338 5960
rect 6776 6326 6854 6332
rect 6776 5960 6782 6326
rect 6848 5960 6854 6326
rect 6776 5954 6854 5960
rect 7292 6326 7370 6332
rect 7292 5960 7298 6326
rect 7364 5960 7370 6326
rect 7292 5954 7370 5960
rect 7808 6326 7886 6332
rect 7808 5960 7814 6326
rect 7880 5960 7886 6326
rect 7808 5954 7886 5960
rect 8324 6326 8402 6332
rect 8324 5960 8330 6326
rect 8396 5960 8402 6326
rect 8324 5954 8402 5960
rect 8840 6326 8918 6332
rect 8840 5960 8846 6326
rect 8912 5960 8918 6326
rect 8840 5954 8918 5960
rect 9356 6326 9434 6332
rect 9356 5960 9362 6326
rect 9428 5960 9434 6326
rect 9356 5954 9434 5960
rect 9872 6326 9950 6332
rect 9872 5960 9878 6326
rect 9944 5960 9950 6326
rect 9872 5954 9950 5960
rect 10388 6326 10466 6332
rect 10388 5960 10394 6326
rect 10460 5960 10466 6326
rect 10388 5954 10466 5960
rect 10904 6326 10982 6332
rect 10904 5960 10910 6326
rect 10976 5960 10982 6326
rect 10904 5954 10982 5960
rect 11420 6326 11498 6332
rect 11420 5960 11426 6326
rect 11492 5960 11498 6326
rect 11420 5954 11498 5960
rect 11936 6326 12014 6332
rect 11936 5960 11942 6326
rect 12008 5960 12014 6326
rect 11936 5954 12014 5960
rect 12330 5964 12348 6932
rect 12384 5964 12396 6932
rect 12330 5950 12396 5964
rect 12482 5920 12548 6984
rect 6330 5874 12548 5920
rect 12334 5824 12400 5832
rect 6260 5818 6338 5824
rect 6260 5452 6266 5818
rect 6332 5452 6338 5818
rect 6260 5446 6338 5452
rect 6776 5818 6854 5824
rect 6776 5452 6782 5818
rect 6848 5452 6854 5818
rect 6776 5446 6854 5452
rect 7292 5818 7370 5824
rect 7292 5452 7298 5818
rect 7364 5452 7370 5818
rect 7292 5446 7370 5452
rect 7808 5818 7886 5824
rect 7808 5452 7814 5818
rect 7880 5452 7886 5818
rect 7808 5446 7886 5452
rect 8324 5818 8402 5824
rect 8324 5452 8330 5818
rect 8396 5452 8402 5818
rect 8324 5446 8402 5452
rect 8840 5818 8918 5824
rect 8840 5452 8846 5818
rect 8912 5452 8918 5818
rect 8840 5446 8918 5452
rect 9356 5818 9434 5824
rect 9356 5452 9362 5818
rect 9428 5452 9434 5818
rect 9356 5446 9434 5452
rect 9872 5818 9950 5824
rect 9872 5452 9878 5818
rect 9944 5452 9950 5818
rect 9872 5446 9950 5452
rect 10388 5818 10466 5824
rect 10388 5452 10394 5818
rect 10460 5452 10466 5818
rect 10388 5446 10466 5452
rect 10904 5818 10982 5824
rect 10904 5452 10910 5818
rect 10976 5452 10982 5818
rect 10904 5446 10982 5452
rect 11420 5818 11498 5824
rect 11420 5452 11426 5818
rect 11492 5452 11498 5818
rect 11420 5446 11498 5452
rect 11936 5818 12014 5824
rect 11936 5452 11942 5818
rect 12008 5452 12014 5818
rect 11936 5446 12014 5452
rect 6518 5186 6596 5192
rect 6518 4852 6524 5186
rect 6590 4852 6596 5186
rect 6518 4846 6596 4852
rect 7034 5186 7112 5192
rect 7034 4852 7040 5186
rect 7106 4852 7112 5186
rect 7034 4846 7112 4852
rect 7550 5186 7628 5192
rect 7550 4852 7556 5186
rect 7622 4852 7628 5186
rect 7550 4846 7628 4852
rect 8066 5186 8144 5192
rect 8066 4852 8072 5186
rect 8138 4852 8144 5186
rect 8066 4846 8144 4852
rect 8582 5186 8660 5192
rect 8582 4852 8588 5186
rect 8654 4852 8660 5186
rect 8582 4846 8660 4852
rect 9098 5186 9176 5192
rect 9098 4852 9104 5186
rect 9170 4852 9176 5186
rect 9098 4846 9176 4852
rect 9614 5186 9692 5192
rect 9614 4852 9620 5186
rect 9686 4852 9692 5186
rect 9614 4846 9692 4852
rect 10130 5186 10208 5192
rect 10130 4852 10136 5186
rect 10202 4852 10208 5186
rect 10130 4846 10208 4852
rect 10646 5186 10724 5192
rect 10646 4852 10652 5186
rect 10718 4852 10724 5186
rect 10646 4846 10724 4852
rect 11162 5186 11240 5192
rect 11162 4852 11168 5186
rect 11234 4852 11240 5186
rect 11162 4846 11240 4852
rect 11678 5186 11756 5192
rect 11678 4852 11684 5186
rect 11750 4852 11756 5186
rect 11678 4846 11756 4852
rect 12194 5186 12272 5192
rect 12194 4852 12200 5186
rect 12266 4852 12272 5186
rect 12194 4846 12272 4852
rect 12334 4856 12348 5824
rect 12384 4856 12400 5824
rect 12334 4842 12400 4856
rect 12482 4810 12548 5874
rect 6334 4764 12548 4810
rect 6518 4722 6596 4728
rect 6518 4388 6524 4722
rect 6590 4388 6596 4722
rect 6518 4382 6596 4388
rect 7034 4722 7112 4728
rect 7034 4388 7040 4722
rect 7106 4388 7112 4722
rect 7034 4382 7112 4388
rect 7550 4722 7628 4728
rect 7550 4388 7556 4722
rect 7622 4388 7628 4722
rect 7550 4382 7628 4388
rect 8066 4722 8144 4728
rect 8066 4388 8072 4722
rect 8138 4388 8144 4722
rect 8066 4382 8144 4388
rect 8582 4722 8660 4728
rect 8582 4388 8588 4722
rect 8654 4388 8660 4722
rect 8582 4382 8660 4388
rect 9098 4722 9176 4728
rect 9098 4388 9104 4722
rect 9170 4388 9176 4722
rect 9098 4382 9176 4388
rect 9614 4722 9692 4728
rect 9614 4388 9620 4722
rect 9686 4388 9692 4722
rect 9614 4382 9692 4388
rect 10130 4722 10208 4728
rect 10130 4388 10136 4722
rect 10202 4388 10208 4722
rect 10130 4382 10208 4388
rect 10646 4722 10724 4728
rect 10646 4388 10652 4722
rect 10718 4388 10724 4722
rect 10646 4382 10724 4388
rect 11162 4722 11240 4728
rect 11162 4388 11168 4722
rect 11234 4388 11240 4722
rect 11162 4382 11240 4388
rect 11678 4722 11756 4728
rect 11678 4388 11684 4722
rect 11750 4388 11756 4722
rect 11678 4382 11756 4388
rect 12194 4722 12272 4728
rect 12194 4388 12200 4722
rect 12266 4388 12272 4722
rect 12194 4382 12272 4388
rect 12334 4716 12400 4726
rect 6260 4122 6338 4128
rect 6260 3756 6266 4122
rect 6332 3756 6338 4122
rect 6260 3750 6338 3756
rect 6776 4122 6854 4128
rect 6776 3756 6782 4122
rect 6848 3756 6854 4122
rect 6776 3750 6854 3756
rect 7292 4122 7370 4128
rect 7292 3756 7298 4122
rect 7364 3756 7370 4122
rect 7292 3750 7370 3756
rect 7808 4122 7886 4128
rect 7808 3756 7814 4122
rect 7880 3756 7886 4122
rect 7808 3750 7886 3756
rect 8324 4122 8402 4128
rect 8324 3756 8330 4122
rect 8396 3756 8402 4122
rect 8324 3750 8402 3756
rect 8840 4122 8918 4128
rect 8840 3756 8846 4122
rect 8912 3756 8918 4122
rect 8840 3750 8918 3756
rect 9356 4122 9434 4128
rect 9356 3756 9362 4122
rect 9428 3756 9434 4122
rect 9356 3750 9434 3756
rect 9872 4122 9950 4128
rect 9872 3756 9878 4122
rect 9944 3756 9950 4122
rect 9872 3750 9950 3756
rect 10388 4122 10466 4128
rect 10388 3756 10394 4122
rect 10460 3756 10466 4122
rect 10388 3750 10466 3756
rect 10904 4122 10982 4128
rect 10904 3756 10910 4122
rect 10976 3756 10982 4122
rect 10904 3750 10982 3756
rect 11420 4122 11498 4128
rect 11420 3756 11426 4122
rect 11492 3756 11498 4122
rect 11420 3750 11498 3756
rect 11936 4122 12014 4128
rect 11936 3756 11942 4122
rect 12008 3756 12014 4122
rect 11936 3750 12014 3756
rect 12334 3748 12348 4716
rect 12384 3748 12400 4716
rect 12334 3730 12400 3748
rect 12482 3700 12548 4764
rect 6316 3654 12548 3700
rect 6260 3614 6338 3620
rect 6260 3248 6266 3614
rect 6332 3248 6338 3614
rect 6260 3242 6338 3248
rect 6776 3614 6854 3620
rect 6776 3248 6782 3614
rect 6848 3248 6854 3614
rect 6776 3242 6854 3248
rect 7292 3614 7370 3620
rect 7292 3248 7298 3614
rect 7364 3248 7370 3614
rect 7292 3242 7370 3248
rect 7808 3614 7886 3620
rect 7808 3248 7814 3614
rect 7880 3248 7886 3614
rect 7808 3242 7886 3248
rect 8324 3614 8402 3620
rect 8324 3248 8330 3614
rect 8396 3248 8402 3614
rect 8324 3242 8402 3248
rect 8840 3614 8918 3620
rect 8840 3248 8846 3614
rect 8912 3248 8918 3614
rect 8840 3242 8918 3248
rect 9356 3614 9434 3620
rect 9356 3248 9362 3614
rect 9428 3248 9434 3614
rect 9356 3242 9434 3248
rect 9872 3614 9950 3620
rect 9872 3248 9878 3614
rect 9944 3248 9950 3614
rect 9872 3242 9950 3248
rect 10388 3614 10466 3620
rect 10388 3248 10394 3614
rect 10460 3248 10466 3614
rect 10388 3242 10466 3248
rect 10904 3614 10982 3620
rect 10904 3248 10910 3614
rect 10976 3248 10982 3614
rect 10904 3242 10982 3248
rect 11420 3614 11498 3620
rect 11420 3248 11426 3614
rect 11492 3248 11498 3614
rect 11420 3242 11498 3248
rect 11936 3614 12014 3620
rect 11936 3248 11942 3614
rect 12008 3248 12014 3614
rect 11936 3242 12014 3248
rect 12332 3602 12398 3614
rect 6518 2966 6596 2972
rect 6518 2632 6524 2966
rect 6590 2632 6596 2966
rect 6518 2626 6596 2632
rect 7034 2966 7112 2972
rect 7034 2632 7040 2966
rect 7106 2632 7112 2966
rect 7034 2626 7112 2632
rect 7550 2966 7628 2972
rect 7550 2632 7556 2966
rect 7622 2632 7628 2966
rect 7550 2626 7628 2632
rect 8066 2966 8144 2972
rect 8066 2632 8072 2966
rect 8138 2632 8144 2966
rect 8066 2626 8144 2632
rect 8582 2966 8660 2972
rect 8582 2632 8588 2966
rect 8654 2632 8660 2966
rect 8582 2626 8660 2632
rect 9098 2966 9176 2972
rect 9098 2632 9104 2966
rect 9170 2632 9176 2966
rect 9098 2626 9176 2632
rect 9614 2966 9692 2972
rect 9614 2632 9620 2966
rect 9686 2632 9692 2966
rect 9614 2626 9692 2632
rect 10130 2966 10208 2972
rect 10130 2632 10136 2966
rect 10202 2632 10208 2966
rect 10130 2626 10208 2632
rect 10646 2966 10724 2972
rect 10646 2632 10652 2966
rect 10718 2632 10724 2966
rect 10646 2626 10724 2632
rect 11162 2966 11240 2972
rect 11162 2632 11168 2966
rect 11234 2632 11240 2966
rect 11162 2626 11240 2632
rect 11678 2966 11756 2972
rect 11678 2632 11684 2966
rect 11750 2632 11756 2966
rect 11678 2626 11756 2632
rect 12194 2966 12272 2972
rect 12194 2632 12200 2966
rect 12266 2632 12272 2966
rect 12194 2626 12272 2632
rect 12332 2634 12348 3602
rect 12384 2634 12398 3602
rect 12332 2618 12398 2634
rect 12482 2590 12548 3654
rect 6324 2544 12548 2590
rect 6132 2460 6196 2509
rect 6132 2444 12434 2460
rect 6132 2386 6184 2444
rect 12402 2386 12434 2444
rect 6132 2338 12434 2386
rect 11184 2304 12054 2308
rect 11184 2300 11828 2304
rect 1876 2266 11828 2300
rect 1876 2194 1918 2266
rect 11306 2194 11828 2266
rect 1876 2164 11828 2194
rect 12036 2164 12054 2304
rect 1876 2158 12054 2164
rect 1876 1826 2010 2158
rect 11184 2156 12054 2158
rect 10706 2044 11138 2060
rect 10706 1938 10723 2044
rect 11120 1938 11138 2044
rect 10706 1922 11138 1938
rect 11234 1826 11368 2156
rect 1876 1822 12020 1826
rect 1876 1788 11830 1822
rect 1876 1716 1922 1788
rect 11310 1716 11830 1788
rect 1876 1714 11830 1716
rect 11998 1714 12020 1822
rect 1876 1690 12020 1714
rect 1876 1684 11370 1690
rect 11234 1680 11368 1684
rect 4674 1498 7750 1554
rect 778 1422 866 1426
rect 3750 1422 3838 1424
rect 778 1396 3838 1422
rect 4290 1412 4356 1440
rect 778 1356 866 1396
rect 3746 1356 3838 1396
rect 778 1332 3838 1356
rect 4058 1356 4170 1404
rect 778 1294 866 1332
rect 778 -904 806 1294
rect 852 -904 866 1294
rect 1010 1234 3994 1280
rect 916 1128 994 1134
rect 916 472 922 1128
rect 988 472 994 1128
rect 916 466 994 472
rect 1138 -124 1254 1192
rect 1416 1132 1532 1192
rect 1406 1126 1548 1132
rect 1406 472 1412 1126
rect 1542 472 1548 1126
rect 1406 466 1548 472
rect 1128 -130 1270 -124
rect 1128 -784 1134 -130
rect 1264 -784 1270 -130
rect 1128 -790 1270 -784
rect 1138 -798 1254 -790
rect 1416 -798 1532 466
rect 1694 -124 1810 1192
rect 1972 1132 2088 1192
rect 1962 1126 2104 1132
rect 1962 472 1968 1126
rect 2098 472 2104 1126
rect 1962 466 2104 472
rect 1684 -130 1826 -124
rect 1684 -784 1690 -130
rect 1820 -784 1826 -130
rect 1684 -790 1826 -784
rect 1694 -798 1810 -790
rect 1972 -798 2088 466
rect 2250 -124 2366 1192
rect 2528 1132 2644 1192
rect 2518 1126 2660 1132
rect 2518 472 2524 1126
rect 2654 472 2660 1126
rect 2518 466 2660 472
rect 2240 -130 2382 -124
rect 2240 -784 2246 -130
rect 2376 -784 2382 -130
rect 2240 -790 2382 -784
rect 2250 -798 2366 -790
rect 2528 -798 2644 466
rect 2806 -124 2922 1192
rect 3084 1132 3200 1192
rect 3362 1132 3478 1192
rect 3750 1182 3838 1202
rect 3618 1134 3696 1140
rect 3074 1126 3216 1132
rect 3074 472 3080 1126
rect 3210 472 3216 1126
rect 3618 478 3624 1134
rect 3690 478 3696 1134
rect 3618 472 3696 478
rect 3074 466 3216 472
rect 2796 -130 2938 -124
rect 2796 -784 2802 -130
rect 2932 -784 2938 -130
rect 2796 -790 2938 -784
rect 2806 -798 2922 -790
rect 3084 -798 3200 466
rect 3362 -124 3478 466
rect 3352 -130 3494 -124
rect 3352 -784 3358 -130
rect 3488 -784 3494 -130
rect 3352 -790 3494 -784
rect 3750 -790 3768 1182
rect 3814 -790 3838 1182
rect 3919 358 3994 1234
rect 3894 348 3994 358
rect 3894 -18 3904 348
rect 3982 -18 3994 348
rect 3894 -30 3994 -18
rect 3362 -798 3478 -790
rect 3750 -810 3838 -790
rect 3919 -848 3994 -30
rect 1010 -894 3994 -848
rect 4058 -786 4074 1356
rect 4152 -786 4170 1356
rect 4290 770 4300 1412
rect 4340 770 4356 1412
rect 4290 734 4356 770
rect 4402 734 4492 1340
rect 4276 728 4360 734
rect 4276 526 4282 728
rect 4356 526 4360 728
rect 4276 520 4360 526
rect 778 -940 866 -904
rect 778 -974 3838 -940
rect 778 -1014 866 -974
rect 3746 -1014 3838 -974
rect 778 -1028 3838 -1014
rect 832 -1030 3838 -1028
rect 4058 -998 4170 -786
rect 4290 482 4356 520
rect 4290 -856 4302 482
rect 4342 -812 4356 482
rect 4402 -766 4492 520
rect 4674 -780 4726 1498
rect 4902 1034 5068 1340
rect 4902 -766 5068 820
rect 5250 -780 5302 1498
rect 5478 734 5644 1340
rect 5478 -766 5644 520
rect 5826 -780 5878 1498
rect 6054 1034 6220 1340
rect 6054 -766 6220 820
rect 6402 -780 6454 1498
rect 6630 734 6796 1340
rect 6630 -766 6796 520
rect 6978 -780 7030 1498
rect 7352 1412 7418 1440
rect 7206 1034 7296 1340
rect 7206 -766 7296 820
rect 7352 770 7364 1412
rect 7404 770 7418 1412
rect 7352 734 7418 770
rect 7528 1394 7638 1422
rect 7336 726 7430 734
rect 7336 530 7344 726
rect 7424 530 7430 726
rect 7336 528 7348 530
rect 7388 528 7430 530
rect 7336 520 7430 528
rect 7352 482 7418 520
rect 7352 -812 7364 482
rect 4342 -830 7364 -812
rect 4342 -856 4410 -830
rect 4292 -872 4410 -856
rect 7290 -856 7364 -830
rect 7404 -856 7418 482
rect 7290 -872 7418 -856
rect 4292 -884 7418 -872
rect 7528 -808 7542 1394
rect 7620 -808 7638 1394
rect 7528 -998 7638 -808
rect 4058 -1016 7638 -998
rect 4058 -1068 4102 -1016
rect 7506 -1068 7638 -1016
rect 4058 -1084 7638 -1068
rect 7694 1226 7750 1498
rect 8402 1490 11490 1546
rect 7798 1404 8358 1432
rect 7798 1334 7834 1404
rect 8322 1334 8358 1404
rect 7798 1282 8358 1334
rect 8402 1226 8458 1490
rect 7694 1180 8006 1226
rect 8142 1220 8458 1226
rect 8142 1186 8156 1220
rect 8210 1186 8458 1220
rect 8142 1180 8458 1186
rect 7694 -384 7750 1180
rect 8072 1032 8160 1046
rect 8072 820 8080 1032
rect 8150 820 8160 1032
rect 8072 810 8160 820
rect 7862 734 7950 744
rect 7862 522 7872 734
rect 7942 522 7950 734
rect 7862 508 7950 522
rect 7998 434 8082 442
rect 7778 428 7848 434
rect 7778 228 7786 428
rect 7838 228 7848 428
rect 7778 220 7848 228
rect 7998 222 8004 434
rect 8078 222 8082 434
rect 7998 212 8082 222
rect 8208 434 8374 442
rect 8208 222 8214 434
rect 8288 222 8328 434
rect 8362 222 8374 434
rect 8208 212 8374 222
rect 8402 -384 8458 1180
rect 7694 -390 8014 -384
rect 7694 -424 7944 -390
rect 8002 -424 8014 -390
rect 7694 -430 8014 -424
rect 8150 -430 8458 -384
rect 7694 -884 7750 -430
rect 7796 -540 8356 -488
rect 7796 -610 7830 -540
rect 8318 -610 8356 -540
rect 7796 -638 8356 -610
rect 8402 -884 8458 -430
rect 7694 -1084 7894 -884
rect 8258 -1084 8458 -884
rect 8520 1398 8630 1428
rect 8520 -804 8534 1398
rect 8612 -804 8630 1398
rect 8756 1420 8822 1442
rect 8756 1086 8768 1420
rect 8812 1086 8822 1420
rect 8756 1034 8822 1086
rect 8870 1034 8958 1362
rect 8738 1030 8832 1034
rect 8738 828 8746 1030
rect 8822 828 8832 1030
rect 8738 820 8832 828
rect 8520 -1002 8630 -804
rect 8756 778 8822 820
rect 8756 -812 8768 778
rect 8810 -812 8822 778
rect 8870 -744 8958 820
rect 9134 -764 9186 1490
rect 9368 734 9534 1362
rect 9368 -744 9534 520
rect 9710 -764 9762 1490
rect 9944 1034 10110 1362
rect 9944 -744 10110 820
rect 10286 -764 10338 1490
rect 10520 734 10686 1362
rect 10520 -744 10686 520
rect 10862 -764 10914 1490
rect 11096 1034 11262 1362
rect 11096 -744 11262 820
rect 11438 -764 11490 1490
rect 11810 1402 11876 1446
rect 11672 734 11758 1362
rect 11810 1068 11822 1402
rect 11866 1068 11876 1402
rect 11810 1034 11876 1068
rect 11968 1416 12078 1526
rect 11804 1028 11902 1034
rect 11804 830 11814 1028
rect 11894 830 11902 1028
rect 11804 820 11902 830
rect 11672 -744 11758 520
rect 11810 776 11876 820
rect 11810 -812 11822 776
rect 8756 -814 11822 -812
rect 11864 -814 11876 776
rect 8756 -828 11876 -814
rect 8756 -866 8872 -828
rect 11768 -866 11876 -828
rect 8756 -880 11876 -866
rect 11968 -826 11984 1416
rect 12062 -180 12078 1416
rect 12062 -198 12212 -180
rect 12062 -606 12106 -198
rect 12062 -628 12212 -606
rect 12062 -826 12078 -628
rect 11968 -1002 12078 -826
rect 8520 -1018 12078 -1002
rect 8520 -1070 8674 -1018
rect 12050 -1070 12078 -1018
rect 4058 -1086 4170 -1084
rect 8520 -1088 12078 -1070
rect 12482 -1079 12548 2544
rect 12590 7980 14981 7988
rect 12590 7946 12692 7980
rect 14878 7946 14981 7980
rect 12590 7938 14981 7946
rect 12590 7884 12636 7938
rect 14932 7884 14981 7938
rect 12590 -180 12596 7884
rect 12588 -526 12596 -180
rect 12630 -526 12636 7884
rect 12794 7838 13128 7884
rect 13586 7838 14904 7884
rect 12670 6338 12770 7792
rect 12670 5960 12680 6338
rect 12670 3758 12770 5960
rect 13734 4080 13834 7792
rect 13734 3798 13834 3808
rect 14792 5844 14892 7792
rect 14792 3788 14892 5482
rect 12670 3602 14822 3758
rect 12666 734 12766 3572
rect 12666 -440 12766 518
rect 13738 3564 13838 3574
rect 13738 -128 13838 3292
rect 13738 -438 13838 -428
rect 14782 1560 14882 3568
rect 14782 -444 14882 1364
rect 12796 -526 13110 -480
rect 13618 -526 14886 -480
rect 14932 -526 14940 7884
rect 14974 -526 14981 7884
rect 12588 -581 12636 -526
rect 14932 -581 14981 -526
rect 12588 -588 14981 -581
rect 12588 -622 12692 -588
rect 14878 -622 14981 -588
rect 12588 -628 14981 -622
rect 12590 -629 14981 -628
rect 12698 -656 14886 -629
rect 12698 -722 12722 -656
rect 14850 -722 14886 -656
rect 12698 -742 14886 -722
<< via1 >>
rect 6178 8240 12314 8278
rect 6178 8220 12314 8240
rect 6264 7590 6330 8058
rect 6780 7590 6846 8058
rect 7296 7590 7362 8058
rect 7812 7590 7878 8058
rect 8328 7590 8394 8058
rect 8844 7590 8910 8058
rect 9360 7590 9426 8058
rect 9876 7590 9942 8058
rect 10392 7590 10458 8058
rect 10908 7590 10974 8058
rect 11424 7590 11490 8058
rect 11940 7590 12006 8058
rect 6524 7072 6590 7406
rect 7040 7072 7106 7406
rect 7556 7072 7622 7406
rect 8072 7072 8138 7406
rect 8588 7072 8654 7406
rect 9104 7072 9170 7406
rect 9620 7072 9686 7406
rect 10136 7072 10202 7406
rect 10652 7072 10718 7406
rect 11168 7072 11234 7406
rect 11684 7072 11750 7406
rect 12200 7072 12266 7406
rect 6524 6608 6590 6942
rect 7040 6608 7106 6942
rect 7556 6608 7622 6942
rect 8072 6608 8138 6942
rect 8588 6608 8654 6942
rect 9104 6608 9170 6942
rect 9620 6608 9686 6942
rect 10136 6608 10202 6942
rect 10652 6608 10718 6942
rect 11168 6608 11234 6942
rect 11684 6608 11750 6942
rect 12200 6608 12266 6942
rect 6266 5960 6332 6326
rect 6782 5960 6848 6326
rect 7298 5960 7364 6326
rect 7814 5960 7880 6326
rect 8330 5960 8396 6326
rect 8846 5960 8912 6326
rect 9362 5960 9428 6326
rect 9878 5960 9944 6326
rect 10394 5960 10460 6326
rect 10910 5960 10976 6326
rect 11426 5960 11492 6326
rect 11942 5960 12008 6326
rect 6266 5452 6332 5818
rect 6782 5452 6848 5818
rect 7298 5452 7364 5818
rect 7814 5452 7880 5818
rect 8330 5452 8396 5818
rect 8846 5452 8912 5818
rect 9362 5452 9428 5818
rect 9878 5452 9944 5818
rect 10394 5452 10460 5818
rect 10910 5452 10976 5818
rect 11426 5452 11492 5818
rect 11942 5452 12008 5818
rect 6524 4852 6590 5186
rect 7040 4852 7106 5186
rect 7556 4852 7622 5186
rect 8072 4852 8138 5186
rect 8588 4852 8654 5186
rect 9104 4852 9170 5186
rect 9620 4852 9686 5186
rect 10136 4852 10202 5186
rect 10652 4852 10718 5186
rect 11168 4852 11234 5186
rect 11684 4852 11750 5186
rect 12200 4852 12266 5186
rect 6524 4388 6590 4722
rect 7040 4388 7106 4722
rect 7556 4388 7622 4722
rect 8072 4388 8138 4722
rect 8588 4388 8654 4722
rect 9104 4388 9170 4722
rect 9620 4388 9686 4722
rect 10136 4388 10202 4722
rect 10652 4388 10718 4722
rect 11168 4388 11234 4722
rect 11684 4388 11750 4722
rect 12200 4388 12266 4722
rect 6266 3756 6332 4122
rect 6782 3756 6848 4122
rect 7298 3756 7364 4122
rect 7814 3756 7880 4122
rect 8330 3756 8396 4122
rect 8846 3756 8912 4122
rect 9362 3756 9428 4122
rect 9878 3756 9944 4122
rect 10394 3756 10460 4122
rect 10910 3756 10976 4122
rect 11426 3756 11492 4122
rect 11942 3756 12008 4122
rect 6266 3248 6332 3614
rect 6782 3248 6848 3614
rect 7298 3248 7364 3614
rect 7814 3248 7880 3614
rect 8330 3248 8396 3614
rect 8846 3248 8912 3614
rect 9362 3248 9428 3614
rect 9878 3248 9944 3614
rect 10394 3248 10460 3614
rect 10910 3248 10976 3614
rect 11426 3248 11492 3614
rect 11942 3248 12008 3614
rect 6524 2632 6590 2966
rect 7040 2632 7106 2966
rect 7556 2632 7622 2966
rect 8072 2632 8138 2966
rect 8588 2632 8654 2966
rect 9104 2632 9170 2966
rect 9620 2632 9686 2966
rect 10136 2632 10202 2966
rect 10652 2632 10718 2966
rect 11168 2632 11234 2966
rect 11684 2632 11750 2966
rect 12200 2632 12266 2966
rect 11828 2164 12036 2304
rect 2126 1940 2516 2042
rect 10723 1938 11120 2044
rect 11830 1714 11998 1822
rect 922 472 988 1128
rect 1412 472 1542 1126
rect 1134 -784 1264 -130
rect 1968 472 2098 1126
rect 1690 -784 1820 -130
rect 2524 472 2654 1126
rect 2246 -784 2376 -130
rect 3080 472 3210 1126
rect 3624 478 3690 1134
rect 2802 -784 2932 -130
rect 3358 -784 3488 -130
rect 3904 -18 3982 348
rect 4282 724 4356 728
rect 4282 528 4308 724
rect 4308 528 4346 724
rect 4346 528 4356 724
rect 4282 526 4356 528
rect 4402 520 4492 734
rect 4902 820 5068 1034
rect 5478 520 5644 734
rect 6054 820 6220 1034
rect 6630 520 6796 734
rect 7206 820 7296 1034
rect 7344 530 7348 726
rect 7348 530 7388 726
rect 7388 530 7424 726
rect 4102 -1018 7506 -1016
rect 4102 -1068 7506 -1018
rect 8080 820 8150 1032
rect 7872 522 7942 734
rect 7786 228 7794 428
rect 7794 228 7830 428
rect 7830 228 7838 428
rect 8004 222 8078 434
rect 8214 222 8288 434
rect 8746 1028 8822 1030
rect 8746 828 8778 1028
rect 8778 828 8818 1028
rect 8818 828 8822 1028
rect 8870 820 8958 1034
rect 9368 520 9534 734
rect 9944 820 10110 1034
rect 10520 520 10686 734
rect 11096 820 11262 1034
rect 11814 830 11818 1028
rect 11818 830 11858 1028
rect 11858 830 11894 1028
rect 11672 520 11758 734
rect 12106 -606 12212 -198
rect 8674 -1020 12050 -1018
rect 8674 -1070 12050 -1020
rect 12680 5960 12770 6338
rect 13734 3808 13834 4080
rect 14792 5482 14892 5844
rect 12666 518 12766 734
rect 13738 3292 13838 3564
rect 13738 -428 13838 -128
rect 14782 1364 14882 1560
rect 12722 -722 14850 -656
<< metal2 >>
rect 6150 8280 14916 8282
rect 6150 8278 12702 8280
rect 6150 8220 6178 8278
rect 12314 8220 12702 8278
rect 6150 8058 12702 8220
rect 6150 7590 6264 8058
rect 6330 7590 6780 8058
rect 6846 7590 7296 8058
rect 7362 7590 7812 8058
rect 7878 7590 8328 8058
rect 8394 7590 8844 8058
rect 8910 7590 9360 8058
rect 9426 7590 9876 8058
rect 9942 7590 10392 8058
rect 10458 7590 10908 8058
rect 10974 7590 11424 8058
rect 11490 7590 11940 8058
rect 12006 7590 12702 8058
rect 6150 7584 12702 7590
rect 12944 7584 14916 8280
rect 6150 7582 14916 7584
rect 628 7406 11364 7414
rect 628 7398 6524 7406
rect 628 6536 644 7398
rect 824 7072 6524 7398
rect 6590 7072 7040 7406
rect 7106 7072 7556 7406
rect 7622 7072 8072 7406
rect 8138 7072 8588 7406
rect 8654 7072 9104 7406
rect 9170 7072 9620 7406
rect 9686 7072 10136 7406
rect 10202 7072 10652 7406
rect 10718 7072 11168 7406
rect 11234 7072 11364 7406
rect 824 6942 11364 7072
rect 824 6608 6524 6942
rect 6590 6608 7040 6942
rect 7106 6608 7556 6942
rect 7622 6608 8072 6942
rect 8138 6608 8588 6942
rect 8654 6608 9104 6942
rect 9170 6608 9620 6942
rect 9686 6608 10136 6942
rect 10202 6608 10652 6942
rect 10718 6608 11168 6942
rect 11234 6608 11364 6942
rect 824 6536 11364 6608
rect 628 6522 11364 6536
rect 11540 7406 14916 7414
rect 11540 7072 11684 7406
rect 11750 7072 12200 7406
rect 12266 7398 14916 7406
rect 12266 7072 13882 7398
rect 11540 6942 13882 7072
rect 11540 6608 11684 6942
rect 11750 6608 12200 6942
rect 12266 6608 13882 6942
rect 11540 6550 13882 6608
rect 14024 6550 14916 7398
rect 11540 6522 14916 6550
rect 6184 6326 12512 6336
rect 6184 5960 6266 6326
rect 6332 5960 6782 6326
rect 6848 5960 7298 6326
rect 7364 5960 7814 6326
rect 7880 5960 8330 6326
rect 8396 5960 8846 6326
rect 8912 5960 9362 6326
rect 9428 5960 9878 6326
rect 9944 5960 10394 6326
rect 10460 5960 10910 6326
rect 10976 5960 11426 6326
rect 11492 5960 11942 6326
rect 12008 5960 12512 6326
rect 12674 5960 12680 6338
rect 12770 5962 14132 6338
rect 14306 5962 14916 6338
rect 12770 5960 14916 5962
rect 6184 5894 12512 5960
rect 6184 5818 12698 5894
rect 6184 5452 6266 5818
rect 6332 5452 6782 5818
rect 6848 5452 7298 5818
rect 7364 5452 7814 5818
rect 7880 5452 8330 5818
rect 8396 5452 8846 5818
rect 8912 5452 9362 5818
rect 9428 5452 9878 5818
rect 9944 5452 10394 5818
rect 10460 5452 10910 5818
rect 10976 5452 11426 5818
rect 11492 5452 11942 5818
rect 12008 5452 12698 5818
rect 6184 5444 12698 5452
rect 12950 5444 12976 5894
rect 13064 5482 13084 5844
rect 13360 5482 14792 5844
rect 14892 5482 14916 5844
rect 628 5238 11382 5254
rect 628 4376 642 5238
rect 822 5186 11382 5238
rect 822 4852 6524 5186
rect 6590 4852 7040 5186
rect 7106 4852 7556 5186
rect 7622 4852 8072 5186
rect 8138 4852 8588 5186
rect 8654 4852 9104 5186
rect 9170 4852 9620 5186
rect 9686 4852 10136 5186
rect 10202 4852 10652 5186
rect 10718 4852 11168 5186
rect 11234 4852 11382 5186
rect 822 4722 11382 4852
rect 822 4388 6524 4722
rect 6590 4388 7040 4722
rect 7106 4388 7556 4722
rect 7622 4388 8072 4722
rect 8138 4388 8588 4722
rect 8654 4388 9104 4722
rect 9170 4388 9620 4722
rect 9686 4388 10136 4722
rect 10202 4388 10652 4722
rect 10718 4388 11168 4722
rect 11234 4388 11382 4722
rect 822 4376 11382 4388
rect 628 4362 11382 4376
rect 11558 5234 14916 5254
rect 11558 5186 13884 5234
rect 11558 4852 11684 5186
rect 11750 4852 12200 5186
rect 12266 4852 13884 5186
rect 11558 4722 13884 4852
rect 11558 4388 11684 4722
rect 11750 4388 12200 4722
rect 12266 4388 13884 4722
rect 11558 4386 13884 4388
rect 14026 4386 14916 5234
rect 11558 4362 14916 4386
rect 6178 4122 12698 4130
rect 6178 3756 6266 4122
rect 6332 3756 6782 4122
rect 6848 3756 7298 4122
rect 7364 3756 7814 4122
rect 7880 3756 8330 4122
rect 8396 3756 8846 4122
rect 8912 3756 9362 4122
rect 9428 3756 9878 4122
rect 9944 3756 10394 4122
rect 10460 3756 10910 4122
rect 10976 3756 11426 4122
rect 11492 3756 11942 4122
rect 12008 3756 12698 4122
rect 6178 3614 12698 3756
rect 6178 3248 6266 3614
rect 6332 3248 6782 3614
rect 6848 3248 7298 3614
rect 7364 3248 7814 3614
rect 7880 3248 8330 3614
rect 8396 3248 8846 3614
rect 8912 3248 9362 3614
rect 9428 3248 9878 3614
rect 9944 3248 10394 3614
rect 10460 3248 10910 3614
rect 10976 3248 11426 3614
rect 11492 3248 11942 3614
rect 12008 3248 12698 3614
rect 6178 3238 12698 3248
rect 12950 3238 12974 4130
rect 13684 4120 14916 4140
rect 13684 4080 14448 4120
rect 13684 3808 13734 4080
rect 13834 3808 14448 4080
rect 13684 3564 14448 3808
rect 13684 3292 13738 3564
rect 13838 3310 14448 3564
rect 14900 3310 14916 4120
rect 13838 3292 14916 3310
rect 13684 3284 14916 3292
rect 628 3046 11376 3060
rect 628 2384 642 3046
rect 822 2966 11376 3046
rect 822 2632 6524 2966
rect 6590 2632 7040 2966
rect 7106 2632 7556 2966
rect 7622 2632 8072 2966
rect 8138 2632 8588 2966
rect 8654 2632 9104 2966
rect 9170 2632 9620 2966
rect 9686 2632 10136 2966
rect 10202 2632 10652 2966
rect 10718 2632 11168 2966
rect 11234 2632 11376 2966
rect 822 2384 11376 2632
rect 628 2368 11376 2384
rect 11552 3044 14916 3060
rect 11552 2966 13884 3044
rect 11552 2632 11684 2966
rect 11750 2632 12200 2966
rect 12266 2632 13884 2966
rect 11552 2390 13884 2632
rect 14024 2390 14916 3044
rect 11552 2368 14916 2390
rect 11814 2304 12702 2306
rect 11814 2164 11828 2304
rect 12036 2164 12702 2304
rect 11814 2162 12702 2164
rect 12946 2162 12956 2306
rect 13472 2214 13772 2238
rect 13472 2106 13498 2214
rect 628 2094 2572 2104
rect 628 1902 638 2094
rect 828 2042 2572 2094
rect 828 1940 2126 2042
rect 2516 1940 2572 2042
rect 828 1902 2572 1940
rect 628 1890 2572 1902
rect 10668 2044 13498 2106
rect 10668 1938 10723 2044
rect 11120 1938 13498 2044
rect 10668 1908 13498 1938
rect 13750 2106 13772 2214
rect 13750 1908 13774 2106
rect 10668 1878 13774 1908
rect 11818 1714 11830 1822
rect 11998 1714 12702 1822
rect 12946 1714 12958 1822
rect 628 1448 3866 1460
rect 628 468 642 1448
rect 822 1134 3866 1448
rect 822 1128 3624 1134
rect 822 472 922 1128
rect 988 1126 3624 1128
rect 988 472 1412 1126
rect 1542 472 1968 1126
rect 2098 472 2524 1126
rect 2654 472 3080 1126
rect 3210 478 3624 1126
rect 3690 478 3866 1134
rect 7348 1364 14126 1560
rect 14316 1364 14782 1560
rect 14882 1364 14926 1560
rect 7348 1034 7544 1364
rect 4276 820 4902 1034
rect 5068 820 6054 1034
rect 6220 820 7206 1034
rect 7296 822 7544 1034
rect 7656 1032 8870 1034
rect 7296 820 7516 822
rect 7656 820 8080 1032
rect 8150 1030 8870 1032
rect 8150 828 8746 1030
rect 8822 828 8870 1030
rect 8150 820 8870 828
rect 8958 820 9944 1034
rect 10110 820 11096 1034
rect 11262 1028 11994 1034
rect 11262 830 11814 1028
rect 11894 830 11994 1028
rect 11262 820 11994 830
rect 4276 728 4402 734
rect 4276 526 4282 728
rect 4356 526 4402 728
rect 4276 520 4402 526
rect 4492 520 5478 734
rect 5644 520 6630 734
rect 6796 726 7872 734
rect 6796 530 7344 726
rect 7424 530 7872 726
rect 6796 522 7872 530
rect 7942 522 8488 734
rect 6796 520 8488 522
rect 8708 520 9368 734
rect 9534 520 10520 734
rect 10686 520 11672 734
rect 11758 520 12666 734
rect 12071 518 12666 520
rect 12766 518 13084 734
rect 13358 518 14926 734
rect 3210 472 3866 478
rect 822 468 3866 472
rect 628 454 3866 468
rect 4276 428 8004 434
rect 3878 348 3994 358
rect 3878 164 3904 348
rect 3982 176 3994 348
rect 4276 228 7786 428
rect 7838 228 8004 428
rect 4276 222 8004 228
rect 8078 222 8214 434
rect 8288 424 14054 434
rect 8288 230 13882 424
rect 14038 230 14054 424
rect 8288 222 14054 230
rect 4276 220 14054 222
rect 3982 164 4082 176
rect 3878 -26 3892 164
rect 4068 -26 4082 164
rect 3878 -38 4082 -26
rect 712 -128 14916 -114
rect 712 -130 13738 -128
rect 712 -784 1134 -130
rect 1264 -784 1690 -130
rect 1820 -784 2246 -130
rect 2376 -784 2802 -130
rect 2932 -784 3358 -130
rect 3488 -198 13738 -130
rect 3488 -606 12106 -198
rect 12212 -428 13738 -198
rect 13838 -132 14916 -128
rect 13838 -428 14438 -132
rect 12212 -606 14438 -428
rect 3488 -656 14438 -606
rect 3488 -722 12722 -656
rect 3488 -784 14438 -722
rect 712 -1016 14438 -784
rect 712 -1068 4102 -1016
rect 7506 -1018 14438 -1016
rect 7506 -1068 8674 -1018
rect 712 -1070 8674 -1068
rect 12050 -1064 14438 -1018
rect 14896 -1064 14916 -132
rect 12050 -1070 14916 -1064
rect 712 -1084 14916 -1070
rect 4052 -1094 7644 -1084
rect 8518 -1086 12096 -1084
rect 8518 -1090 12080 -1086
<< via2 >>
rect 12702 7584 12944 8280
rect 644 6536 824 7398
rect 13882 6550 14024 7398
rect 14132 5962 14306 6338
rect 12698 5444 12950 5894
rect 13084 5482 13360 5844
rect 642 4376 822 5238
rect 13884 4386 14026 5234
rect 12698 3238 12950 4130
rect 14448 3310 14900 4120
rect 642 2384 822 3046
rect 13884 2390 14024 3044
rect 12702 2162 12946 2306
rect 638 1902 828 2094
rect 13498 1908 13750 2214
rect 12702 1714 12946 1822
rect 642 468 822 1448
rect 14126 1364 14316 1560
rect 13084 518 13358 734
rect 13882 230 14038 424
rect 3892 -18 3904 164
rect 3904 -18 3982 164
rect 3982 -18 4068 164
rect 3892 -26 4068 -18
rect 14438 -656 14896 -132
rect 14438 -722 14850 -656
rect 14850 -722 14896 -656
rect 14438 -1064 14896 -722
<< metal3 >>
rect 12690 8280 12960 8290
rect 12690 7584 12702 8280
rect 12944 7584 12960 8280
rect 13474 8076 13774 8132
rect 13474 7852 13514 8076
rect 13734 7852 13774 8076
rect 628 7398 840 7456
rect 628 6536 644 7398
rect 824 6536 840 7398
rect 628 5238 840 6536
rect 628 4376 642 5238
rect 822 4376 840 5238
rect 628 3046 840 4376
rect 628 2384 642 3046
rect 822 2384 840 3046
rect 628 2094 840 2384
rect 628 1902 638 2094
rect 828 1902 840 2094
rect 628 1448 840 1902
rect 628 468 642 1448
rect 822 468 840 1448
rect 628 374 840 468
rect 12690 5894 12960 7584
rect 12690 5444 12698 5894
rect 12950 5444 12960 5894
rect 12690 4130 12960 5444
rect 12690 3238 12698 4130
rect 12950 3238 12960 4130
rect 12690 2306 12960 3238
rect 12690 2162 12702 2306
rect 12946 2162 12960 2306
rect 12690 1822 12960 2162
rect 12690 1714 12702 1822
rect 12946 1714 12960 1822
rect 4256 176 4586 178
rect 3878 164 4586 176
rect 3878 -26 3892 164
rect 4068 158 4586 164
rect 4068 -26 4284 158
rect 3878 -38 4284 -26
rect 4256 -94 4284 -38
rect 4562 -94 4586 158
rect 12690 124 12960 1714
rect 13074 6794 13374 7750
rect 13074 6570 13114 6794
rect 13334 6570 13374 6794
rect 13074 5844 13374 6570
rect 13074 5482 13084 5844
rect 13360 5482 13374 5844
rect 13074 4188 13374 5482
rect 13074 3964 13114 4188
rect 13334 3964 13374 4188
rect 13074 1572 13374 3964
rect 13074 1348 13114 1572
rect 13334 1348 13374 1572
rect 13074 734 13374 1348
rect 13074 518 13084 734
rect 13358 518 13374 734
rect 13074 340 13374 518
rect 13474 5464 13774 7852
rect 13474 5240 13514 5464
rect 13734 5240 13774 5464
rect 13474 2856 13774 5240
rect 13474 2632 13514 2856
rect 13734 2632 13774 2856
rect 13474 2214 13774 2632
rect 13474 1908 13498 2214
rect 13750 1908 13774 2214
rect 4256 -126 4586 -94
rect 13474 -636 13774 1908
rect 13870 7398 14050 7762
rect 13870 6550 13882 7398
rect 14024 6550 14050 7398
rect 13870 5234 14050 6550
rect 13870 4386 13884 5234
rect 14026 4386 14050 5234
rect 13870 3044 14050 4386
rect 13870 2390 13884 3044
rect 14024 2390 14050 3044
rect 13870 424 14050 2390
rect 13870 230 13882 424
rect 14038 230 14050 424
rect 13870 204 14050 230
rect 14120 6338 14322 8154
rect 14120 5962 14132 6338
rect 14306 5962 14322 6338
rect 14120 1560 14322 5962
rect 14120 1364 14126 1560
rect 14316 1364 14322 1560
rect 14120 -940 14322 1364
rect 14422 4120 14922 8284
rect 14422 3310 14448 4120
rect 14900 3310 14922 4120
rect 14422 -132 14922 3310
rect 14422 -1064 14438 -132
rect 14896 -1064 14922 -132
rect 14422 -1090 14922 -1064
<< via3 >>
rect 13514 7852 13734 8076
rect 4284 -94 4562 158
rect 13114 6570 13334 6794
rect 13114 3964 13334 4188
rect 13114 1348 13334 1572
rect 13514 5240 13734 5464
rect 13514 2632 13734 2856
<< metal4 >>
rect 13474 8076 13774 8116
rect 13474 8012 13514 8076
rect 12458 7908 13514 8012
rect 13474 7852 13514 7908
rect 13734 7852 13774 8076
rect 13474 7814 13774 7852
rect 13074 6794 13374 6834
rect 13074 6732 13114 6794
rect 12466 6628 13114 6732
rect 13074 6570 13114 6628
rect 13334 6570 13374 6794
rect 13074 6530 13374 6570
rect 13474 5464 13774 5504
rect 13474 5400 13514 5464
rect 12466 5296 13514 5400
rect 13474 5240 13514 5296
rect 13734 5240 13774 5464
rect 13474 5200 13774 5240
rect 13074 4188 13374 4228
rect 13074 4120 13114 4188
rect 12466 4016 13114 4120
rect 13074 3964 13114 4016
rect 13334 3964 13374 4188
rect 13074 3924 13374 3964
rect 13474 2856 13774 2896
rect 13474 2788 13514 2856
rect 12466 2684 13514 2788
rect 13474 2632 13514 2684
rect 13734 2632 13774 2856
rect 13474 2592 13774 2632
rect 13074 1572 13374 1612
rect 13074 1508 13114 1572
rect 12466 1404 13114 1508
rect 13074 1348 13114 1404
rect 13334 1348 13374 1572
rect 13074 1308 13374 1348
rect 4366 178 4468 512
rect 4256 158 4586 178
rect 4256 -94 4284 158
rect 4562 -94 4586 158
rect 4256 -126 4586 -94
use sky130_fd_pr__cap_mim_m3_1_BHK9HY  sky130_fd_pr__cap_mim_m3_1_BHK9HY_0 paramcells
timestamp 1748311075
transform 0 1 6770 1 0 4214
box -3798 -5800 3798 5800
use sky130_fd_pr__nfet_05v0_nvt_FEJX3A  sky130_fd_pr__nfet_05v0_nvt_FEJX3A_0 paramcells
timestamp 1748311075
transform -1 0 10317 0 1 293
box -1580 -1194 1580 1194
use sky130_fd_pr__nfet_g5v0d10v5_NZU856  sky130_fd_pr__nfet_g5v0d10v5_NZU856_0 paramcells
timestamp 1748311075
transform 1 0 9265 0 1 5343
box -3166 -2978 3166 2978
use sky130_fd_pr__nfet_01v8_lvt_AJ3MPE  XM2 paramcells
timestamp 1748311075
transform -1 0 8078 0 1 398
box -320 -960 320 960
use sky130_fd_pr__pfet_01v8_lvt_UX3DP3  XM6 paramcells
timestamp 1748311075
transform 1 0 13785 0 1 3679
box -1225 -4337 1225 4337
use sky130_fd_pr__pfet_g5v0d10v5_8UL4MK  XM8 paramcells
timestamp 1748311075
transform 1 0 2311 0 1 193
box -1559 -1297 1559 1297
use sky130_fd_pr__nfet_05v0_nvt_FEJX3A  XM10
timestamp 1748311075
transform 1 0 5849 0 1 293
box -1580 -1194 1580 1194
use sky130_fd_pr__res_high_po_0p69_FJD3D2  XR1 paramcells
timestamp 1748311075
transform 0 1 6622 -1 0 1991
box -235 -4682 235 4682
<< labels >>
flabel metal2 13062 -1020 13262 -820 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal2 13052 8032 13252 8232 0 FreeSans 256 0 0 0 VSS
port 5 nsew
flabel metal1 12482 8108 12682 8308 0 FreeSans 256 0 0 0 VBIAS
port 4 nsew
flabel metal3 628 1502 840 1702 0 FreeSans 256 0 0 0 VOUT
port 1 nsew
flabel metal1 7694 -1084 7894 -884 0 FreeSans 256 0 0 0 VINN
port 2 nsew
flabel metal1 8258 -1084 8458 -884 0 FreeSans 256 0 0 0 VINP
port 3 nsew
<< end >>
