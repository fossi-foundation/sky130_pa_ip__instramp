magic
tech sky130A
magscale 1 2
timestamp 1729620069
<< pwell >>
rect -30070 -3082 30070 3082
<< psubdiff >>
rect -30034 3012 -29938 3046
rect 29938 3012 30034 3046
rect -30034 2950 -30000 3012
rect 30000 2950 30034 3012
rect -30034 -3012 -30000 -2950
rect 30000 -3012 30034 -2950
rect -30034 -3046 -29938 -3012
rect 29938 -3046 30034 -3012
<< psubdiffcont >>
rect -29938 3012 29938 3046
rect -30034 -2950 -30000 2950
rect 30000 -2950 30034 2950
rect -29938 -3046 29938 -3012
<< xpolycontact >>
rect -29904 2484 -29766 2916
rect -29904 -2916 -29766 -2484
rect -29670 2484 -29532 2916
rect -29670 -2916 -29532 -2484
rect -29436 2484 -29298 2916
rect -29436 -2916 -29298 -2484
rect -29202 2484 -29064 2916
rect -29202 -2916 -29064 -2484
rect -28968 2484 -28830 2916
rect -28968 -2916 -28830 -2484
rect -28734 2484 -28596 2916
rect -28734 -2916 -28596 -2484
rect -28500 2484 -28362 2916
rect -28500 -2916 -28362 -2484
rect -28266 2484 -28128 2916
rect -28266 -2916 -28128 -2484
rect -28032 2484 -27894 2916
rect -28032 -2916 -27894 -2484
rect -27798 2484 -27660 2916
rect -27798 -2916 -27660 -2484
rect -27564 2484 -27426 2916
rect -27564 -2916 -27426 -2484
rect -27330 2484 -27192 2916
rect -27330 -2916 -27192 -2484
rect -27096 2484 -26958 2916
rect -27096 -2916 -26958 -2484
rect -26862 2484 -26724 2916
rect -26862 -2916 -26724 -2484
rect -26628 2484 -26490 2916
rect -26628 -2916 -26490 -2484
rect -26394 2484 -26256 2916
rect -26394 -2916 -26256 -2484
rect -26160 2484 -26022 2916
rect -26160 -2916 -26022 -2484
rect -25926 2484 -25788 2916
rect -25926 -2916 -25788 -2484
rect -25692 2484 -25554 2916
rect -25692 -2916 -25554 -2484
rect -25458 2484 -25320 2916
rect -25458 -2916 -25320 -2484
rect -25224 2484 -25086 2916
rect -25224 -2916 -25086 -2484
rect -24990 2484 -24852 2916
rect -24990 -2916 -24852 -2484
rect -24756 2484 -24618 2916
rect -24756 -2916 -24618 -2484
rect -24522 2484 -24384 2916
rect -24522 -2916 -24384 -2484
rect -24288 2484 -24150 2916
rect -24288 -2916 -24150 -2484
rect -24054 2484 -23916 2916
rect -24054 -2916 -23916 -2484
rect -23820 2484 -23682 2916
rect -23820 -2916 -23682 -2484
rect -23586 2484 -23448 2916
rect -23586 -2916 -23448 -2484
rect -23352 2484 -23214 2916
rect -23352 -2916 -23214 -2484
rect -23118 2484 -22980 2916
rect -23118 -2916 -22980 -2484
rect -22884 2484 -22746 2916
rect -22884 -2916 -22746 -2484
rect -22650 2484 -22512 2916
rect -22650 -2916 -22512 -2484
rect -22416 2484 -22278 2916
rect -22416 -2916 -22278 -2484
rect -22182 2484 -22044 2916
rect -22182 -2916 -22044 -2484
rect -21948 2484 -21810 2916
rect -21948 -2916 -21810 -2484
rect -21714 2484 -21576 2916
rect -21714 -2916 -21576 -2484
rect -21480 2484 -21342 2916
rect -21480 -2916 -21342 -2484
rect -21246 2484 -21108 2916
rect -21246 -2916 -21108 -2484
rect -21012 2484 -20874 2916
rect -21012 -2916 -20874 -2484
rect -20778 2484 -20640 2916
rect -20778 -2916 -20640 -2484
rect -20544 2484 -20406 2916
rect -20544 -2916 -20406 -2484
rect -20310 2484 -20172 2916
rect -20310 -2916 -20172 -2484
rect -20076 2484 -19938 2916
rect -20076 -2916 -19938 -2484
rect -19842 2484 -19704 2916
rect -19842 -2916 -19704 -2484
rect -19608 2484 -19470 2916
rect -19608 -2916 -19470 -2484
rect -19374 2484 -19236 2916
rect -19374 -2916 -19236 -2484
rect -19140 2484 -19002 2916
rect -19140 -2916 -19002 -2484
rect -18906 2484 -18768 2916
rect -18906 -2916 -18768 -2484
rect -18672 2484 -18534 2916
rect -18672 -2916 -18534 -2484
rect -18438 2484 -18300 2916
rect -18438 -2916 -18300 -2484
rect -18204 2484 -18066 2916
rect -18204 -2916 -18066 -2484
rect -17970 2484 -17832 2916
rect -17970 -2916 -17832 -2484
rect -17736 2484 -17598 2916
rect -17736 -2916 -17598 -2484
rect -17502 2484 -17364 2916
rect -17502 -2916 -17364 -2484
rect -17268 2484 -17130 2916
rect -17268 -2916 -17130 -2484
rect -17034 2484 -16896 2916
rect -17034 -2916 -16896 -2484
rect -16800 2484 -16662 2916
rect -16800 -2916 -16662 -2484
rect -16566 2484 -16428 2916
rect -16566 -2916 -16428 -2484
rect -16332 2484 -16194 2916
rect -16332 -2916 -16194 -2484
rect -16098 2484 -15960 2916
rect -16098 -2916 -15960 -2484
rect -15864 2484 -15726 2916
rect -15864 -2916 -15726 -2484
rect -15630 2484 -15492 2916
rect -15630 -2916 -15492 -2484
rect -15396 2484 -15258 2916
rect -15396 -2916 -15258 -2484
rect -15162 2484 -15024 2916
rect -15162 -2916 -15024 -2484
rect -14928 2484 -14790 2916
rect -14928 -2916 -14790 -2484
rect -14694 2484 -14556 2916
rect -14694 -2916 -14556 -2484
rect -14460 2484 -14322 2916
rect -14460 -2916 -14322 -2484
rect -14226 2484 -14088 2916
rect -14226 -2916 -14088 -2484
rect -13992 2484 -13854 2916
rect -13992 -2916 -13854 -2484
rect -13758 2484 -13620 2916
rect -13758 -2916 -13620 -2484
rect -13524 2484 -13386 2916
rect -13524 -2916 -13386 -2484
rect -13290 2484 -13152 2916
rect -13290 -2916 -13152 -2484
rect -13056 2484 -12918 2916
rect -13056 -2916 -12918 -2484
rect -12822 2484 -12684 2916
rect -12822 -2916 -12684 -2484
rect -12588 2484 -12450 2916
rect -12588 -2916 -12450 -2484
rect -12354 2484 -12216 2916
rect -12354 -2916 -12216 -2484
rect -12120 2484 -11982 2916
rect -12120 -2916 -11982 -2484
rect -11886 2484 -11748 2916
rect -11886 -2916 -11748 -2484
rect -11652 2484 -11514 2916
rect -11652 -2916 -11514 -2484
rect -11418 2484 -11280 2916
rect -11418 -2916 -11280 -2484
rect -11184 2484 -11046 2916
rect -11184 -2916 -11046 -2484
rect -10950 2484 -10812 2916
rect -10950 -2916 -10812 -2484
rect -10716 2484 -10578 2916
rect -10716 -2916 -10578 -2484
rect -10482 2484 -10344 2916
rect -10482 -2916 -10344 -2484
rect -10248 2484 -10110 2916
rect -10248 -2916 -10110 -2484
rect -10014 2484 -9876 2916
rect -10014 -2916 -9876 -2484
rect -9780 2484 -9642 2916
rect -9780 -2916 -9642 -2484
rect -9546 2484 -9408 2916
rect -9546 -2916 -9408 -2484
rect -9312 2484 -9174 2916
rect -9312 -2916 -9174 -2484
rect -9078 2484 -8940 2916
rect -9078 -2916 -8940 -2484
rect -8844 2484 -8706 2916
rect -8844 -2916 -8706 -2484
rect -8610 2484 -8472 2916
rect -8610 -2916 -8472 -2484
rect -8376 2484 -8238 2916
rect -8376 -2916 -8238 -2484
rect -8142 2484 -8004 2916
rect -8142 -2916 -8004 -2484
rect -7908 2484 -7770 2916
rect -7908 -2916 -7770 -2484
rect -7674 2484 -7536 2916
rect -7674 -2916 -7536 -2484
rect -7440 2484 -7302 2916
rect -7440 -2916 -7302 -2484
rect -7206 2484 -7068 2916
rect -7206 -2916 -7068 -2484
rect -6972 2484 -6834 2916
rect -6972 -2916 -6834 -2484
rect -6738 2484 -6600 2916
rect -6738 -2916 -6600 -2484
rect -6504 2484 -6366 2916
rect -6504 -2916 -6366 -2484
rect -6270 2484 -6132 2916
rect -6270 -2916 -6132 -2484
rect -6036 2484 -5898 2916
rect -6036 -2916 -5898 -2484
rect -5802 2484 -5664 2916
rect -5802 -2916 -5664 -2484
rect -5568 2484 -5430 2916
rect -5568 -2916 -5430 -2484
rect -5334 2484 -5196 2916
rect -5334 -2916 -5196 -2484
rect -5100 2484 -4962 2916
rect -5100 -2916 -4962 -2484
rect -4866 2484 -4728 2916
rect -4866 -2916 -4728 -2484
rect -4632 2484 -4494 2916
rect -4632 -2916 -4494 -2484
rect -4398 2484 -4260 2916
rect -4398 -2916 -4260 -2484
rect -4164 2484 -4026 2916
rect -4164 -2916 -4026 -2484
rect -3930 2484 -3792 2916
rect -3930 -2916 -3792 -2484
rect -3696 2484 -3558 2916
rect -3696 -2916 -3558 -2484
rect -3462 2484 -3324 2916
rect -3462 -2916 -3324 -2484
rect -3228 2484 -3090 2916
rect -3228 -2916 -3090 -2484
rect -2994 2484 -2856 2916
rect -2994 -2916 -2856 -2484
rect -2760 2484 -2622 2916
rect -2760 -2916 -2622 -2484
rect -2526 2484 -2388 2916
rect -2526 -2916 -2388 -2484
rect -2292 2484 -2154 2916
rect -2292 -2916 -2154 -2484
rect -2058 2484 -1920 2916
rect -2058 -2916 -1920 -2484
rect -1824 2484 -1686 2916
rect -1824 -2916 -1686 -2484
rect -1590 2484 -1452 2916
rect -1590 -2916 -1452 -2484
rect -1356 2484 -1218 2916
rect -1356 -2916 -1218 -2484
rect -1122 2484 -984 2916
rect -1122 -2916 -984 -2484
rect -888 2484 -750 2916
rect -888 -2916 -750 -2484
rect -654 2484 -516 2916
rect -654 -2916 -516 -2484
rect -420 2484 -282 2916
rect -420 -2916 -282 -2484
rect -186 2484 -48 2916
rect -186 -2916 -48 -2484
rect 48 2484 186 2916
rect 48 -2916 186 -2484
rect 282 2484 420 2916
rect 282 -2916 420 -2484
rect 516 2484 654 2916
rect 516 -2916 654 -2484
rect 750 2484 888 2916
rect 750 -2916 888 -2484
rect 984 2484 1122 2916
rect 984 -2916 1122 -2484
rect 1218 2484 1356 2916
rect 1218 -2916 1356 -2484
rect 1452 2484 1590 2916
rect 1452 -2916 1590 -2484
rect 1686 2484 1824 2916
rect 1686 -2916 1824 -2484
rect 1920 2484 2058 2916
rect 1920 -2916 2058 -2484
rect 2154 2484 2292 2916
rect 2154 -2916 2292 -2484
rect 2388 2484 2526 2916
rect 2388 -2916 2526 -2484
rect 2622 2484 2760 2916
rect 2622 -2916 2760 -2484
rect 2856 2484 2994 2916
rect 2856 -2916 2994 -2484
rect 3090 2484 3228 2916
rect 3090 -2916 3228 -2484
rect 3324 2484 3462 2916
rect 3324 -2916 3462 -2484
rect 3558 2484 3696 2916
rect 3558 -2916 3696 -2484
rect 3792 2484 3930 2916
rect 3792 -2916 3930 -2484
rect 4026 2484 4164 2916
rect 4026 -2916 4164 -2484
rect 4260 2484 4398 2916
rect 4260 -2916 4398 -2484
rect 4494 2484 4632 2916
rect 4494 -2916 4632 -2484
rect 4728 2484 4866 2916
rect 4728 -2916 4866 -2484
rect 4962 2484 5100 2916
rect 4962 -2916 5100 -2484
rect 5196 2484 5334 2916
rect 5196 -2916 5334 -2484
rect 5430 2484 5568 2916
rect 5430 -2916 5568 -2484
rect 5664 2484 5802 2916
rect 5664 -2916 5802 -2484
rect 5898 2484 6036 2916
rect 5898 -2916 6036 -2484
rect 6132 2484 6270 2916
rect 6132 -2916 6270 -2484
rect 6366 2484 6504 2916
rect 6366 -2916 6504 -2484
rect 6600 2484 6738 2916
rect 6600 -2916 6738 -2484
rect 6834 2484 6972 2916
rect 6834 -2916 6972 -2484
rect 7068 2484 7206 2916
rect 7068 -2916 7206 -2484
rect 7302 2484 7440 2916
rect 7302 -2916 7440 -2484
rect 7536 2484 7674 2916
rect 7536 -2916 7674 -2484
rect 7770 2484 7908 2916
rect 7770 -2916 7908 -2484
rect 8004 2484 8142 2916
rect 8004 -2916 8142 -2484
rect 8238 2484 8376 2916
rect 8238 -2916 8376 -2484
rect 8472 2484 8610 2916
rect 8472 -2916 8610 -2484
rect 8706 2484 8844 2916
rect 8706 -2916 8844 -2484
rect 8940 2484 9078 2916
rect 8940 -2916 9078 -2484
rect 9174 2484 9312 2916
rect 9174 -2916 9312 -2484
rect 9408 2484 9546 2916
rect 9408 -2916 9546 -2484
rect 9642 2484 9780 2916
rect 9642 -2916 9780 -2484
rect 9876 2484 10014 2916
rect 9876 -2916 10014 -2484
rect 10110 2484 10248 2916
rect 10110 -2916 10248 -2484
rect 10344 2484 10482 2916
rect 10344 -2916 10482 -2484
rect 10578 2484 10716 2916
rect 10578 -2916 10716 -2484
rect 10812 2484 10950 2916
rect 10812 -2916 10950 -2484
rect 11046 2484 11184 2916
rect 11046 -2916 11184 -2484
rect 11280 2484 11418 2916
rect 11280 -2916 11418 -2484
rect 11514 2484 11652 2916
rect 11514 -2916 11652 -2484
rect 11748 2484 11886 2916
rect 11748 -2916 11886 -2484
rect 11982 2484 12120 2916
rect 11982 -2916 12120 -2484
rect 12216 2484 12354 2916
rect 12216 -2916 12354 -2484
rect 12450 2484 12588 2916
rect 12450 -2916 12588 -2484
rect 12684 2484 12822 2916
rect 12684 -2916 12822 -2484
rect 12918 2484 13056 2916
rect 12918 -2916 13056 -2484
rect 13152 2484 13290 2916
rect 13152 -2916 13290 -2484
rect 13386 2484 13524 2916
rect 13386 -2916 13524 -2484
rect 13620 2484 13758 2916
rect 13620 -2916 13758 -2484
rect 13854 2484 13992 2916
rect 13854 -2916 13992 -2484
rect 14088 2484 14226 2916
rect 14088 -2916 14226 -2484
rect 14322 2484 14460 2916
rect 14322 -2916 14460 -2484
rect 14556 2484 14694 2916
rect 14556 -2916 14694 -2484
rect 14790 2484 14928 2916
rect 14790 -2916 14928 -2484
rect 15024 2484 15162 2916
rect 15024 -2916 15162 -2484
rect 15258 2484 15396 2916
rect 15258 -2916 15396 -2484
rect 15492 2484 15630 2916
rect 15492 -2916 15630 -2484
rect 15726 2484 15864 2916
rect 15726 -2916 15864 -2484
rect 15960 2484 16098 2916
rect 15960 -2916 16098 -2484
rect 16194 2484 16332 2916
rect 16194 -2916 16332 -2484
rect 16428 2484 16566 2916
rect 16428 -2916 16566 -2484
rect 16662 2484 16800 2916
rect 16662 -2916 16800 -2484
rect 16896 2484 17034 2916
rect 16896 -2916 17034 -2484
rect 17130 2484 17268 2916
rect 17130 -2916 17268 -2484
rect 17364 2484 17502 2916
rect 17364 -2916 17502 -2484
rect 17598 2484 17736 2916
rect 17598 -2916 17736 -2484
rect 17832 2484 17970 2916
rect 17832 -2916 17970 -2484
rect 18066 2484 18204 2916
rect 18066 -2916 18204 -2484
rect 18300 2484 18438 2916
rect 18300 -2916 18438 -2484
rect 18534 2484 18672 2916
rect 18534 -2916 18672 -2484
rect 18768 2484 18906 2916
rect 18768 -2916 18906 -2484
rect 19002 2484 19140 2916
rect 19002 -2916 19140 -2484
rect 19236 2484 19374 2916
rect 19236 -2916 19374 -2484
rect 19470 2484 19608 2916
rect 19470 -2916 19608 -2484
rect 19704 2484 19842 2916
rect 19704 -2916 19842 -2484
rect 19938 2484 20076 2916
rect 19938 -2916 20076 -2484
rect 20172 2484 20310 2916
rect 20172 -2916 20310 -2484
rect 20406 2484 20544 2916
rect 20406 -2916 20544 -2484
rect 20640 2484 20778 2916
rect 20640 -2916 20778 -2484
rect 20874 2484 21012 2916
rect 20874 -2916 21012 -2484
rect 21108 2484 21246 2916
rect 21108 -2916 21246 -2484
rect 21342 2484 21480 2916
rect 21342 -2916 21480 -2484
rect 21576 2484 21714 2916
rect 21576 -2916 21714 -2484
rect 21810 2484 21948 2916
rect 21810 -2916 21948 -2484
rect 22044 2484 22182 2916
rect 22044 -2916 22182 -2484
rect 22278 2484 22416 2916
rect 22278 -2916 22416 -2484
rect 22512 2484 22650 2916
rect 22512 -2916 22650 -2484
rect 22746 2484 22884 2916
rect 22746 -2916 22884 -2484
rect 22980 2484 23118 2916
rect 22980 -2916 23118 -2484
rect 23214 2484 23352 2916
rect 23214 -2916 23352 -2484
rect 23448 2484 23586 2916
rect 23448 -2916 23586 -2484
rect 23682 2484 23820 2916
rect 23682 -2916 23820 -2484
rect 23916 2484 24054 2916
rect 23916 -2916 24054 -2484
rect 24150 2484 24288 2916
rect 24150 -2916 24288 -2484
rect 24384 2484 24522 2916
rect 24384 -2916 24522 -2484
rect 24618 2484 24756 2916
rect 24618 -2916 24756 -2484
rect 24852 2484 24990 2916
rect 24852 -2916 24990 -2484
rect 25086 2484 25224 2916
rect 25086 -2916 25224 -2484
rect 25320 2484 25458 2916
rect 25320 -2916 25458 -2484
rect 25554 2484 25692 2916
rect 25554 -2916 25692 -2484
rect 25788 2484 25926 2916
rect 25788 -2916 25926 -2484
rect 26022 2484 26160 2916
rect 26022 -2916 26160 -2484
rect 26256 2484 26394 2916
rect 26256 -2916 26394 -2484
rect 26490 2484 26628 2916
rect 26490 -2916 26628 -2484
rect 26724 2484 26862 2916
rect 26724 -2916 26862 -2484
rect 26958 2484 27096 2916
rect 26958 -2916 27096 -2484
rect 27192 2484 27330 2916
rect 27192 -2916 27330 -2484
rect 27426 2484 27564 2916
rect 27426 -2916 27564 -2484
rect 27660 2484 27798 2916
rect 27660 -2916 27798 -2484
rect 27894 2484 28032 2916
rect 27894 -2916 28032 -2484
rect 28128 2484 28266 2916
rect 28128 -2916 28266 -2484
rect 28362 2484 28500 2916
rect 28362 -2916 28500 -2484
rect 28596 2484 28734 2916
rect 28596 -2916 28734 -2484
rect 28830 2484 28968 2916
rect 28830 -2916 28968 -2484
rect 29064 2484 29202 2916
rect 29064 -2916 29202 -2484
rect 29298 2484 29436 2916
rect 29298 -2916 29436 -2484
rect 29532 2484 29670 2916
rect 29532 -2916 29670 -2484
rect 29766 2484 29904 2916
rect 29766 -2916 29904 -2484
<< ppolyres >>
rect -29904 -2484 -29766 2484
rect -29670 -2484 -29532 2484
rect -29436 -2484 -29298 2484
rect -29202 -2484 -29064 2484
rect -28968 -2484 -28830 2484
rect -28734 -2484 -28596 2484
rect -28500 -2484 -28362 2484
rect -28266 -2484 -28128 2484
rect -28032 -2484 -27894 2484
rect -27798 -2484 -27660 2484
rect -27564 -2484 -27426 2484
rect -27330 -2484 -27192 2484
rect -27096 -2484 -26958 2484
rect -26862 -2484 -26724 2484
rect -26628 -2484 -26490 2484
rect -26394 -2484 -26256 2484
rect -26160 -2484 -26022 2484
rect -25926 -2484 -25788 2484
rect -25692 -2484 -25554 2484
rect -25458 -2484 -25320 2484
rect -25224 -2484 -25086 2484
rect -24990 -2484 -24852 2484
rect -24756 -2484 -24618 2484
rect -24522 -2484 -24384 2484
rect -24288 -2484 -24150 2484
rect -24054 -2484 -23916 2484
rect -23820 -2484 -23682 2484
rect -23586 -2484 -23448 2484
rect -23352 -2484 -23214 2484
rect -23118 -2484 -22980 2484
rect -22884 -2484 -22746 2484
rect -22650 -2484 -22512 2484
rect -22416 -2484 -22278 2484
rect -22182 -2484 -22044 2484
rect -21948 -2484 -21810 2484
rect -21714 -2484 -21576 2484
rect -21480 -2484 -21342 2484
rect -21246 -2484 -21108 2484
rect -21012 -2484 -20874 2484
rect -20778 -2484 -20640 2484
rect -20544 -2484 -20406 2484
rect -20310 -2484 -20172 2484
rect -20076 -2484 -19938 2484
rect -19842 -2484 -19704 2484
rect -19608 -2484 -19470 2484
rect -19374 -2484 -19236 2484
rect -19140 -2484 -19002 2484
rect -18906 -2484 -18768 2484
rect -18672 -2484 -18534 2484
rect -18438 -2484 -18300 2484
rect -18204 -2484 -18066 2484
rect -17970 -2484 -17832 2484
rect -17736 -2484 -17598 2484
rect -17502 -2484 -17364 2484
rect -17268 -2484 -17130 2484
rect -17034 -2484 -16896 2484
rect -16800 -2484 -16662 2484
rect -16566 -2484 -16428 2484
rect -16332 -2484 -16194 2484
rect -16098 -2484 -15960 2484
rect -15864 -2484 -15726 2484
rect -15630 -2484 -15492 2484
rect -15396 -2484 -15258 2484
rect -15162 -2484 -15024 2484
rect -14928 -2484 -14790 2484
rect -14694 -2484 -14556 2484
rect -14460 -2484 -14322 2484
rect -14226 -2484 -14088 2484
rect -13992 -2484 -13854 2484
rect -13758 -2484 -13620 2484
rect -13524 -2484 -13386 2484
rect -13290 -2484 -13152 2484
rect -13056 -2484 -12918 2484
rect -12822 -2484 -12684 2484
rect -12588 -2484 -12450 2484
rect -12354 -2484 -12216 2484
rect -12120 -2484 -11982 2484
rect -11886 -2484 -11748 2484
rect -11652 -2484 -11514 2484
rect -11418 -2484 -11280 2484
rect -11184 -2484 -11046 2484
rect -10950 -2484 -10812 2484
rect -10716 -2484 -10578 2484
rect -10482 -2484 -10344 2484
rect -10248 -2484 -10110 2484
rect -10014 -2484 -9876 2484
rect -9780 -2484 -9642 2484
rect -9546 -2484 -9408 2484
rect -9312 -2484 -9174 2484
rect -9078 -2484 -8940 2484
rect -8844 -2484 -8706 2484
rect -8610 -2484 -8472 2484
rect -8376 -2484 -8238 2484
rect -8142 -2484 -8004 2484
rect -7908 -2484 -7770 2484
rect -7674 -2484 -7536 2484
rect -7440 -2484 -7302 2484
rect -7206 -2484 -7068 2484
rect -6972 -2484 -6834 2484
rect -6738 -2484 -6600 2484
rect -6504 -2484 -6366 2484
rect -6270 -2484 -6132 2484
rect -6036 -2484 -5898 2484
rect -5802 -2484 -5664 2484
rect -5568 -2484 -5430 2484
rect -5334 -2484 -5196 2484
rect -5100 -2484 -4962 2484
rect -4866 -2484 -4728 2484
rect -4632 -2484 -4494 2484
rect -4398 -2484 -4260 2484
rect -4164 -2484 -4026 2484
rect -3930 -2484 -3792 2484
rect -3696 -2484 -3558 2484
rect -3462 -2484 -3324 2484
rect -3228 -2484 -3090 2484
rect -2994 -2484 -2856 2484
rect -2760 -2484 -2622 2484
rect -2526 -2484 -2388 2484
rect -2292 -2484 -2154 2484
rect -2058 -2484 -1920 2484
rect -1824 -2484 -1686 2484
rect -1590 -2484 -1452 2484
rect -1356 -2484 -1218 2484
rect -1122 -2484 -984 2484
rect -888 -2484 -750 2484
rect -654 -2484 -516 2484
rect -420 -2484 -282 2484
rect -186 -2484 -48 2484
rect 48 -2484 186 2484
rect 282 -2484 420 2484
rect 516 -2484 654 2484
rect 750 -2484 888 2484
rect 984 -2484 1122 2484
rect 1218 -2484 1356 2484
rect 1452 -2484 1590 2484
rect 1686 -2484 1824 2484
rect 1920 -2484 2058 2484
rect 2154 -2484 2292 2484
rect 2388 -2484 2526 2484
rect 2622 -2484 2760 2484
rect 2856 -2484 2994 2484
rect 3090 -2484 3228 2484
rect 3324 -2484 3462 2484
rect 3558 -2484 3696 2484
rect 3792 -2484 3930 2484
rect 4026 -2484 4164 2484
rect 4260 -2484 4398 2484
rect 4494 -2484 4632 2484
rect 4728 -2484 4866 2484
rect 4962 -2484 5100 2484
rect 5196 -2484 5334 2484
rect 5430 -2484 5568 2484
rect 5664 -2484 5802 2484
rect 5898 -2484 6036 2484
rect 6132 -2484 6270 2484
rect 6366 -2484 6504 2484
rect 6600 -2484 6738 2484
rect 6834 -2484 6972 2484
rect 7068 -2484 7206 2484
rect 7302 -2484 7440 2484
rect 7536 -2484 7674 2484
rect 7770 -2484 7908 2484
rect 8004 -2484 8142 2484
rect 8238 -2484 8376 2484
rect 8472 -2484 8610 2484
rect 8706 -2484 8844 2484
rect 8940 -2484 9078 2484
rect 9174 -2484 9312 2484
rect 9408 -2484 9546 2484
rect 9642 -2484 9780 2484
rect 9876 -2484 10014 2484
rect 10110 -2484 10248 2484
rect 10344 -2484 10482 2484
rect 10578 -2484 10716 2484
rect 10812 -2484 10950 2484
rect 11046 -2484 11184 2484
rect 11280 -2484 11418 2484
rect 11514 -2484 11652 2484
rect 11748 -2484 11886 2484
rect 11982 -2484 12120 2484
rect 12216 -2484 12354 2484
rect 12450 -2484 12588 2484
rect 12684 -2484 12822 2484
rect 12918 -2484 13056 2484
rect 13152 -2484 13290 2484
rect 13386 -2484 13524 2484
rect 13620 -2484 13758 2484
rect 13854 -2484 13992 2484
rect 14088 -2484 14226 2484
rect 14322 -2484 14460 2484
rect 14556 -2484 14694 2484
rect 14790 -2484 14928 2484
rect 15024 -2484 15162 2484
rect 15258 -2484 15396 2484
rect 15492 -2484 15630 2484
rect 15726 -2484 15864 2484
rect 15960 -2484 16098 2484
rect 16194 -2484 16332 2484
rect 16428 -2484 16566 2484
rect 16662 -2484 16800 2484
rect 16896 -2484 17034 2484
rect 17130 -2484 17268 2484
rect 17364 -2484 17502 2484
rect 17598 -2484 17736 2484
rect 17832 -2484 17970 2484
rect 18066 -2484 18204 2484
rect 18300 -2484 18438 2484
rect 18534 -2484 18672 2484
rect 18768 -2484 18906 2484
rect 19002 -2484 19140 2484
rect 19236 -2484 19374 2484
rect 19470 -2484 19608 2484
rect 19704 -2484 19842 2484
rect 19938 -2484 20076 2484
rect 20172 -2484 20310 2484
rect 20406 -2484 20544 2484
rect 20640 -2484 20778 2484
rect 20874 -2484 21012 2484
rect 21108 -2484 21246 2484
rect 21342 -2484 21480 2484
rect 21576 -2484 21714 2484
rect 21810 -2484 21948 2484
rect 22044 -2484 22182 2484
rect 22278 -2484 22416 2484
rect 22512 -2484 22650 2484
rect 22746 -2484 22884 2484
rect 22980 -2484 23118 2484
rect 23214 -2484 23352 2484
rect 23448 -2484 23586 2484
rect 23682 -2484 23820 2484
rect 23916 -2484 24054 2484
rect 24150 -2484 24288 2484
rect 24384 -2484 24522 2484
rect 24618 -2484 24756 2484
rect 24852 -2484 24990 2484
rect 25086 -2484 25224 2484
rect 25320 -2484 25458 2484
rect 25554 -2484 25692 2484
rect 25788 -2484 25926 2484
rect 26022 -2484 26160 2484
rect 26256 -2484 26394 2484
rect 26490 -2484 26628 2484
rect 26724 -2484 26862 2484
rect 26958 -2484 27096 2484
rect 27192 -2484 27330 2484
rect 27426 -2484 27564 2484
rect 27660 -2484 27798 2484
rect 27894 -2484 28032 2484
rect 28128 -2484 28266 2484
rect 28362 -2484 28500 2484
rect 28596 -2484 28734 2484
rect 28830 -2484 28968 2484
rect 29064 -2484 29202 2484
rect 29298 -2484 29436 2484
rect 29532 -2484 29670 2484
rect 29766 -2484 29904 2484
<< locali >>
rect -30034 3012 -29938 3046
rect 29938 3012 30034 3046
rect -30034 2950 -30000 3012
rect 30000 2950 30034 3012
rect -30034 -3012 -30000 -2950
rect 30000 -3012 30034 -2950
rect -30034 -3046 -29938 -3012
rect 29938 -3046 30034 -3012
<< viali >>
rect -29888 2501 -29782 2898
rect -29654 2501 -29548 2898
rect -29420 2501 -29314 2898
rect -29186 2501 -29080 2898
rect -28952 2501 -28846 2898
rect -28718 2501 -28612 2898
rect -28484 2501 -28378 2898
rect -28250 2501 -28144 2898
rect -28016 2501 -27910 2898
rect -27782 2501 -27676 2898
rect -27548 2501 -27442 2898
rect -27314 2501 -27208 2898
rect -27080 2501 -26974 2898
rect -26846 2501 -26740 2898
rect -26612 2501 -26506 2898
rect -26378 2501 -26272 2898
rect -26144 2501 -26038 2898
rect -25910 2501 -25804 2898
rect -25676 2501 -25570 2898
rect -25442 2501 -25336 2898
rect -25208 2501 -25102 2898
rect -24974 2501 -24868 2898
rect -24740 2501 -24634 2898
rect -24506 2501 -24400 2898
rect -24272 2501 -24166 2898
rect -24038 2501 -23932 2898
rect -23804 2501 -23698 2898
rect -23570 2501 -23464 2898
rect -23336 2501 -23230 2898
rect -23102 2501 -22996 2898
rect -22868 2501 -22762 2898
rect -22634 2501 -22528 2898
rect -22400 2501 -22294 2898
rect -22166 2501 -22060 2898
rect -21932 2501 -21826 2898
rect -21698 2501 -21592 2898
rect -21464 2501 -21358 2898
rect -21230 2501 -21124 2898
rect -20996 2501 -20890 2898
rect -20762 2501 -20656 2898
rect -20528 2501 -20422 2898
rect -20294 2501 -20188 2898
rect -20060 2501 -19954 2898
rect -19826 2501 -19720 2898
rect -19592 2501 -19486 2898
rect -19358 2501 -19252 2898
rect -19124 2501 -19018 2898
rect -18890 2501 -18784 2898
rect -18656 2501 -18550 2898
rect -18422 2501 -18316 2898
rect -18188 2501 -18082 2898
rect -17954 2501 -17848 2898
rect -17720 2501 -17614 2898
rect -17486 2501 -17380 2898
rect -17252 2501 -17146 2898
rect -17018 2501 -16912 2898
rect -16784 2501 -16678 2898
rect -16550 2501 -16444 2898
rect -16316 2501 -16210 2898
rect -16082 2501 -15976 2898
rect -15848 2501 -15742 2898
rect -15614 2501 -15508 2898
rect -15380 2501 -15274 2898
rect -15146 2501 -15040 2898
rect -14912 2501 -14806 2898
rect -14678 2501 -14572 2898
rect -14444 2501 -14338 2898
rect -14210 2501 -14104 2898
rect -13976 2501 -13870 2898
rect -13742 2501 -13636 2898
rect -13508 2501 -13402 2898
rect -13274 2501 -13168 2898
rect -13040 2501 -12934 2898
rect -12806 2501 -12700 2898
rect -12572 2501 -12466 2898
rect -12338 2501 -12232 2898
rect -12104 2501 -11998 2898
rect -11870 2501 -11764 2898
rect -11636 2501 -11530 2898
rect -11402 2501 -11296 2898
rect -11168 2501 -11062 2898
rect -10934 2501 -10828 2898
rect -10700 2501 -10594 2898
rect -10466 2501 -10360 2898
rect -10232 2501 -10126 2898
rect -9998 2501 -9892 2898
rect -9764 2501 -9658 2898
rect -9530 2501 -9424 2898
rect -9296 2501 -9190 2898
rect -9062 2501 -8956 2898
rect -8828 2501 -8722 2898
rect -8594 2501 -8488 2898
rect -8360 2501 -8254 2898
rect -8126 2501 -8020 2898
rect -7892 2501 -7786 2898
rect -7658 2501 -7552 2898
rect -7424 2501 -7318 2898
rect -7190 2501 -7084 2898
rect -6956 2501 -6850 2898
rect -6722 2501 -6616 2898
rect -6488 2501 -6382 2898
rect -6254 2501 -6148 2898
rect -6020 2501 -5914 2898
rect -5786 2501 -5680 2898
rect -5552 2501 -5446 2898
rect -5318 2501 -5212 2898
rect -5084 2501 -4978 2898
rect -4850 2501 -4744 2898
rect -4616 2501 -4510 2898
rect -4382 2501 -4276 2898
rect -4148 2501 -4042 2898
rect -3914 2501 -3808 2898
rect -3680 2501 -3574 2898
rect -3446 2501 -3340 2898
rect -3212 2501 -3106 2898
rect -2978 2501 -2872 2898
rect -2744 2501 -2638 2898
rect -2510 2501 -2404 2898
rect -2276 2501 -2170 2898
rect -2042 2501 -1936 2898
rect -1808 2501 -1702 2898
rect -1574 2501 -1468 2898
rect -1340 2501 -1234 2898
rect -1106 2501 -1000 2898
rect -872 2501 -766 2898
rect -638 2501 -532 2898
rect -404 2501 -298 2898
rect -170 2501 -64 2898
rect 64 2501 170 2898
rect 298 2501 404 2898
rect 532 2501 638 2898
rect 766 2501 872 2898
rect 1000 2501 1106 2898
rect 1234 2501 1340 2898
rect 1468 2501 1574 2898
rect 1702 2501 1808 2898
rect 1936 2501 2042 2898
rect 2170 2501 2276 2898
rect 2404 2501 2510 2898
rect 2638 2501 2744 2898
rect 2872 2501 2978 2898
rect 3106 2501 3212 2898
rect 3340 2501 3446 2898
rect 3574 2501 3680 2898
rect 3808 2501 3914 2898
rect 4042 2501 4148 2898
rect 4276 2501 4382 2898
rect 4510 2501 4616 2898
rect 4744 2501 4850 2898
rect 4978 2501 5084 2898
rect 5212 2501 5318 2898
rect 5446 2501 5552 2898
rect 5680 2501 5786 2898
rect 5914 2501 6020 2898
rect 6148 2501 6254 2898
rect 6382 2501 6488 2898
rect 6616 2501 6722 2898
rect 6850 2501 6956 2898
rect 7084 2501 7190 2898
rect 7318 2501 7424 2898
rect 7552 2501 7658 2898
rect 7786 2501 7892 2898
rect 8020 2501 8126 2898
rect 8254 2501 8360 2898
rect 8488 2501 8594 2898
rect 8722 2501 8828 2898
rect 8956 2501 9062 2898
rect 9190 2501 9296 2898
rect 9424 2501 9530 2898
rect 9658 2501 9764 2898
rect 9892 2501 9998 2898
rect 10126 2501 10232 2898
rect 10360 2501 10466 2898
rect 10594 2501 10700 2898
rect 10828 2501 10934 2898
rect 11062 2501 11168 2898
rect 11296 2501 11402 2898
rect 11530 2501 11636 2898
rect 11764 2501 11870 2898
rect 11998 2501 12104 2898
rect 12232 2501 12338 2898
rect 12466 2501 12572 2898
rect 12700 2501 12806 2898
rect 12934 2501 13040 2898
rect 13168 2501 13274 2898
rect 13402 2501 13508 2898
rect 13636 2501 13742 2898
rect 13870 2501 13976 2898
rect 14104 2501 14210 2898
rect 14338 2501 14444 2898
rect 14572 2501 14678 2898
rect 14806 2501 14912 2898
rect 15040 2501 15146 2898
rect 15274 2501 15380 2898
rect 15508 2501 15614 2898
rect 15742 2501 15848 2898
rect 15976 2501 16082 2898
rect 16210 2501 16316 2898
rect 16444 2501 16550 2898
rect 16678 2501 16784 2898
rect 16912 2501 17018 2898
rect 17146 2501 17252 2898
rect 17380 2501 17486 2898
rect 17614 2501 17720 2898
rect 17848 2501 17954 2898
rect 18082 2501 18188 2898
rect 18316 2501 18422 2898
rect 18550 2501 18656 2898
rect 18784 2501 18890 2898
rect 19018 2501 19124 2898
rect 19252 2501 19358 2898
rect 19486 2501 19592 2898
rect 19720 2501 19826 2898
rect 19954 2501 20060 2898
rect 20188 2501 20294 2898
rect 20422 2501 20528 2898
rect 20656 2501 20762 2898
rect 20890 2501 20996 2898
rect 21124 2501 21230 2898
rect 21358 2501 21464 2898
rect 21592 2501 21698 2898
rect 21826 2501 21932 2898
rect 22060 2501 22166 2898
rect 22294 2501 22400 2898
rect 22528 2501 22634 2898
rect 22762 2501 22868 2898
rect 22996 2501 23102 2898
rect 23230 2501 23336 2898
rect 23464 2501 23570 2898
rect 23698 2501 23804 2898
rect 23932 2501 24038 2898
rect 24166 2501 24272 2898
rect 24400 2501 24506 2898
rect 24634 2501 24740 2898
rect 24868 2501 24974 2898
rect 25102 2501 25208 2898
rect 25336 2501 25442 2898
rect 25570 2501 25676 2898
rect 25804 2501 25910 2898
rect 26038 2501 26144 2898
rect 26272 2501 26378 2898
rect 26506 2501 26612 2898
rect 26740 2501 26846 2898
rect 26974 2501 27080 2898
rect 27208 2501 27314 2898
rect 27442 2501 27548 2898
rect 27676 2501 27782 2898
rect 27910 2501 28016 2898
rect 28144 2501 28250 2898
rect 28378 2501 28484 2898
rect 28612 2501 28718 2898
rect 28846 2501 28952 2898
rect 29080 2501 29186 2898
rect 29314 2501 29420 2898
rect 29548 2501 29654 2898
rect 29782 2501 29888 2898
rect -29888 -2898 -29782 -2501
rect -29654 -2898 -29548 -2501
rect -29420 -2898 -29314 -2501
rect -29186 -2898 -29080 -2501
rect -28952 -2898 -28846 -2501
rect -28718 -2898 -28612 -2501
rect -28484 -2898 -28378 -2501
rect -28250 -2898 -28144 -2501
rect -28016 -2898 -27910 -2501
rect -27782 -2898 -27676 -2501
rect -27548 -2898 -27442 -2501
rect -27314 -2898 -27208 -2501
rect -27080 -2898 -26974 -2501
rect -26846 -2898 -26740 -2501
rect -26612 -2898 -26506 -2501
rect -26378 -2898 -26272 -2501
rect -26144 -2898 -26038 -2501
rect -25910 -2898 -25804 -2501
rect -25676 -2898 -25570 -2501
rect -25442 -2898 -25336 -2501
rect -25208 -2898 -25102 -2501
rect -24974 -2898 -24868 -2501
rect -24740 -2898 -24634 -2501
rect -24506 -2898 -24400 -2501
rect -24272 -2898 -24166 -2501
rect -24038 -2898 -23932 -2501
rect -23804 -2898 -23698 -2501
rect -23570 -2898 -23464 -2501
rect -23336 -2898 -23230 -2501
rect -23102 -2898 -22996 -2501
rect -22868 -2898 -22762 -2501
rect -22634 -2898 -22528 -2501
rect -22400 -2898 -22294 -2501
rect -22166 -2898 -22060 -2501
rect -21932 -2898 -21826 -2501
rect -21698 -2898 -21592 -2501
rect -21464 -2898 -21358 -2501
rect -21230 -2898 -21124 -2501
rect -20996 -2898 -20890 -2501
rect -20762 -2898 -20656 -2501
rect -20528 -2898 -20422 -2501
rect -20294 -2898 -20188 -2501
rect -20060 -2898 -19954 -2501
rect -19826 -2898 -19720 -2501
rect -19592 -2898 -19486 -2501
rect -19358 -2898 -19252 -2501
rect -19124 -2898 -19018 -2501
rect -18890 -2898 -18784 -2501
rect -18656 -2898 -18550 -2501
rect -18422 -2898 -18316 -2501
rect -18188 -2898 -18082 -2501
rect -17954 -2898 -17848 -2501
rect -17720 -2898 -17614 -2501
rect -17486 -2898 -17380 -2501
rect -17252 -2898 -17146 -2501
rect -17018 -2898 -16912 -2501
rect -16784 -2898 -16678 -2501
rect -16550 -2898 -16444 -2501
rect -16316 -2898 -16210 -2501
rect -16082 -2898 -15976 -2501
rect -15848 -2898 -15742 -2501
rect -15614 -2898 -15508 -2501
rect -15380 -2898 -15274 -2501
rect -15146 -2898 -15040 -2501
rect -14912 -2898 -14806 -2501
rect -14678 -2898 -14572 -2501
rect -14444 -2898 -14338 -2501
rect -14210 -2898 -14104 -2501
rect -13976 -2898 -13870 -2501
rect -13742 -2898 -13636 -2501
rect -13508 -2898 -13402 -2501
rect -13274 -2898 -13168 -2501
rect -13040 -2898 -12934 -2501
rect -12806 -2898 -12700 -2501
rect -12572 -2898 -12466 -2501
rect -12338 -2898 -12232 -2501
rect -12104 -2898 -11998 -2501
rect -11870 -2898 -11764 -2501
rect -11636 -2898 -11530 -2501
rect -11402 -2898 -11296 -2501
rect -11168 -2898 -11062 -2501
rect -10934 -2898 -10828 -2501
rect -10700 -2898 -10594 -2501
rect -10466 -2898 -10360 -2501
rect -10232 -2898 -10126 -2501
rect -9998 -2898 -9892 -2501
rect -9764 -2898 -9658 -2501
rect -9530 -2898 -9424 -2501
rect -9296 -2898 -9190 -2501
rect -9062 -2898 -8956 -2501
rect -8828 -2898 -8722 -2501
rect -8594 -2898 -8488 -2501
rect -8360 -2898 -8254 -2501
rect -8126 -2898 -8020 -2501
rect -7892 -2898 -7786 -2501
rect -7658 -2898 -7552 -2501
rect -7424 -2898 -7318 -2501
rect -7190 -2898 -7084 -2501
rect -6956 -2898 -6850 -2501
rect -6722 -2898 -6616 -2501
rect -6488 -2898 -6382 -2501
rect -6254 -2898 -6148 -2501
rect -6020 -2898 -5914 -2501
rect -5786 -2898 -5680 -2501
rect -5552 -2898 -5446 -2501
rect -5318 -2898 -5212 -2501
rect -5084 -2898 -4978 -2501
rect -4850 -2898 -4744 -2501
rect -4616 -2898 -4510 -2501
rect -4382 -2898 -4276 -2501
rect -4148 -2898 -4042 -2501
rect -3914 -2898 -3808 -2501
rect -3680 -2898 -3574 -2501
rect -3446 -2898 -3340 -2501
rect -3212 -2898 -3106 -2501
rect -2978 -2898 -2872 -2501
rect -2744 -2898 -2638 -2501
rect -2510 -2898 -2404 -2501
rect -2276 -2898 -2170 -2501
rect -2042 -2898 -1936 -2501
rect -1808 -2898 -1702 -2501
rect -1574 -2898 -1468 -2501
rect -1340 -2898 -1234 -2501
rect -1106 -2898 -1000 -2501
rect -872 -2898 -766 -2501
rect -638 -2898 -532 -2501
rect -404 -2898 -298 -2501
rect -170 -2898 -64 -2501
rect 64 -2898 170 -2501
rect 298 -2898 404 -2501
rect 532 -2898 638 -2501
rect 766 -2898 872 -2501
rect 1000 -2898 1106 -2501
rect 1234 -2898 1340 -2501
rect 1468 -2898 1574 -2501
rect 1702 -2898 1808 -2501
rect 1936 -2898 2042 -2501
rect 2170 -2898 2276 -2501
rect 2404 -2898 2510 -2501
rect 2638 -2898 2744 -2501
rect 2872 -2898 2978 -2501
rect 3106 -2898 3212 -2501
rect 3340 -2898 3446 -2501
rect 3574 -2898 3680 -2501
rect 3808 -2898 3914 -2501
rect 4042 -2898 4148 -2501
rect 4276 -2898 4382 -2501
rect 4510 -2898 4616 -2501
rect 4744 -2898 4850 -2501
rect 4978 -2898 5084 -2501
rect 5212 -2898 5318 -2501
rect 5446 -2898 5552 -2501
rect 5680 -2898 5786 -2501
rect 5914 -2898 6020 -2501
rect 6148 -2898 6254 -2501
rect 6382 -2898 6488 -2501
rect 6616 -2898 6722 -2501
rect 6850 -2898 6956 -2501
rect 7084 -2898 7190 -2501
rect 7318 -2898 7424 -2501
rect 7552 -2898 7658 -2501
rect 7786 -2898 7892 -2501
rect 8020 -2898 8126 -2501
rect 8254 -2898 8360 -2501
rect 8488 -2898 8594 -2501
rect 8722 -2898 8828 -2501
rect 8956 -2898 9062 -2501
rect 9190 -2898 9296 -2501
rect 9424 -2898 9530 -2501
rect 9658 -2898 9764 -2501
rect 9892 -2898 9998 -2501
rect 10126 -2898 10232 -2501
rect 10360 -2898 10466 -2501
rect 10594 -2898 10700 -2501
rect 10828 -2898 10934 -2501
rect 11062 -2898 11168 -2501
rect 11296 -2898 11402 -2501
rect 11530 -2898 11636 -2501
rect 11764 -2898 11870 -2501
rect 11998 -2898 12104 -2501
rect 12232 -2898 12338 -2501
rect 12466 -2898 12572 -2501
rect 12700 -2898 12806 -2501
rect 12934 -2898 13040 -2501
rect 13168 -2898 13274 -2501
rect 13402 -2898 13508 -2501
rect 13636 -2898 13742 -2501
rect 13870 -2898 13976 -2501
rect 14104 -2898 14210 -2501
rect 14338 -2898 14444 -2501
rect 14572 -2898 14678 -2501
rect 14806 -2898 14912 -2501
rect 15040 -2898 15146 -2501
rect 15274 -2898 15380 -2501
rect 15508 -2898 15614 -2501
rect 15742 -2898 15848 -2501
rect 15976 -2898 16082 -2501
rect 16210 -2898 16316 -2501
rect 16444 -2898 16550 -2501
rect 16678 -2898 16784 -2501
rect 16912 -2898 17018 -2501
rect 17146 -2898 17252 -2501
rect 17380 -2898 17486 -2501
rect 17614 -2898 17720 -2501
rect 17848 -2898 17954 -2501
rect 18082 -2898 18188 -2501
rect 18316 -2898 18422 -2501
rect 18550 -2898 18656 -2501
rect 18784 -2898 18890 -2501
rect 19018 -2898 19124 -2501
rect 19252 -2898 19358 -2501
rect 19486 -2898 19592 -2501
rect 19720 -2898 19826 -2501
rect 19954 -2898 20060 -2501
rect 20188 -2898 20294 -2501
rect 20422 -2898 20528 -2501
rect 20656 -2898 20762 -2501
rect 20890 -2898 20996 -2501
rect 21124 -2898 21230 -2501
rect 21358 -2898 21464 -2501
rect 21592 -2898 21698 -2501
rect 21826 -2898 21932 -2501
rect 22060 -2898 22166 -2501
rect 22294 -2898 22400 -2501
rect 22528 -2898 22634 -2501
rect 22762 -2898 22868 -2501
rect 22996 -2898 23102 -2501
rect 23230 -2898 23336 -2501
rect 23464 -2898 23570 -2501
rect 23698 -2898 23804 -2501
rect 23932 -2898 24038 -2501
rect 24166 -2898 24272 -2501
rect 24400 -2898 24506 -2501
rect 24634 -2898 24740 -2501
rect 24868 -2898 24974 -2501
rect 25102 -2898 25208 -2501
rect 25336 -2898 25442 -2501
rect 25570 -2898 25676 -2501
rect 25804 -2898 25910 -2501
rect 26038 -2898 26144 -2501
rect 26272 -2898 26378 -2501
rect 26506 -2898 26612 -2501
rect 26740 -2898 26846 -2501
rect 26974 -2898 27080 -2501
rect 27208 -2898 27314 -2501
rect 27442 -2898 27548 -2501
rect 27676 -2898 27782 -2501
rect 27910 -2898 28016 -2501
rect 28144 -2898 28250 -2501
rect 28378 -2898 28484 -2501
rect 28612 -2898 28718 -2501
rect 28846 -2898 28952 -2501
rect 29080 -2898 29186 -2501
rect 29314 -2898 29420 -2501
rect 29548 -2898 29654 -2501
rect 29782 -2898 29888 -2501
<< metal1 >>
rect -29894 2898 -29776 2910
rect -29894 2501 -29888 2898
rect -29782 2501 -29776 2898
rect -29894 2489 -29776 2501
rect -29660 2898 -29542 2910
rect -29660 2501 -29654 2898
rect -29548 2501 -29542 2898
rect -29660 2489 -29542 2501
rect -29426 2898 -29308 2910
rect -29426 2501 -29420 2898
rect -29314 2501 -29308 2898
rect -29426 2489 -29308 2501
rect -29192 2898 -29074 2910
rect -29192 2501 -29186 2898
rect -29080 2501 -29074 2898
rect -29192 2489 -29074 2501
rect -28958 2898 -28840 2910
rect -28958 2501 -28952 2898
rect -28846 2501 -28840 2898
rect -28958 2489 -28840 2501
rect -28724 2898 -28606 2910
rect -28724 2501 -28718 2898
rect -28612 2501 -28606 2898
rect -28724 2489 -28606 2501
rect -28490 2898 -28372 2910
rect -28490 2501 -28484 2898
rect -28378 2501 -28372 2898
rect -28490 2489 -28372 2501
rect -28256 2898 -28138 2910
rect -28256 2501 -28250 2898
rect -28144 2501 -28138 2898
rect -28256 2489 -28138 2501
rect -28022 2898 -27904 2910
rect -28022 2501 -28016 2898
rect -27910 2501 -27904 2898
rect -28022 2489 -27904 2501
rect -27788 2898 -27670 2910
rect -27788 2501 -27782 2898
rect -27676 2501 -27670 2898
rect -27788 2489 -27670 2501
rect -27554 2898 -27436 2910
rect -27554 2501 -27548 2898
rect -27442 2501 -27436 2898
rect -27554 2489 -27436 2501
rect -27320 2898 -27202 2910
rect -27320 2501 -27314 2898
rect -27208 2501 -27202 2898
rect -27320 2489 -27202 2501
rect -27086 2898 -26968 2910
rect -27086 2501 -27080 2898
rect -26974 2501 -26968 2898
rect -27086 2489 -26968 2501
rect -26852 2898 -26734 2910
rect -26852 2501 -26846 2898
rect -26740 2501 -26734 2898
rect -26852 2489 -26734 2501
rect -26618 2898 -26500 2910
rect -26618 2501 -26612 2898
rect -26506 2501 -26500 2898
rect -26618 2489 -26500 2501
rect -26384 2898 -26266 2910
rect -26384 2501 -26378 2898
rect -26272 2501 -26266 2898
rect -26384 2489 -26266 2501
rect -26150 2898 -26032 2910
rect -26150 2501 -26144 2898
rect -26038 2501 -26032 2898
rect -26150 2489 -26032 2501
rect -25916 2898 -25798 2910
rect -25916 2501 -25910 2898
rect -25804 2501 -25798 2898
rect -25916 2489 -25798 2501
rect -25682 2898 -25564 2910
rect -25682 2501 -25676 2898
rect -25570 2501 -25564 2898
rect -25682 2489 -25564 2501
rect -25448 2898 -25330 2910
rect -25448 2501 -25442 2898
rect -25336 2501 -25330 2898
rect -25448 2489 -25330 2501
rect -25214 2898 -25096 2910
rect -25214 2501 -25208 2898
rect -25102 2501 -25096 2898
rect -25214 2489 -25096 2501
rect -24980 2898 -24862 2910
rect -24980 2501 -24974 2898
rect -24868 2501 -24862 2898
rect -24980 2489 -24862 2501
rect -24746 2898 -24628 2910
rect -24746 2501 -24740 2898
rect -24634 2501 -24628 2898
rect -24746 2489 -24628 2501
rect -24512 2898 -24394 2910
rect -24512 2501 -24506 2898
rect -24400 2501 -24394 2898
rect -24512 2489 -24394 2501
rect -24278 2898 -24160 2910
rect -24278 2501 -24272 2898
rect -24166 2501 -24160 2898
rect -24278 2489 -24160 2501
rect -24044 2898 -23926 2910
rect -24044 2501 -24038 2898
rect -23932 2501 -23926 2898
rect -24044 2489 -23926 2501
rect -23810 2898 -23692 2910
rect -23810 2501 -23804 2898
rect -23698 2501 -23692 2898
rect -23810 2489 -23692 2501
rect -23576 2898 -23458 2910
rect -23576 2501 -23570 2898
rect -23464 2501 -23458 2898
rect -23576 2489 -23458 2501
rect -23342 2898 -23224 2910
rect -23342 2501 -23336 2898
rect -23230 2501 -23224 2898
rect -23342 2489 -23224 2501
rect -23108 2898 -22990 2910
rect -23108 2501 -23102 2898
rect -22996 2501 -22990 2898
rect -23108 2489 -22990 2501
rect -22874 2898 -22756 2910
rect -22874 2501 -22868 2898
rect -22762 2501 -22756 2898
rect -22874 2489 -22756 2501
rect -22640 2898 -22522 2910
rect -22640 2501 -22634 2898
rect -22528 2501 -22522 2898
rect -22640 2489 -22522 2501
rect -22406 2898 -22288 2910
rect -22406 2501 -22400 2898
rect -22294 2501 -22288 2898
rect -22406 2489 -22288 2501
rect -22172 2898 -22054 2910
rect -22172 2501 -22166 2898
rect -22060 2501 -22054 2898
rect -22172 2489 -22054 2501
rect -21938 2898 -21820 2910
rect -21938 2501 -21932 2898
rect -21826 2501 -21820 2898
rect -21938 2489 -21820 2501
rect -21704 2898 -21586 2910
rect -21704 2501 -21698 2898
rect -21592 2501 -21586 2898
rect -21704 2489 -21586 2501
rect -21470 2898 -21352 2910
rect -21470 2501 -21464 2898
rect -21358 2501 -21352 2898
rect -21470 2489 -21352 2501
rect -21236 2898 -21118 2910
rect -21236 2501 -21230 2898
rect -21124 2501 -21118 2898
rect -21236 2489 -21118 2501
rect -21002 2898 -20884 2910
rect -21002 2501 -20996 2898
rect -20890 2501 -20884 2898
rect -21002 2489 -20884 2501
rect -20768 2898 -20650 2910
rect -20768 2501 -20762 2898
rect -20656 2501 -20650 2898
rect -20768 2489 -20650 2501
rect -20534 2898 -20416 2910
rect -20534 2501 -20528 2898
rect -20422 2501 -20416 2898
rect -20534 2489 -20416 2501
rect -20300 2898 -20182 2910
rect -20300 2501 -20294 2898
rect -20188 2501 -20182 2898
rect -20300 2489 -20182 2501
rect -20066 2898 -19948 2910
rect -20066 2501 -20060 2898
rect -19954 2501 -19948 2898
rect -20066 2489 -19948 2501
rect -19832 2898 -19714 2910
rect -19832 2501 -19826 2898
rect -19720 2501 -19714 2898
rect -19832 2489 -19714 2501
rect -19598 2898 -19480 2910
rect -19598 2501 -19592 2898
rect -19486 2501 -19480 2898
rect -19598 2489 -19480 2501
rect -19364 2898 -19246 2910
rect -19364 2501 -19358 2898
rect -19252 2501 -19246 2898
rect -19364 2489 -19246 2501
rect -19130 2898 -19012 2910
rect -19130 2501 -19124 2898
rect -19018 2501 -19012 2898
rect -19130 2489 -19012 2501
rect -18896 2898 -18778 2910
rect -18896 2501 -18890 2898
rect -18784 2501 -18778 2898
rect -18896 2489 -18778 2501
rect -18662 2898 -18544 2910
rect -18662 2501 -18656 2898
rect -18550 2501 -18544 2898
rect -18662 2489 -18544 2501
rect -18428 2898 -18310 2910
rect -18428 2501 -18422 2898
rect -18316 2501 -18310 2898
rect -18428 2489 -18310 2501
rect -18194 2898 -18076 2910
rect -18194 2501 -18188 2898
rect -18082 2501 -18076 2898
rect -18194 2489 -18076 2501
rect -17960 2898 -17842 2910
rect -17960 2501 -17954 2898
rect -17848 2501 -17842 2898
rect -17960 2489 -17842 2501
rect -17726 2898 -17608 2910
rect -17726 2501 -17720 2898
rect -17614 2501 -17608 2898
rect -17726 2489 -17608 2501
rect -17492 2898 -17374 2910
rect -17492 2501 -17486 2898
rect -17380 2501 -17374 2898
rect -17492 2489 -17374 2501
rect -17258 2898 -17140 2910
rect -17258 2501 -17252 2898
rect -17146 2501 -17140 2898
rect -17258 2489 -17140 2501
rect -17024 2898 -16906 2910
rect -17024 2501 -17018 2898
rect -16912 2501 -16906 2898
rect -17024 2489 -16906 2501
rect -16790 2898 -16672 2910
rect -16790 2501 -16784 2898
rect -16678 2501 -16672 2898
rect -16790 2489 -16672 2501
rect -16556 2898 -16438 2910
rect -16556 2501 -16550 2898
rect -16444 2501 -16438 2898
rect -16556 2489 -16438 2501
rect -16322 2898 -16204 2910
rect -16322 2501 -16316 2898
rect -16210 2501 -16204 2898
rect -16322 2489 -16204 2501
rect -16088 2898 -15970 2910
rect -16088 2501 -16082 2898
rect -15976 2501 -15970 2898
rect -16088 2489 -15970 2501
rect -15854 2898 -15736 2910
rect -15854 2501 -15848 2898
rect -15742 2501 -15736 2898
rect -15854 2489 -15736 2501
rect -15620 2898 -15502 2910
rect -15620 2501 -15614 2898
rect -15508 2501 -15502 2898
rect -15620 2489 -15502 2501
rect -15386 2898 -15268 2910
rect -15386 2501 -15380 2898
rect -15274 2501 -15268 2898
rect -15386 2489 -15268 2501
rect -15152 2898 -15034 2910
rect -15152 2501 -15146 2898
rect -15040 2501 -15034 2898
rect -15152 2489 -15034 2501
rect -14918 2898 -14800 2910
rect -14918 2501 -14912 2898
rect -14806 2501 -14800 2898
rect -14918 2489 -14800 2501
rect -14684 2898 -14566 2910
rect -14684 2501 -14678 2898
rect -14572 2501 -14566 2898
rect -14684 2489 -14566 2501
rect -14450 2898 -14332 2910
rect -14450 2501 -14444 2898
rect -14338 2501 -14332 2898
rect -14450 2489 -14332 2501
rect -14216 2898 -14098 2910
rect -14216 2501 -14210 2898
rect -14104 2501 -14098 2898
rect -14216 2489 -14098 2501
rect -13982 2898 -13864 2910
rect -13982 2501 -13976 2898
rect -13870 2501 -13864 2898
rect -13982 2489 -13864 2501
rect -13748 2898 -13630 2910
rect -13748 2501 -13742 2898
rect -13636 2501 -13630 2898
rect -13748 2489 -13630 2501
rect -13514 2898 -13396 2910
rect -13514 2501 -13508 2898
rect -13402 2501 -13396 2898
rect -13514 2489 -13396 2501
rect -13280 2898 -13162 2910
rect -13280 2501 -13274 2898
rect -13168 2501 -13162 2898
rect -13280 2489 -13162 2501
rect -13046 2898 -12928 2910
rect -13046 2501 -13040 2898
rect -12934 2501 -12928 2898
rect -13046 2489 -12928 2501
rect -12812 2898 -12694 2910
rect -12812 2501 -12806 2898
rect -12700 2501 -12694 2898
rect -12812 2489 -12694 2501
rect -12578 2898 -12460 2910
rect -12578 2501 -12572 2898
rect -12466 2501 -12460 2898
rect -12578 2489 -12460 2501
rect -12344 2898 -12226 2910
rect -12344 2501 -12338 2898
rect -12232 2501 -12226 2898
rect -12344 2489 -12226 2501
rect -12110 2898 -11992 2910
rect -12110 2501 -12104 2898
rect -11998 2501 -11992 2898
rect -12110 2489 -11992 2501
rect -11876 2898 -11758 2910
rect -11876 2501 -11870 2898
rect -11764 2501 -11758 2898
rect -11876 2489 -11758 2501
rect -11642 2898 -11524 2910
rect -11642 2501 -11636 2898
rect -11530 2501 -11524 2898
rect -11642 2489 -11524 2501
rect -11408 2898 -11290 2910
rect -11408 2501 -11402 2898
rect -11296 2501 -11290 2898
rect -11408 2489 -11290 2501
rect -11174 2898 -11056 2910
rect -11174 2501 -11168 2898
rect -11062 2501 -11056 2898
rect -11174 2489 -11056 2501
rect -10940 2898 -10822 2910
rect -10940 2501 -10934 2898
rect -10828 2501 -10822 2898
rect -10940 2489 -10822 2501
rect -10706 2898 -10588 2910
rect -10706 2501 -10700 2898
rect -10594 2501 -10588 2898
rect -10706 2489 -10588 2501
rect -10472 2898 -10354 2910
rect -10472 2501 -10466 2898
rect -10360 2501 -10354 2898
rect -10472 2489 -10354 2501
rect -10238 2898 -10120 2910
rect -10238 2501 -10232 2898
rect -10126 2501 -10120 2898
rect -10238 2489 -10120 2501
rect -10004 2898 -9886 2910
rect -10004 2501 -9998 2898
rect -9892 2501 -9886 2898
rect -10004 2489 -9886 2501
rect -9770 2898 -9652 2910
rect -9770 2501 -9764 2898
rect -9658 2501 -9652 2898
rect -9770 2489 -9652 2501
rect -9536 2898 -9418 2910
rect -9536 2501 -9530 2898
rect -9424 2501 -9418 2898
rect -9536 2489 -9418 2501
rect -9302 2898 -9184 2910
rect -9302 2501 -9296 2898
rect -9190 2501 -9184 2898
rect -9302 2489 -9184 2501
rect -9068 2898 -8950 2910
rect -9068 2501 -9062 2898
rect -8956 2501 -8950 2898
rect -9068 2489 -8950 2501
rect -8834 2898 -8716 2910
rect -8834 2501 -8828 2898
rect -8722 2501 -8716 2898
rect -8834 2489 -8716 2501
rect -8600 2898 -8482 2910
rect -8600 2501 -8594 2898
rect -8488 2501 -8482 2898
rect -8600 2489 -8482 2501
rect -8366 2898 -8248 2910
rect -8366 2501 -8360 2898
rect -8254 2501 -8248 2898
rect -8366 2489 -8248 2501
rect -8132 2898 -8014 2910
rect -8132 2501 -8126 2898
rect -8020 2501 -8014 2898
rect -8132 2489 -8014 2501
rect -7898 2898 -7780 2910
rect -7898 2501 -7892 2898
rect -7786 2501 -7780 2898
rect -7898 2489 -7780 2501
rect -7664 2898 -7546 2910
rect -7664 2501 -7658 2898
rect -7552 2501 -7546 2898
rect -7664 2489 -7546 2501
rect -7430 2898 -7312 2910
rect -7430 2501 -7424 2898
rect -7318 2501 -7312 2898
rect -7430 2489 -7312 2501
rect -7196 2898 -7078 2910
rect -7196 2501 -7190 2898
rect -7084 2501 -7078 2898
rect -7196 2489 -7078 2501
rect -6962 2898 -6844 2910
rect -6962 2501 -6956 2898
rect -6850 2501 -6844 2898
rect -6962 2489 -6844 2501
rect -6728 2898 -6610 2910
rect -6728 2501 -6722 2898
rect -6616 2501 -6610 2898
rect -6728 2489 -6610 2501
rect -6494 2898 -6376 2910
rect -6494 2501 -6488 2898
rect -6382 2501 -6376 2898
rect -6494 2489 -6376 2501
rect -6260 2898 -6142 2910
rect -6260 2501 -6254 2898
rect -6148 2501 -6142 2898
rect -6260 2489 -6142 2501
rect -6026 2898 -5908 2910
rect -6026 2501 -6020 2898
rect -5914 2501 -5908 2898
rect -6026 2489 -5908 2501
rect -5792 2898 -5674 2910
rect -5792 2501 -5786 2898
rect -5680 2501 -5674 2898
rect -5792 2489 -5674 2501
rect -5558 2898 -5440 2910
rect -5558 2501 -5552 2898
rect -5446 2501 -5440 2898
rect -5558 2489 -5440 2501
rect -5324 2898 -5206 2910
rect -5324 2501 -5318 2898
rect -5212 2501 -5206 2898
rect -5324 2489 -5206 2501
rect -5090 2898 -4972 2910
rect -5090 2501 -5084 2898
rect -4978 2501 -4972 2898
rect -5090 2489 -4972 2501
rect -4856 2898 -4738 2910
rect -4856 2501 -4850 2898
rect -4744 2501 -4738 2898
rect -4856 2489 -4738 2501
rect -4622 2898 -4504 2910
rect -4622 2501 -4616 2898
rect -4510 2501 -4504 2898
rect -4622 2489 -4504 2501
rect -4388 2898 -4270 2910
rect -4388 2501 -4382 2898
rect -4276 2501 -4270 2898
rect -4388 2489 -4270 2501
rect -4154 2898 -4036 2910
rect -4154 2501 -4148 2898
rect -4042 2501 -4036 2898
rect -4154 2489 -4036 2501
rect -3920 2898 -3802 2910
rect -3920 2501 -3914 2898
rect -3808 2501 -3802 2898
rect -3920 2489 -3802 2501
rect -3686 2898 -3568 2910
rect -3686 2501 -3680 2898
rect -3574 2501 -3568 2898
rect -3686 2489 -3568 2501
rect -3452 2898 -3334 2910
rect -3452 2501 -3446 2898
rect -3340 2501 -3334 2898
rect -3452 2489 -3334 2501
rect -3218 2898 -3100 2910
rect -3218 2501 -3212 2898
rect -3106 2501 -3100 2898
rect -3218 2489 -3100 2501
rect -2984 2898 -2866 2910
rect -2984 2501 -2978 2898
rect -2872 2501 -2866 2898
rect -2984 2489 -2866 2501
rect -2750 2898 -2632 2910
rect -2750 2501 -2744 2898
rect -2638 2501 -2632 2898
rect -2750 2489 -2632 2501
rect -2516 2898 -2398 2910
rect -2516 2501 -2510 2898
rect -2404 2501 -2398 2898
rect -2516 2489 -2398 2501
rect -2282 2898 -2164 2910
rect -2282 2501 -2276 2898
rect -2170 2501 -2164 2898
rect -2282 2489 -2164 2501
rect -2048 2898 -1930 2910
rect -2048 2501 -2042 2898
rect -1936 2501 -1930 2898
rect -2048 2489 -1930 2501
rect -1814 2898 -1696 2910
rect -1814 2501 -1808 2898
rect -1702 2501 -1696 2898
rect -1814 2489 -1696 2501
rect -1580 2898 -1462 2910
rect -1580 2501 -1574 2898
rect -1468 2501 -1462 2898
rect -1580 2489 -1462 2501
rect -1346 2898 -1228 2910
rect -1346 2501 -1340 2898
rect -1234 2501 -1228 2898
rect -1346 2489 -1228 2501
rect -1112 2898 -994 2910
rect -1112 2501 -1106 2898
rect -1000 2501 -994 2898
rect -1112 2489 -994 2501
rect -878 2898 -760 2910
rect -878 2501 -872 2898
rect -766 2501 -760 2898
rect -878 2489 -760 2501
rect -644 2898 -526 2910
rect -644 2501 -638 2898
rect -532 2501 -526 2898
rect -644 2489 -526 2501
rect -410 2898 -292 2910
rect -410 2501 -404 2898
rect -298 2501 -292 2898
rect -410 2489 -292 2501
rect -176 2898 -58 2910
rect -176 2501 -170 2898
rect -64 2501 -58 2898
rect -176 2489 -58 2501
rect 58 2898 176 2910
rect 58 2501 64 2898
rect 170 2501 176 2898
rect 58 2489 176 2501
rect 292 2898 410 2910
rect 292 2501 298 2898
rect 404 2501 410 2898
rect 292 2489 410 2501
rect 526 2898 644 2910
rect 526 2501 532 2898
rect 638 2501 644 2898
rect 526 2489 644 2501
rect 760 2898 878 2910
rect 760 2501 766 2898
rect 872 2501 878 2898
rect 760 2489 878 2501
rect 994 2898 1112 2910
rect 994 2501 1000 2898
rect 1106 2501 1112 2898
rect 994 2489 1112 2501
rect 1228 2898 1346 2910
rect 1228 2501 1234 2898
rect 1340 2501 1346 2898
rect 1228 2489 1346 2501
rect 1462 2898 1580 2910
rect 1462 2501 1468 2898
rect 1574 2501 1580 2898
rect 1462 2489 1580 2501
rect 1696 2898 1814 2910
rect 1696 2501 1702 2898
rect 1808 2501 1814 2898
rect 1696 2489 1814 2501
rect 1930 2898 2048 2910
rect 1930 2501 1936 2898
rect 2042 2501 2048 2898
rect 1930 2489 2048 2501
rect 2164 2898 2282 2910
rect 2164 2501 2170 2898
rect 2276 2501 2282 2898
rect 2164 2489 2282 2501
rect 2398 2898 2516 2910
rect 2398 2501 2404 2898
rect 2510 2501 2516 2898
rect 2398 2489 2516 2501
rect 2632 2898 2750 2910
rect 2632 2501 2638 2898
rect 2744 2501 2750 2898
rect 2632 2489 2750 2501
rect 2866 2898 2984 2910
rect 2866 2501 2872 2898
rect 2978 2501 2984 2898
rect 2866 2489 2984 2501
rect 3100 2898 3218 2910
rect 3100 2501 3106 2898
rect 3212 2501 3218 2898
rect 3100 2489 3218 2501
rect 3334 2898 3452 2910
rect 3334 2501 3340 2898
rect 3446 2501 3452 2898
rect 3334 2489 3452 2501
rect 3568 2898 3686 2910
rect 3568 2501 3574 2898
rect 3680 2501 3686 2898
rect 3568 2489 3686 2501
rect 3802 2898 3920 2910
rect 3802 2501 3808 2898
rect 3914 2501 3920 2898
rect 3802 2489 3920 2501
rect 4036 2898 4154 2910
rect 4036 2501 4042 2898
rect 4148 2501 4154 2898
rect 4036 2489 4154 2501
rect 4270 2898 4388 2910
rect 4270 2501 4276 2898
rect 4382 2501 4388 2898
rect 4270 2489 4388 2501
rect 4504 2898 4622 2910
rect 4504 2501 4510 2898
rect 4616 2501 4622 2898
rect 4504 2489 4622 2501
rect 4738 2898 4856 2910
rect 4738 2501 4744 2898
rect 4850 2501 4856 2898
rect 4738 2489 4856 2501
rect 4972 2898 5090 2910
rect 4972 2501 4978 2898
rect 5084 2501 5090 2898
rect 4972 2489 5090 2501
rect 5206 2898 5324 2910
rect 5206 2501 5212 2898
rect 5318 2501 5324 2898
rect 5206 2489 5324 2501
rect 5440 2898 5558 2910
rect 5440 2501 5446 2898
rect 5552 2501 5558 2898
rect 5440 2489 5558 2501
rect 5674 2898 5792 2910
rect 5674 2501 5680 2898
rect 5786 2501 5792 2898
rect 5674 2489 5792 2501
rect 5908 2898 6026 2910
rect 5908 2501 5914 2898
rect 6020 2501 6026 2898
rect 5908 2489 6026 2501
rect 6142 2898 6260 2910
rect 6142 2501 6148 2898
rect 6254 2501 6260 2898
rect 6142 2489 6260 2501
rect 6376 2898 6494 2910
rect 6376 2501 6382 2898
rect 6488 2501 6494 2898
rect 6376 2489 6494 2501
rect 6610 2898 6728 2910
rect 6610 2501 6616 2898
rect 6722 2501 6728 2898
rect 6610 2489 6728 2501
rect 6844 2898 6962 2910
rect 6844 2501 6850 2898
rect 6956 2501 6962 2898
rect 6844 2489 6962 2501
rect 7078 2898 7196 2910
rect 7078 2501 7084 2898
rect 7190 2501 7196 2898
rect 7078 2489 7196 2501
rect 7312 2898 7430 2910
rect 7312 2501 7318 2898
rect 7424 2501 7430 2898
rect 7312 2489 7430 2501
rect 7546 2898 7664 2910
rect 7546 2501 7552 2898
rect 7658 2501 7664 2898
rect 7546 2489 7664 2501
rect 7780 2898 7898 2910
rect 7780 2501 7786 2898
rect 7892 2501 7898 2898
rect 7780 2489 7898 2501
rect 8014 2898 8132 2910
rect 8014 2501 8020 2898
rect 8126 2501 8132 2898
rect 8014 2489 8132 2501
rect 8248 2898 8366 2910
rect 8248 2501 8254 2898
rect 8360 2501 8366 2898
rect 8248 2489 8366 2501
rect 8482 2898 8600 2910
rect 8482 2501 8488 2898
rect 8594 2501 8600 2898
rect 8482 2489 8600 2501
rect 8716 2898 8834 2910
rect 8716 2501 8722 2898
rect 8828 2501 8834 2898
rect 8716 2489 8834 2501
rect 8950 2898 9068 2910
rect 8950 2501 8956 2898
rect 9062 2501 9068 2898
rect 8950 2489 9068 2501
rect 9184 2898 9302 2910
rect 9184 2501 9190 2898
rect 9296 2501 9302 2898
rect 9184 2489 9302 2501
rect 9418 2898 9536 2910
rect 9418 2501 9424 2898
rect 9530 2501 9536 2898
rect 9418 2489 9536 2501
rect 9652 2898 9770 2910
rect 9652 2501 9658 2898
rect 9764 2501 9770 2898
rect 9652 2489 9770 2501
rect 9886 2898 10004 2910
rect 9886 2501 9892 2898
rect 9998 2501 10004 2898
rect 9886 2489 10004 2501
rect 10120 2898 10238 2910
rect 10120 2501 10126 2898
rect 10232 2501 10238 2898
rect 10120 2489 10238 2501
rect 10354 2898 10472 2910
rect 10354 2501 10360 2898
rect 10466 2501 10472 2898
rect 10354 2489 10472 2501
rect 10588 2898 10706 2910
rect 10588 2501 10594 2898
rect 10700 2501 10706 2898
rect 10588 2489 10706 2501
rect 10822 2898 10940 2910
rect 10822 2501 10828 2898
rect 10934 2501 10940 2898
rect 10822 2489 10940 2501
rect 11056 2898 11174 2910
rect 11056 2501 11062 2898
rect 11168 2501 11174 2898
rect 11056 2489 11174 2501
rect 11290 2898 11408 2910
rect 11290 2501 11296 2898
rect 11402 2501 11408 2898
rect 11290 2489 11408 2501
rect 11524 2898 11642 2910
rect 11524 2501 11530 2898
rect 11636 2501 11642 2898
rect 11524 2489 11642 2501
rect 11758 2898 11876 2910
rect 11758 2501 11764 2898
rect 11870 2501 11876 2898
rect 11758 2489 11876 2501
rect 11992 2898 12110 2910
rect 11992 2501 11998 2898
rect 12104 2501 12110 2898
rect 11992 2489 12110 2501
rect 12226 2898 12344 2910
rect 12226 2501 12232 2898
rect 12338 2501 12344 2898
rect 12226 2489 12344 2501
rect 12460 2898 12578 2910
rect 12460 2501 12466 2898
rect 12572 2501 12578 2898
rect 12460 2489 12578 2501
rect 12694 2898 12812 2910
rect 12694 2501 12700 2898
rect 12806 2501 12812 2898
rect 12694 2489 12812 2501
rect 12928 2898 13046 2910
rect 12928 2501 12934 2898
rect 13040 2501 13046 2898
rect 12928 2489 13046 2501
rect 13162 2898 13280 2910
rect 13162 2501 13168 2898
rect 13274 2501 13280 2898
rect 13162 2489 13280 2501
rect 13396 2898 13514 2910
rect 13396 2501 13402 2898
rect 13508 2501 13514 2898
rect 13396 2489 13514 2501
rect 13630 2898 13748 2910
rect 13630 2501 13636 2898
rect 13742 2501 13748 2898
rect 13630 2489 13748 2501
rect 13864 2898 13982 2910
rect 13864 2501 13870 2898
rect 13976 2501 13982 2898
rect 13864 2489 13982 2501
rect 14098 2898 14216 2910
rect 14098 2501 14104 2898
rect 14210 2501 14216 2898
rect 14098 2489 14216 2501
rect 14332 2898 14450 2910
rect 14332 2501 14338 2898
rect 14444 2501 14450 2898
rect 14332 2489 14450 2501
rect 14566 2898 14684 2910
rect 14566 2501 14572 2898
rect 14678 2501 14684 2898
rect 14566 2489 14684 2501
rect 14800 2898 14918 2910
rect 14800 2501 14806 2898
rect 14912 2501 14918 2898
rect 14800 2489 14918 2501
rect 15034 2898 15152 2910
rect 15034 2501 15040 2898
rect 15146 2501 15152 2898
rect 15034 2489 15152 2501
rect 15268 2898 15386 2910
rect 15268 2501 15274 2898
rect 15380 2501 15386 2898
rect 15268 2489 15386 2501
rect 15502 2898 15620 2910
rect 15502 2501 15508 2898
rect 15614 2501 15620 2898
rect 15502 2489 15620 2501
rect 15736 2898 15854 2910
rect 15736 2501 15742 2898
rect 15848 2501 15854 2898
rect 15736 2489 15854 2501
rect 15970 2898 16088 2910
rect 15970 2501 15976 2898
rect 16082 2501 16088 2898
rect 15970 2489 16088 2501
rect 16204 2898 16322 2910
rect 16204 2501 16210 2898
rect 16316 2501 16322 2898
rect 16204 2489 16322 2501
rect 16438 2898 16556 2910
rect 16438 2501 16444 2898
rect 16550 2501 16556 2898
rect 16438 2489 16556 2501
rect 16672 2898 16790 2910
rect 16672 2501 16678 2898
rect 16784 2501 16790 2898
rect 16672 2489 16790 2501
rect 16906 2898 17024 2910
rect 16906 2501 16912 2898
rect 17018 2501 17024 2898
rect 16906 2489 17024 2501
rect 17140 2898 17258 2910
rect 17140 2501 17146 2898
rect 17252 2501 17258 2898
rect 17140 2489 17258 2501
rect 17374 2898 17492 2910
rect 17374 2501 17380 2898
rect 17486 2501 17492 2898
rect 17374 2489 17492 2501
rect 17608 2898 17726 2910
rect 17608 2501 17614 2898
rect 17720 2501 17726 2898
rect 17608 2489 17726 2501
rect 17842 2898 17960 2910
rect 17842 2501 17848 2898
rect 17954 2501 17960 2898
rect 17842 2489 17960 2501
rect 18076 2898 18194 2910
rect 18076 2501 18082 2898
rect 18188 2501 18194 2898
rect 18076 2489 18194 2501
rect 18310 2898 18428 2910
rect 18310 2501 18316 2898
rect 18422 2501 18428 2898
rect 18310 2489 18428 2501
rect 18544 2898 18662 2910
rect 18544 2501 18550 2898
rect 18656 2501 18662 2898
rect 18544 2489 18662 2501
rect 18778 2898 18896 2910
rect 18778 2501 18784 2898
rect 18890 2501 18896 2898
rect 18778 2489 18896 2501
rect 19012 2898 19130 2910
rect 19012 2501 19018 2898
rect 19124 2501 19130 2898
rect 19012 2489 19130 2501
rect 19246 2898 19364 2910
rect 19246 2501 19252 2898
rect 19358 2501 19364 2898
rect 19246 2489 19364 2501
rect 19480 2898 19598 2910
rect 19480 2501 19486 2898
rect 19592 2501 19598 2898
rect 19480 2489 19598 2501
rect 19714 2898 19832 2910
rect 19714 2501 19720 2898
rect 19826 2501 19832 2898
rect 19714 2489 19832 2501
rect 19948 2898 20066 2910
rect 19948 2501 19954 2898
rect 20060 2501 20066 2898
rect 19948 2489 20066 2501
rect 20182 2898 20300 2910
rect 20182 2501 20188 2898
rect 20294 2501 20300 2898
rect 20182 2489 20300 2501
rect 20416 2898 20534 2910
rect 20416 2501 20422 2898
rect 20528 2501 20534 2898
rect 20416 2489 20534 2501
rect 20650 2898 20768 2910
rect 20650 2501 20656 2898
rect 20762 2501 20768 2898
rect 20650 2489 20768 2501
rect 20884 2898 21002 2910
rect 20884 2501 20890 2898
rect 20996 2501 21002 2898
rect 20884 2489 21002 2501
rect 21118 2898 21236 2910
rect 21118 2501 21124 2898
rect 21230 2501 21236 2898
rect 21118 2489 21236 2501
rect 21352 2898 21470 2910
rect 21352 2501 21358 2898
rect 21464 2501 21470 2898
rect 21352 2489 21470 2501
rect 21586 2898 21704 2910
rect 21586 2501 21592 2898
rect 21698 2501 21704 2898
rect 21586 2489 21704 2501
rect 21820 2898 21938 2910
rect 21820 2501 21826 2898
rect 21932 2501 21938 2898
rect 21820 2489 21938 2501
rect 22054 2898 22172 2910
rect 22054 2501 22060 2898
rect 22166 2501 22172 2898
rect 22054 2489 22172 2501
rect 22288 2898 22406 2910
rect 22288 2501 22294 2898
rect 22400 2501 22406 2898
rect 22288 2489 22406 2501
rect 22522 2898 22640 2910
rect 22522 2501 22528 2898
rect 22634 2501 22640 2898
rect 22522 2489 22640 2501
rect 22756 2898 22874 2910
rect 22756 2501 22762 2898
rect 22868 2501 22874 2898
rect 22756 2489 22874 2501
rect 22990 2898 23108 2910
rect 22990 2501 22996 2898
rect 23102 2501 23108 2898
rect 22990 2489 23108 2501
rect 23224 2898 23342 2910
rect 23224 2501 23230 2898
rect 23336 2501 23342 2898
rect 23224 2489 23342 2501
rect 23458 2898 23576 2910
rect 23458 2501 23464 2898
rect 23570 2501 23576 2898
rect 23458 2489 23576 2501
rect 23692 2898 23810 2910
rect 23692 2501 23698 2898
rect 23804 2501 23810 2898
rect 23692 2489 23810 2501
rect 23926 2898 24044 2910
rect 23926 2501 23932 2898
rect 24038 2501 24044 2898
rect 23926 2489 24044 2501
rect 24160 2898 24278 2910
rect 24160 2501 24166 2898
rect 24272 2501 24278 2898
rect 24160 2489 24278 2501
rect 24394 2898 24512 2910
rect 24394 2501 24400 2898
rect 24506 2501 24512 2898
rect 24394 2489 24512 2501
rect 24628 2898 24746 2910
rect 24628 2501 24634 2898
rect 24740 2501 24746 2898
rect 24628 2489 24746 2501
rect 24862 2898 24980 2910
rect 24862 2501 24868 2898
rect 24974 2501 24980 2898
rect 24862 2489 24980 2501
rect 25096 2898 25214 2910
rect 25096 2501 25102 2898
rect 25208 2501 25214 2898
rect 25096 2489 25214 2501
rect 25330 2898 25448 2910
rect 25330 2501 25336 2898
rect 25442 2501 25448 2898
rect 25330 2489 25448 2501
rect 25564 2898 25682 2910
rect 25564 2501 25570 2898
rect 25676 2501 25682 2898
rect 25564 2489 25682 2501
rect 25798 2898 25916 2910
rect 25798 2501 25804 2898
rect 25910 2501 25916 2898
rect 25798 2489 25916 2501
rect 26032 2898 26150 2910
rect 26032 2501 26038 2898
rect 26144 2501 26150 2898
rect 26032 2489 26150 2501
rect 26266 2898 26384 2910
rect 26266 2501 26272 2898
rect 26378 2501 26384 2898
rect 26266 2489 26384 2501
rect 26500 2898 26618 2910
rect 26500 2501 26506 2898
rect 26612 2501 26618 2898
rect 26500 2489 26618 2501
rect 26734 2898 26852 2910
rect 26734 2501 26740 2898
rect 26846 2501 26852 2898
rect 26734 2489 26852 2501
rect 26968 2898 27086 2910
rect 26968 2501 26974 2898
rect 27080 2501 27086 2898
rect 26968 2489 27086 2501
rect 27202 2898 27320 2910
rect 27202 2501 27208 2898
rect 27314 2501 27320 2898
rect 27202 2489 27320 2501
rect 27436 2898 27554 2910
rect 27436 2501 27442 2898
rect 27548 2501 27554 2898
rect 27436 2489 27554 2501
rect 27670 2898 27788 2910
rect 27670 2501 27676 2898
rect 27782 2501 27788 2898
rect 27670 2489 27788 2501
rect 27904 2898 28022 2910
rect 27904 2501 27910 2898
rect 28016 2501 28022 2898
rect 27904 2489 28022 2501
rect 28138 2898 28256 2910
rect 28138 2501 28144 2898
rect 28250 2501 28256 2898
rect 28138 2489 28256 2501
rect 28372 2898 28490 2910
rect 28372 2501 28378 2898
rect 28484 2501 28490 2898
rect 28372 2489 28490 2501
rect 28606 2898 28724 2910
rect 28606 2501 28612 2898
rect 28718 2501 28724 2898
rect 28606 2489 28724 2501
rect 28840 2898 28958 2910
rect 28840 2501 28846 2898
rect 28952 2501 28958 2898
rect 28840 2489 28958 2501
rect 29074 2898 29192 2910
rect 29074 2501 29080 2898
rect 29186 2501 29192 2898
rect 29074 2489 29192 2501
rect 29308 2898 29426 2910
rect 29308 2501 29314 2898
rect 29420 2501 29426 2898
rect 29308 2489 29426 2501
rect 29542 2898 29660 2910
rect 29542 2501 29548 2898
rect 29654 2501 29660 2898
rect 29542 2489 29660 2501
rect 29776 2898 29894 2910
rect 29776 2501 29782 2898
rect 29888 2501 29894 2898
rect 29776 2489 29894 2501
rect -29894 -2501 -29776 -2489
rect -29894 -2898 -29888 -2501
rect -29782 -2898 -29776 -2501
rect -29894 -2910 -29776 -2898
rect -29660 -2501 -29542 -2489
rect -29660 -2898 -29654 -2501
rect -29548 -2898 -29542 -2501
rect -29660 -2910 -29542 -2898
rect -29426 -2501 -29308 -2489
rect -29426 -2898 -29420 -2501
rect -29314 -2898 -29308 -2501
rect -29426 -2910 -29308 -2898
rect -29192 -2501 -29074 -2489
rect -29192 -2898 -29186 -2501
rect -29080 -2898 -29074 -2501
rect -29192 -2910 -29074 -2898
rect -28958 -2501 -28840 -2489
rect -28958 -2898 -28952 -2501
rect -28846 -2898 -28840 -2501
rect -28958 -2910 -28840 -2898
rect -28724 -2501 -28606 -2489
rect -28724 -2898 -28718 -2501
rect -28612 -2898 -28606 -2501
rect -28724 -2910 -28606 -2898
rect -28490 -2501 -28372 -2489
rect -28490 -2898 -28484 -2501
rect -28378 -2898 -28372 -2501
rect -28490 -2910 -28372 -2898
rect -28256 -2501 -28138 -2489
rect -28256 -2898 -28250 -2501
rect -28144 -2898 -28138 -2501
rect -28256 -2910 -28138 -2898
rect -28022 -2501 -27904 -2489
rect -28022 -2898 -28016 -2501
rect -27910 -2898 -27904 -2501
rect -28022 -2910 -27904 -2898
rect -27788 -2501 -27670 -2489
rect -27788 -2898 -27782 -2501
rect -27676 -2898 -27670 -2501
rect -27788 -2910 -27670 -2898
rect -27554 -2501 -27436 -2489
rect -27554 -2898 -27548 -2501
rect -27442 -2898 -27436 -2501
rect -27554 -2910 -27436 -2898
rect -27320 -2501 -27202 -2489
rect -27320 -2898 -27314 -2501
rect -27208 -2898 -27202 -2501
rect -27320 -2910 -27202 -2898
rect -27086 -2501 -26968 -2489
rect -27086 -2898 -27080 -2501
rect -26974 -2898 -26968 -2501
rect -27086 -2910 -26968 -2898
rect -26852 -2501 -26734 -2489
rect -26852 -2898 -26846 -2501
rect -26740 -2898 -26734 -2501
rect -26852 -2910 -26734 -2898
rect -26618 -2501 -26500 -2489
rect -26618 -2898 -26612 -2501
rect -26506 -2898 -26500 -2501
rect -26618 -2910 -26500 -2898
rect -26384 -2501 -26266 -2489
rect -26384 -2898 -26378 -2501
rect -26272 -2898 -26266 -2501
rect -26384 -2910 -26266 -2898
rect -26150 -2501 -26032 -2489
rect -26150 -2898 -26144 -2501
rect -26038 -2898 -26032 -2501
rect -26150 -2910 -26032 -2898
rect -25916 -2501 -25798 -2489
rect -25916 -2898 -25910 -2501
rect -25804 -2898 -25798 -2501
rect -25916 -2910 -25798 -2898
rect -25682 -2501 -25564 -2489
rect -25682 -2898 -25676 -2501
rect -25570 -2898 -25564 -2501
rect -25682 -2910 -25564 -2898
rect -25448 -2501 -25330 -2489
rect -25448 -2898 -25442 -2501
rect -25336 -2898 -25330 -2501
rect -25448 -2910 -25330 -2898
rect -25214 -2501 -25096 -2489
rect -25214 -2898 -25208 -2501
rect -25102 -2898 -25096 -2501
rect -25214 -2910 -25096 -2898
rect -24980 -2501 -24862 -2489
rect -24980 -2898 -24974 -2501
rect -24868 -2898 -24862 -2501
rect -24980 -2910 -24862 -2898
rect -24746 -2501 -24628 -2489
rect -24746 -2898 -24740 -2501
rect -24634 -2898 -24628 -2501
rect -24746 -2910 -24628 -2898
rect -24512 -2501 -24394 -2489
rect -24512 -2898 -24506 -2501
rect -24400 -2898 -24394 -2501
rect -24512 -2910 -24394 -2898
rect -24278 -2501 -24160 -2489
rect -24278 -2898 -24272 -2501
rect -24166 -2898 -24160 -2501
rect -24278 -2910 -24160 -2898
rect -24044 -2501 -23926 -2489
rect -24044 -2898 -24038 -2501
rect -23932 -2898 -23926 -2501
rect -24044 -2910 -23926 -2898
rect -23810 -2501 -23692 -2489
rect -23810 -2898 -23804 -2501
rect -23698 -2898 -23692 -2501
rect -23810 -2910 -23692 -2898
rect -23576 -2501 -23458 -2489
rect -23576 -2898 -23570 -2501
rect -23464 -2898 -23458 -2501
rect -23576 -2910 -23458 -2898
rect -23342 -2501 -23224 -2489
rect -23342 -2898 -23336 -2501
rect -23230 -2898 -23224 -2501
rect -23342 -2910 -23224 -2898
rect -23108 -2501 -22990 -2489
rect -23108 -2898 -23102 -2501
rect -22996 -2898 -22990 -2501
rect -23108 -2910 -22990 -2898
rect -22874 -2501 -22756 -2489
rect -22874 -2898 -22868 -2501
rect -22762 -2898 -22756 -2501
rect -22874 -2910 -22756 -2898
rect -22640 -2501 -22522 -2489
rect -22640 -2898 -22634 -2501
rect -22528 -2898 -22522 -2501
rect -22640 -2910 -22522 -2898
rect -22406 -2501 -22288 -2489
rect -22406 -2898 -22400 -2501
rect -22294 -2898 -22288 -2501
rect -22406 -2910 -22288 -2898
rect -22172 -2501 -22054 -2489
rect -22172 -2898 -22166 -2501
rect -22060 -2898 -22054 -2501
rect -22172 -2910 -22054 -2898
rect -21938 -2501 -21820 -2489
rect -21938 -2898 -21932 -2501
rect -21826 -2898 -21820 -2501
rect -21938 -2910 -21820 -2898
rect -21704 -2501 -21586 -2489
rect -21704 -2898 -21698 -2501
rect -21592 -2898 -21586 -2501
rect -21704 -2910 -21586 -2898
rect -21470 -2501 -21352 -2489
rect -21470 -2898 -21464 -2501
rect -21358 -2898 -21352 -2501
rect -21470 -2910 -21352 -2898
rect -21236 -2501 -21118 -2489
rect -21236 -2898 -21230 -2501
rect -21124 -2898 -21118 -2501
rect -21236 -2910 -21118 -2898
rect -21002 -2501 -20884 -2489
rect -21002 -2898 -20996 -2501
rect -20890 -2898 -20884 -2501
rect -21002 -2910 -20884 -2898
rect -20768 -2501 -20650 -2489
rect -20768 -2898 -20762 -2501
rect -20656 -2898 -20650 -2501
rect -20768 -2910 -20650 -2898
rect -20534 -2501 -20416 -2489
rect -20534 -2898 -20528 -2501
rect -20422 -2898 -20416 -2501
rect -20534 -2910 -20416 -2898
rect -20300 -2501 -20182 -2489
rect -20300 -2898 -20294 -2501
rect -20188 -2898 -20182 -2501
rect -20300 -2910 -20182 -2898
rect -20066 -2501 -19948 -2489
rect -20066 -2898 -20060 -2501
rect -19954 -2898 -19948 -2501
rect -20066 -2910 -19948 -2898
rect -19832 -2501 -19714 -2489
rect -19832 -2898 -19826 -2501
rect -19720 -2898 -19714 -2501
rect -19832 -2910 -19714 -2898
rect -19598 -2501 -19480 -2489
rect -19598 -2898 -19592 -2501
rect -19486 -2898 -19480 -2501
rect -19598 -2910 -19480 -2898
rect -19364 -2501 -19246 -2489
rect -19364 -2898 -19358 -2501
rect -19252 -2898 -19246 -2501
rect -19364 -2910 -19246 -2898
rect -19130 -2501 -19012 -2489
rect -19130 -2898 -19124 -2501
rect -19018 -2898 -19012 -2501
rect -19130 -2910 -19012 -2898
rect -18896 -2501 -18778 -2489
rect -18896 -2898 -18890 -2501
rect -18784 -2898 -18778 -2501
rect -18896 -2910 -18778 -2898
rect -18662 -2501 -18544 -2489
rect -18662 -2898 -18656 -2501
rect -18550 -2898 -18544 -2501
rect -18662 -2910 -18544 -2898
rect -18428 -2501 -18310 -2489
rect -18428 -2898 -18422 -2501
rect -18316 -2898 -18310 -2501
rect -18428 -2910 -18310 -2898
rect -18194 -2501 -18076 -2489
rect -18194 -2898 -18188 -2501
rect -18082 -2898 -18076 -2501
rect -18194 -2910 -18076 -2898
rect -17960 -2501 -17842 -2489
rect -17960 -2898 -17954 -2501
rect -17848 -2898 -17842 -2501
rect -17960 -2910 -17842 -2898
rect -17726 -2501 -17608 -2489
rect -17726 -2898 -17720 -2501
rect -17614 -2898 -17608 -2501
rect -17726 -2910 -17608 -2898
rect -17492 -2501 -17374 -2489
rect -17492 -2898 -17486 -2501
rect -17380 -2898 -17374 -2501
rect -17492 -2910 -17374 -2898
rect -17258 -2501 -17140 -2489
rect -17258 -2898 -17252 -2501
rect -17146 -2898 -17140 -2501
rect -17258 -2910 -17140 -2898
rect -17024 -2501 -16906 -2489
rect -17024 -2898 -17018 -2501
rect -16912 -2898 -16906 -2501
rect -17024 -2910 -16906 -2898
rect -16790 -2501 -16672 -2489
rect -16790 -2898 -16784 -2501
rect -16678 -2898 -16672 -2501
rect -16790 -2910 -16672 -2898
rect -16556 -2501 -16438 -2489
rect -16556 -2898 -16550 -2501
rect -16444 -2898 -16438 -2501
rect -16556 -2910 -16438 -2898
rect -16322 -2501 -16204 -2489
rect -16322 -2898 -16316 -2501
rect -16210 -2898 -16204 -2501
rect -16322 -2910 -16204 -2898
rect -16088 -2501 -15970 -2489
rect -16088 -2898 -16082 -2501
rect -15976 -2898 -15970 -2501
rect -16088 -2910 -15970 -2898
rect -15854 -2501 -15736 -2489
rect -15854 -2898 -15848 -2501
rect -15742 -2898 -15736 -2501
rect -15854 -2910 -15736 -2898
rect -15620 -2501 -15502 -2489
rect -15620 -2898 -15614 -2501
rect -15508 -2898 -15502 -2501
rect -15620 -2910 -15502 -2898
rect -15386 -2501 -15268 -2489
rect -15386 -2898 -15380 -2501
rect -15274 -2898 -15268 -2501
rect -15386 -2910 -15268 -2898
rect -15152 -2501 -15034 -2489
rect -15152 -2898 -15146 -2501
rect -15040 -2898 -15034 -2501
rect -15152 -2910 -15034 -2898
rect -14918 -2501 -14800 -2489
rect -14918 -2898 -14912 -2501
rect -14806 -2898 -14800 -2501
rect -14918 -2910 -14800 -2898
rect -14684 -2501 -14566 -2489
rect -14684 -2898 -14678 -2501
rect -14572 -2898 -14566 -2501
rect -14684 -2910 -14566 -2898
rect -14450 -2501 -14332 -2489
rect -14450 -2898 -14444 -2501
rect -14338 -2898 -14332 -2501
rect -14450 -2910 -14332 -2898
rect -14216 -2501 -14098 -2489
rect -14216 -2898 -14210 -2501
rect -14104 -2898 -14098 -2501
rect -14216 -2910 -14098 -2898
rect -13982 -2501 -13864 -2489
rect -13982 -2898 -13976 -2501
rect -13870 -2898 -13864 -2501
rect -13982 -2910 -13864 -2898
rect -13748 -2501 -13630 -2489
rect -13748 -2898 -13742 -2501
rect -13636 -2898 -13630 -2501
rect -13748 -2910 -13630 -2898
rect -13514 -2501 -13396 -2489
rect -13514 -2898 -13508 -2501
rect -13402 -2898 -13396 -2501
rect -13514 -2910 -13396 -2898
rect -13280 -2501 -13162 -2489
rect -13280 -2898 -13274 -2501
rect -13168 -2898 -13162 -2501
rect -13280 -2910 -13162 -2898
rect -13046 -2501 -12928 -2489
rect -13046 -2898 -13040 -2501
rect -12934 -2898 -12928 -2501
rect -13046 -2910 -12928 -2898
rect -12812 -2501 -12694 -2489
rect -12812 -2898 -12806 -2501
rect -12700 -2898 -12694 -2501
rect -12812 -2910 -12694 -2898
rect -12578 -2501 -12460 -2489
rect -12578 -2898 -12572 -2501
rect -12466 -2898 -12460 -2501
rect -12578 -2910 -12460 -2898
rect -12344 -2501 -12226 -2489
rect -12344 -2898 -12338 -2501
rect -12232 -2898 -12226 -2501
rect -12344 -2910 -12226 -2898
rect -12110 -2501 -11992 -2489
rect -12110 -2898 -12104 -2501
rect -11998 -2898 -11992 -2501
rect -12110 -2910 -11992 -2898
rect -11876 -2501 -11758 -2489
rect -11876 -2898 -11870 -2501
rect -11764 -2898 -11758 -2501
rect -11876 -2910 -11758 -2898
rect -11642 -2501 -11524 -2489
rect -11642 -2898 -11636 -2501
rect -11530 -2898 -11524 -2501
rect -11642 -2910 -11524 -2898
rect -11408 -2501 -11290 -2489
rect -11408 -2898 -11402 -2501
rect -11296 -2898 -11290 -2501
rect -11408 -2910 -11290 -2898
rect -11174 -2501 -11056 -2489
rect -11174 -2898 -11168 -2501
rect -11062 -2898 -11056 -2501
rect -11174 -2910 -11056 -2898
rect -10940 -2501 -10822 -2489
rect -10940 -2898 -10934 -2501
rect -10828 -2898 -10822 -2501
rect -10940 -2910 -10822 -2898
rect -10706 -2501 -10588 -2489
rect -10706 -2898 -10700 -2501
rect -10594 -2898 -10588 -2501
rect -10706 -2910 -10588 -2898
rect -10472 -2501 -10354 -2489
rect -10472 -2898 -10466 -2501
rect -10360 -2898 -10354 -2501
rect -10472 -2910 -10354 -2898
rect -10238 -2501 -10120 -2489
rect -10238 -2898 -10232 -2501
rect -10126 -2898 -10120 -2501
rect -10238 -2910 -10120 -2898
rect -10004 -2501 -9886 -2489
rect -10004 -2898 -9998 -2501
rect -9892 -2898 -9886 -2501
rect -10004 -2910 -9886 -2898
rect -9770 -2501 -9652 -2489
rect -9770 -2898 -9764 -2501
rect -9658 -2898 -9652 -2501
rect -9770 -2910 -9652 -2898
rect -9536 -2501 -9418 -2489
rect -9536 -2898 -9530 -2501
rect -9424 -2898 -9418 -2501
rect -9536 -2910 -9418 -2898
rect -9302 -2501 -9184 -2489
rect -9302 -2898 -9296 -2501
rect -9190 -2898 -9184 -2501
rect -9302 -2910 -9184 -2898
rect -9068 -2501 -8950 -2489
rect -9068 -2898 -9062 -2501
rect -8956 -2898 -8950 -2501
rect -9068 -2910 -8950 -2898
rect -8834 -2501 -8716 -2489
rect -8834 -2898 -8828 -2501
rect -8722 -2898 -8716 -2501
rect -8834 -2910 -8716 -2898
rect -8600 -2501 -8482 -2489
rect -8600 -2898 -8594 -2501
rect -8488 -2898 -8482 -2501
rect -8600 -2910 -8482 -2898
rect -8366 -2501 -8248 -2489
rect -8366 -2898 -8360 -2501
rect -8254 -2898 -8248 -2501
rect -8366 -2910 -8248 -2898
rect -8132 -2501 -8014 -2489
rect -8132 -2898 -8126 -2501
rect -8020 -2898 -8014 -2501
rect -8132 -2910 -8014 -2898
rect -7898 -2501 -7780 -2489
rect -7898 -2898 -7892 -2501
rect -7786 -2898 -7780 -2501
rect -7898 -2910 -7780 -2898
rect -7664 -2501 -7546 -2489
rect -7664 -2898 -7658 -2501
rect -7552 -2898 -7546 -2501
rect -7664 -2910 -7546 -2898
rect -7430 -2501 -7312 -2489
rect -7430 -2898 -7424 -2501
rect -7318 -2898 -7312 -2501
rect -7430 -2910 -7312 -2898
rect -7196 -2501 -7078 -2489
rect -7196 -2898 -7190 -2501
rect -7084 -2898 -7078 -2501
rect -7196 -2910 -7078 -2898
rect -6962 -2501 -6844 -2489
rect -6962 -2898 -6956 -2501
rect -6850 -2898 -6844 -2501
rect -6962 -2910 -6844 -2898
rect -6728 -2501 -6610 -2489
rect -6728 -2898 -6722 -2501
rect -6616 -2898 -6610 -2501
rect -6728 -2910 -6610 -2898
rect -6494 -2501 -6376 -2489
rect -6494 -2898 -6488 -2501
rect -6382 -2898 -6376 -2501
rect -6494 -2910 -6376 -2898
rect -6260 -2501 -6142 -2489
rect -6260 -2898 -6254 -2501
rect -6148 -2898 -6142 -2501
rect -6260 -2910 -6142 -2898
rect -6026 -2501 -5908 -2489
rect -6026 -2898 -6020 -2501
rect -5914 -2898 -5908 -2501
rect -6026 -2910 -5908 -2898
rect -5792 -2501 -5674 -2489
rect -5792 -2898 -5786 -2501
rect -5680 -2898 -5674 -2501
rect -5792 -2910 -5674 -2898
rect -5558 -2501 -5440 -2489
rect -5558 -2898 -5552 -2501
rect -5446 -2898 -5440 -2501
rect -5558 -2910 -5440 -2898
rect -5324 -2501 -5206 -2489
rect -5324 -2898 -5318 -2501
rect -5212 -2898 -5206 -2501
rect -5324 -2910 -5206 -2898
rect -5090 -2501 -4972 -2489
rect -5090 -2898 -5084 -2501
rect -4978 -2898 -4972 -2501
rect -5090 -2910 -4972 -2898
rect -4856 -2501 -4738 -2489
rect -4856 -2898 -4850 -2501
rect -4744 -2898 -4738 -2501
rect -4856 -2910 -4738 -2898
rect -4622 -2501 -4504 -2489
rect -4622 -2898 -4616 -2501
rect -4510 -2898 -4504 -2501
rect -4622 -2910 -4504 -2898
rect -4388 -2501 -4270 -2489
rect -4388 -2898 -4382 -2501
rect -4276 -2898 -4270 -2501
rect -4388 -2910 -4270 -2898
rect -4154 -2501 -4036 -2489
rect -4154 -2898 -4148 -2501
rect -4042 -2898 -4036 -2501
rect -4154 -2910 -4036 -2898
rect -3920 -2501 -3802 -2489
rect -3920 -2898 -3914 -2501
rect -3808 -2898 -3802 -2501
rect -3920 -2910 -3802 -2898
rect -3686 -2501 -3568 -2489
rect -3686 -2898 -3680 -2501
rect -3574 -2898 -3568 -2501
rect -3686 -2910 -3568 -2898
rect -3452 -2501 -3334 -2489
rect -3452 -2898 -3446 -2501
rect -3340 -2898 -3334 -2501
rect -3452 -2910 -3334 -2898
rect -3218 -2501 -3100 -2489
rect -3218 -2898 -3212 -2501
rect -3106 -2898 -3100 -2501
rect -3218 -2910 -3100 -2898
rect -2984 -2501 -2866 -2489
rect -2984 -2898 -2978 -2501
rect -2872 -2898 -2866 -2501
rect -2984 -2910 -2866 -2898
rect -2750 -2501 -2632 -2489
rect -2750 -2898 -2744 -2501
rect -2638 -2898 -2632 -2501
rect -2750 -2910 -2632 -2898
rect -2516 -2501 -2398 -2489
rect -2516 -2898 -2510 -2501
rect -2404 -2898 -2398 -2501
rect -2516 -2910 -2398 -2898
rect -2282 -2501 -2164 -2489
rect -2282 -2898 -2276 -2501
rect -2170 -2898 -2164 -2501
rect -2282 -2910 -2164 -2898
rect -2048 -2501 -1930 -2489
rect -2048 -2898 -2042 -2501
rect -1936 -2898 -1930 -2501
rect -2048 -2910 -1930 -2898
rect -1814 -2501 -1696 -2489
rect -1814 -2898 -1808 -2501
rect -1702 -2898 -1696 -2501
rect -1814 -2910 -1696 -2898
rect -1580 -2501 -1462 -2489
rect -1580 -2898 -1574 -2501
rect -1468 -2898 -1462 -2501
rect -1580 -2910 -1462 -2898
rect -1346 -2501 -1228 -2489
rect -1346 -2898 -1340 -2501
rect -1234 -2898 -1228 -2501
rect -1346 -2910 -1228 -2898
rect -1112 -2501 -994 -2489
rect -1112 -2898 -1106 -2501
rect -1000 -2898 -994 -2501
rect -1112 -2910 -994 -2898
rect -878 -2501 -760 -2489
rect -878 -2898 -872 -2501
rect -766 -2898 -760 -2501
rect -878 -2910 -760 -2898
rect -644 -2501 -526 -2489
rect -644 -2898 -638 -2501
rect -532 -2898 -526 -2501
rect -644 -2910 -526 -2898
rect -410 -2501 -292 -2489
rect -410 -2898 -404 -2501
rect -298 -2898 -292 -2501
rect -410 -2910 -292 -2898
rect -176 -2501 -58 -2489
rect -176 -2898 -170 -2501
rect -64 -2898 -58 -2501
rect -176 -2910 -58 -2898
rect 58 -2501 176 -2489
rect 58 -2898 64 -2501
rect 170 -2898 176 -2501
rect 58 -2910 176 -2898
rect 292 -2501 410 -2489
rect 292 -2898 298 -2501
rect 404 -2898 410 -2501
rect 292 -2910 410 -2898
rect 526 -2501 644 -2489
rect 526 -2898 532 -2501
rect 638 -2898 644 -2501
rect 526 -2910 644 -2898
rect 760 -2501 878 -2489
rect 760 -2898 766 -2501
rect 872 -2898 878 -2501
rect 760 -2910 878 -2898
rect 994 -2501 1112 -2489
rect 994 -2898 1000 -2501
rect 1106 -2898 1112 -2501
rect 994 -2910 1112 -2898
rect 1228 -2501 1346 -2489
rect 1228 -2898 1234 -2501
rect 1340 -2898 1346 -2501
rect 1228 -2910 1346 -2898
rect 1462 -2501 1580 -2489
rect 1462 -2898 1468 -2501
rect 1574 -2898 1580 -2501
rect 1462 -2910 1580 -2898
rect 1696 -2501 1814 -2489
rect 1696 -2898 1702 -2501
rect 1808 -2898 1814 -2501
rect 1696 -2910 1814 -2898
rect 1930 -2501 2048 -2489
rect 1930 -2898 1936 -2501
rect 2042 -2898 2048 -2501
rect 1930 -2910 2048 -2898
rect 2164 -2501 2282 -2489
rect 2164 -2898 2170 -2501
rect 2276 -2898 2282 -2501
rect 2164 -2910 2282 -2898
rect 2398 -2501 2516 -2489
rect 2398 -2898 2404 -2501
rect 2510 -2898 2516 -2501
rect 2398 -2910 2516 -2898
rect 2632 -2501 2750 -2489
rect 2632 -2898 2638 -2501
rect 2744 -2898 2750 -2501
rect 2632 -2910 2750 -2898
rect 2866 -2501 2984 -2489
rect 2866 -2898 2872 -2501
rect 2978 -2898 2984 -2501
rect 2866 -2910 2984 -2898
rect 3100 -2501 3218 -2489
rect 3100 -2898 3106 -2501
rect 3212 -2898 3218 -2501
rect 3100 -2910 3218 -2898
rect 3334 -2501 3452 -2489
rect 3334 -2898 3340 -2501
rect 3446 -2898 3452 -2501
rect 3334 -2910 3452 -2898
rect 3568 -2501 3686 -2489
rect 3568 -2898 3574 -2501
rect 3680 -2898 3686 -2501
rect 3568 -2910 3686 -2898
rect 3802 -2501 3920 -2489
rect 3802 -2898 3808 -2501
rect 3914 -2898 3920 -2501
rect 3802 -2910 3920 -2898
rect 4036 -2501 4154 -2489
rect 4036 -2898 4042 -2501
rect 4148 -2898 4154 -2501
rect 4036 -2910 4154 -2898
rect 4270 -2501 4388 -2489
rect 4270 -2898 4276 -2501
rect 4382 -2898 4388 -2501
rect 4270 -2910 4388 -2898
rect 4504 -2501 4622 -2489
rect 4504 -2898 4510 -2501
rect 4616 -2898 4622 -2501
rect 4504 -2910 4622 -2898
rect 4738 -2501 4856 -2489
rect 4738 -2898 4744 -2501
rect 4850 -2898 4856 -2501
rect 4738 -2910 4856 -2898
rect 4972 -2501 5090 -2489
rect 4972 -2898 4978 -2501
rect 5084 -2898 5090 -2501
rect 4972 -2910 5090 -2898
rect 5206 -2501 5324 -2489
rect 5206 -2898 5212 -2501
rect 5318 -2898 5324 -2501
rect 5206 -2910 5324 -2898
rect 5440 -2501 5558 -2489
rect 5440 -2898 5446 -2501
rect 5552 -2898 5558 -2501
rect 5440 -2910 5558 -2898
rect 5674 -2501 5792 -2489
rect 5674 -2898 5680 -2501
rect 5786 -2898 5792 -2501
rect 5674 -2910 5792 -2898
rect 5908 -2501 6026 -2489
rect 5908 -2898 5914 -2501
rect 6020 -2898 6026 -2501
rect 5908 -2910 6026 -2898
rect 6142 -2501 6260 -2489
rect 6142 -2898 6148 -2501
rect 6254 -2898 6260 -2501
rect 6142 -2910 6260 -2898
rect 6376 -2501 6494 -2489
rect 6376 -2898 6382 -2501
rect 6488 -2898 6494 -2501
rect 6376 -2910 6494 -2898
rect 6610 -2501 6728 -2489
rect 6610 -2898 6616 -2501
rect 6722 -2898 6728 -2501
rect 6610 -2910 6728 -2898
rect 6844 -2501 6962 -2489
rect 6844 -2898 6850 -2501
rect 6956 -2898 6962 -2501
rect 6844 -2910 6962 -2898
rect 7078 -2501 7196 -2489
rect 7078 -2898 7084 -2501
rect 7190 -2898 7196 -2501
rect 7078 -2910 7196 -2898
rect 7312 -2501 7430 -2489
rect 7312 -2898 7318 -2501
rect 7424 -2898 7430 -2501
rect 7312 -2910 7430 -2898
rect 7546 -2501 7664 -2489
rect 7546 -2898 7552 -2501
rect 7658 -2898 7664 -2501
rect 7546 -2910 7664 -2898
rect 7780 -2501 7898 -2489
rect 7780 -2898 7786 -2501
rect 7892 -2898 7898 -2501
rect 7780 -2910 7898 -2898
rect 8014 -2501 8132 -2489
rect 8014 -2898 8020 -2501
rect 8126 -2898 8132 -2501
rect 8014 -2910 8132 -2898
rect 8248 -2501 8366 -2489
rect 8248 -2898 8254 -2501
rect 8360 -2898 8366 -2501
rect 8248 -2910 8366 -2898
rect 8482 -2501 8600 -2489
rect 8482 -2898 8488 -2501
rect 8594 -2898 8600 -2501
rect 8482 -2910 8600 -2898
rect 8716 -2501 8834 -2489
rect 8716 -2898 8722 -2501
rect 8828 -2898 8834 -2501
rect 8716 -2910 8834 -2898
rect 8950 -2501 9068 -2489
rect 8950 -2898 8956 -2501
rect 9062 -2898 9068 -2501
rect 8950 -2910 9068 -2898
rect 9184 -2501 9302 -2489
rect 9184 -2898 9190 -2501
rect 9296 -2898 9302 -2501
rect 9184 -2910 9302 -2898
rect 9418 -2501 9536 -2489
rect 9418 -2898 9424 -2501
rect 9530 -2898 9536 -2501
rect 9418 -2910 9536 -2898
rect 9652 -2501 9770 -2489
rect 9652 -2898 9658 -2501
rect 9764 -2898 9770 -2501
rect 9652 -2910 9770 -2898
rect 9886 -2501 10004 -2489
rect 9886 -2898 9892 -2501
rect 9998 -2898 10004 -2501
rect 9886 -2910 10004 -2898
rect 10120 -2501 10238 -2489
rect 10120 -2898 10126 -2501
rect 10232 -2898 10238 -2501
rect 10120 -2910 10238 -2898
rect 10354 -2501 10472 -2489
rect 10354 -2898 10360 -2501
rect 10466 -2898 10472 -2501
rect 10354 -2910 10472 -2898
rect 10588 -2501 10706 -2489
rect 10588 -2898 10594 -2501
rect 10700 -2898 10706 -2501
rect 10588 -2910 10706 -2898
rect 10822 -2501 10940 -2489
rect 10822 -2898 10828 -2501
rect 10934 -2898 10940 -2501
rect 10822 -2910 10940 -2898
rect 11056 -2501 11174 -2489
rect 11056 -2898 11062 -2501
rect 11168 -2898 11174 -2501
rect 11056 -2910 11174 -2898
rect 11290 -2501 11408 -2489
rect 11290 -2898 11296 -2501
rect 11402 -2898 11408 -2501
rect 11290 -2910 11408 -2898
rect 11524 -2501 11642 -2489
rect 11524 -2898 11530 -2501
rect 11636 -2898 11642 -2501
rect 11524 -2910 11642 -2898
rect 11758 -2501 11876 -2489
rect 11758 -2898 11764 -2501
rect 11870 -2898 11876 -2501
rect 11758 -2910 11876 -2898
rect 11992 -2501 12110 -2489
rect 11992 -2898 11998 -2501
rect 12104 -2898 12110 -2501
rect 11992 -2910 12110 -2898
rect 12226 -2501 12344 -2489
rect 12226 -2898 12232 -2501
rect 12338 -2898 12344 -2501
rect 12226 -2910 12344 -2898
rect 12460 -2501 12578 -2489
rect 12460 -2898 12466 -2501
rect 12572 -2898 12578 -2501
rect 12460 -2910 12578 -2898
rect 12694 -2501 12812 -2489
rect 12694 -2898 12700 -2501
rect 12806 -2898 12812 -2501
rect 12694 -2910 12812 -2898
rect 12928 -2501 13046 -2489
rect 12928 -2898 12934 -2501
rect 13040 -2898 13046 -2501
rect 12928 -2910 13046 -2898
rect 13162 -2501 13280 -2489
rect 13162 -2898 13168 -2501
rect 13274 -2898 13280 -2501
rect 13162 -2910 13280 -2898
rect 13396 -2501 13514 -2489
rect 13396 -2898 13402 -2501
rect 13508 -2898 13514 -2501
rect 13396 -2910 13514 -2898
rect 13630 -2501 13748 -2489
rect 13630 -2898 13636 -2501
rect 13742 -2898 13748 -2501
rect 13630 -2910 13748 -2898
rect 13864 -2501 13982 -2489
rect 13864 -2898 13870 -2501
rect 13976 -2898 13982 -2501
rect 13864 -2910 13982 -2898
rect 14098 -2501 14216 -2489
rect 14098 -2898 14104 -2501
rect 14210 -2898 14216 -2501
rect 14098 -2910 14216 -2898
rect 14332 -2501 14450 -2489
rect 14332 -2898 14338 -2501
rect 14444 -2898 14450 -2501
rect 14332 -2910 14450 -2898
rect 14566 -2501 14684 -2489
rect 14566 -2898 14572 -2501
rect 14678 -2898 14684 -2501
rect 14566 -2910 14684 -2898
rect 14800 -2501 14918 -2489
rect 14800 -2898 14806 -2501
rect 14912 -2898 14918 -2501
rect 14800 -2910 14918 -2898
rect 15034 -2501 15152 -2489
rect 15034 -2898 15040 -2501
rect 15146 -2898 15152 -2501
rect 15034 -2910 15152 -2898
rect 15268 -2501 15386 -2489
rect 15268 -2898 15274 -2501
rect 15380 -2898 15386 -2501
rect 15268 -2910 15386 -2898
rect 15502 -2501 15620 -2489
rect 15502 -2898 15508 -2501
rect 15614 -2898 15620 -2501
rect 15502 -2910 15620 -2898
rect 15736 -2501 15854 -2489
rect 15736 -2898 15742 -2501
rect 15848 -2898 15854 -2501
rect 15736 -2910 15854 -2898
rect 15970 -2501 16088 -2489
rect 15970 -2898 15976 -2501
rect 16082 -2898 16088 -2501
rect 15970 -2910 16088 -2898
rect 16204 -2501 16322 -2489
rect 16204 -2898 16210 -2501
rect 16316 -2898 16322 -2501
rect 16204 -2910 16322 -2898
rect 16438 -2501 16556 -2489
rect 16438 -2898 16444 -2501
rect 16550 -2898 16556 -2501
rect 16438 -2910 16556 -2898
rect 16672 -2501 16790 -2489
rect 16672 -2898 16678 -2501
rect 16784 -2898 16790 -2501
rect 16672 -2910 16790 -2898
rect 16906 -2501 17024 -2489
rect 16906 -2898 16912 -2501
rect 17018 -2898 17024 -2501
rect 16906 -2910 17024 -2898
rect 17140 -2501 17258 -2489
rect 17140 -2898 17146 -2501
rect 17252 -2898 17258 -2501
rect 17140 -2910 17258 -2898
rect 17374 -2501 17492 -2489
rect 17374 -2898 17380 -2501
rect 17486 -2898 17492 -2501
rect 17374 -2910 17492 -2898
rect 17608 -2501 17726 -2489
rect 17608 -2898 17614 -2501
rect 17720 -2898 17726 -2501
rect 17608 -2910 17726 -2898
rect 17842 -2501 17960 -2489
rect 17842 -2898 17848 -2501
rect 17954 -2898 17960 -2501
rect 17842 -2910 17960 -2898
rect 18076 -2501 18194 -2489
rect 18076 -2898 18082 -2501
rect 18188 -2898 18194 -2501
rect 18076 -2910 18194 -2898
rect 18310 -2501 18428 -2489
rect 18310 -2898 18316 -2501
rect 18422 -2898 18428 -2501
rect 18310 -2910 18428 -2898
rect 18544 -2501 18662 -2489
rect 18544 -2898 18550 -2501
rect 18656 -2898 18662 -2501
rect 18544 -2910 18662 -2898
rect 18778 -2501 18896 -2489
rect 18778 -2898 18784 -2501
rect 18890 -2898 18896 -2501
rect 18778 -2910 18896 -2898
rect 19012 -2501 19130 -2489
rect 19012 -2898 19018 -2501
rect 19124 -2898 19130 -2501
rect 19012 -2910 19130 -2898
rect 19246 -2501 19364 -2489
rect 19246 -2898 19252 -2501
rect 19358 -2898 19364 -2501
rect 19246 -2910 19364 -2898
rect 19480 -2501 19598 -2489
rect 19480 -2898 19486 -2501
rect 19592 -2898 19598 -2501
rect 19480 -2910 19598 -2898
rect 19714 -2501 19832 -2489
rect 19714 -2898 19720 -2501
rect 19826 -2898 19832 -2501
rect 19714 -2910 19832 -2898
rect 19948 -2501 20066 -2489
rect 19948 -2898 19954 -2501
rect 20060 -2898 20066 -2501
rect 19948 -2910 20066 -2898
rect 20182 -2501 20300 -2489
rect 20182 -2898 20188 -2501
rect 20294 -2898 20300 -2501
rect 20182 -2910 20300 -2898
rect 20416 -2501 20534 -2489
rect 20416 -2898 20422 -2501
rect 20528 -2898 20534 -2501
rect 20416 -2910 20534 -2898
rect 20650 -2501 20768 -2489
rect 20650 -2898 20656 -2501
rect 20762 -2898 20768 -2501
rect 20650 -2910 20768 -2898
rect 20884 -2501 21002 -2489
rect 20884 -2898 20890 -2501
rect 20996 -2898 21002 -2501
rect 20884 -2910 21002 -2898
rect 21118 -2501 21236 -2489
rect 21118 -2898 21124 -2501
rect 21230 -2898 21236 -2501
rect 21118 -2910 21236 -2898
rect 21352 -2501 21470 -2489
rect 21352 -2898 21358 -2501
rect 21464 -2898 21470 -2501
rect 21352 -2910 21470 -2898
rect 21586 -2501 21704 -2489
rect 21586 -2898 21592 -2501
rect 21698 -2898 21704 -2501
rect 21586 -2910 21704 -2898
rect 21820 -2501 21938 -2489
rect 21820 -2898 21826 -2501
rect 21932 -2898 21938 -2501
rect 21820 -2910 21938 -2898
rect 22054 -2501 22172 -2489
rect 22054 -2898 22060 -2501
rect 22166 -2898 22172 -2501
rect 22054 -2910 22172 -2898
rect 22288 -2501 22406 -2489
rect 22288 -2898 22294 -2501
rect 22400 -2898 22406 -2501
rect 22288 -2910 22406 -2898
rect 22522 -2501 22640 -2489
rect 22522 -2898 22528 -2501
rect 22634 -2898 22640 -2501
rect 22522 -2910 22640 -2898
rect 22756 -2501 22874 -2489
rect 22756 -2898 22762 -2501
rect 22868 -2898 22874 -2501
rect 22756 -2910 22874 -2898
rect 22990 -2501 23108 -2489
rect 22990 -2898 22996 -2501
rect 23102 -2898 23108 -2501
rect 22990 -2910 23108 -2898
rect 23224 -2501 23342 -2489
rect 23224 -2898 23230 -2501
rect 23336 -2898 23342 -2501
rect 23224 -2910 23342 -2898
rect 23458 -2501 23576 -2489
rect 23458 -2898 23464 -2501
rect 23570 -2898 23576 -2501
rect 23458 -2910 23576 -2898
rect 23692 -2501 23810 -2489
rect 23692 -2898 23698 -2501
rect 23804 -2898 23810 -2501
rect 23692 -2910 23810 -2898
rect 23926 -2501 24044 -2489
rect 23926 -2898 23932 -2501
rect 24038 -2898 24044 -2501
rect 23926 -2910 24044 -2898
rect 24160 -2501 24278 -2489
rect 24160 -2898 24166 -2501
rect 24272 -2898 24278 -2501
rect 24160 -2910 24278 -2898
rect 24394 -2501 24512 -2489
rect 24394 -2898 24400 -2501
rect 24506 -2898 24512 -2501
rect 24394 -2910 24512 -2898
rect 24628 -2501 24746 -2489
rect 24628 -2898 24634 -2501
rect 24740 -2898 24746 -2501
rect 24628 -2910 24746 -2898
rect 24862 -2501 24980 -2489
rect 24862 -2898 24868 -2501
rect 24974 -2898 24980 -2501
rect 24862 -2910 24980 -2898
rect 25096 -2501 25214 -2489
rect 25096 -2898 25102 -2501
rect 25208 -2898 25214 -2501
rect 25096 -2910 25214 -2898
rect 25330 -2501 25448 -2489
rect 25330 -2898 25336 -2501
rect 25442 -2898 25448 -2501
rect 25330 -2910 25448 -2898
rect 25564 -2501 25682 -2489
rect 25564 -2898 25570 -2501
rect 25676 -2898 25682 -2501
rect 25564 -2910 25682 -2898
rect 25798 -2501 25916 -2489
rect 25798 -2898 25804 -2501
rect 25910 -2898 25916 -2501
rect 25798 -2910 25916 -2898
rect 26032 -2501 26150 -2489
rect 26032 -2898 26038 -2501
rect 26144 -2898 26150 -2501
rect 26032 -2910 26150 -2898
rect 26266 -2501 26384 -2489
rect 26266 -2898 26272 -2501
rect 26378 -2898 26384 -2501
rect 26266 -2910 26384 -2898
rect 26500 -2501 26618 -2489
rect 26500 -2898 26506 -2501
rect 26612 -2898 26618 -2501
rect 26500 -2910 26618 -2898
rect 26734 -2501 26852 -2489
rect 26734 -2898 26740 -2501
rect 26846 -2898 26852 -2501
rect 26734 -2910 26852 -2898
rect 26968 -2501 27086 -2489
rect 26968 -2898 26974 -2501
rect 27080 -2898 27086 -2501
rect 26968 -2910 27086 -2898
rect 27202 -2501 27320 -2489
rect 27202 -2898 27208 -2501
rect 27314 -2898 27320 -2501
rect 27202 -2910 27320 -2898
rect 27436 -2501 27554 -2489
rect 27436 -2898 27442 -2501
rect 27548 -2898 27554 -2501
rect 27436 -2910 27554 -2898
rect 27670 -2501 27788 -2489
rect 27670 -2898 27676 -2501
rect 27782 -2898 27788 -2501
rect 27670 -2910 27788 -2898
rect 27904 -2501 28022 -2489
rect 27904 -2898 27910 -2501
rect 28016 -2898 28022 -2501
rect 27904 -2910 28022 -2898
rect 28138 -2501 28256 -2489
rect 28138 -2898 28144 -2501
rect 28250 -2898 28256 -2501
rect 28138 -2910 28256 -2898
rect 28372 -2501 28490 -2489
rect 28372 -2898 28378 -2501
rect 28484 -2898 28490 -2501
rect 28372 -2910 28490 -2898
rect 28606 -2501 28724 -2489
rect 28606 -2898 28612 -2501
rect 28718 -2898 28724 -2501
rect 28606 -2910 28724 -2898
rect 28840 -2501 28958 -2489
rect 28840 -2898 28846 -2501
rect 28952 -2898 28958 -2501
rect 28840 -2910 28958 -2898
rect 29074 -2501 29192 -2489
rect 29074 -2898 29080 -2501
rect 29186 -2898 29192 -2501
rect 29074 -2910 29192 -2898
rect 29308 -2501 29426 -2489
rect 29308 -2898 29314 -2501
rect 29420 -2898 29426 -2501
rect 29308 -2910 29426 -2898
rect 29542 -2501 29660 -2489
rect 29542 -2898 29548 -2501
rect 29654 -2898 29660 -2501
rect 29542 -2910 29660 -2898
rect 29776 -2501 29894 -2489
rect 29776 -2898 29782 -2501
rect 29888 -2898 29894 -2501
rect 29776 -2910 29894 -2898
<< properties >>
string FIXED_BBOX -30017 -3029 30017 3029
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 25.0 m 1 nx 256 wmin 0.690 lmin 0.50 class resistor rho 319.8 val 12.151k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
