magic
tech sky130A
magscale 1 2
timestamp 1729620069
<< pwell >>
rect -1054 -3082 1054 3082
<< psubdiff >>
rect -1018 3012 -922 3046
rect 922 3012 1018 3046
rect -1018 2950 -984 3012
rect 984 2950 1018 3012
rect -1018 -3012 -984 -2950
rect 984 -3012 1018 -2950
rect -1018 -3046 -922 -3012
rect 922 -3046 1018 -3012
<< psubdiffcont >>
rect -922 3012 922 3046
rect -1018 -2950 -984 2950
rect 984 -2950 1018 2950
rect -922 -3046 922 -3012
<< xpolycontact >>
rect -888 2484 -750 2916
rect -888 -2916 -750 -2484
rect -654 2484 -516 2916
rect -654 -2916 -516 -2484
rect -420 2484 -282 2916
rect -420 -2916 -282 -2484
rect -186 2484 -48 2916
rect -186 -2916 -48 -2484
rect 48 2484 186 2916
rect 48 -2916 186 -2484
rect 282 2484 420 2916
rect 282 -2916 420 -2484
rect 516 2484 654 2916
rect 516 -2916 654 -2484
rect 750 2484 888 2916
rect 750 -2916 888 -2484
<< ppolyres >>
rect -888 -2484 -750 2484
rect -654 -2484 -516 2484
rect -420 -2484 -282 2484
rect -186 -2484 -48 2484
rect 48 -2484 186 2484
rect 282 -2484 420 2484
rect 516 -2484 654 2484
rect 750 -2484 888 2484
<< locali >>
rect -1018 3012 -922 3046
rect 922 3012 1018 3046
rect -1018 2950 -984 3012
rect 984 2950 1018 3012
rect -1018 -3012 -984 -2950
rect 984 -3012 1018 -2950
rect -1018 -3046 -922 -3012
rect 922 -3046 1018 -3012
<< viali >>
rect -872 2501 -766 2898
rect -638 2501 -532 2898
rect -404 2501 -298 2898
rect -170 2501 -64 2898
rect 64 2501 170 2898
rect 298 2501 404 2898
rect 532 2501 638 2898
rect 766 2501 872 2898
rect -872 -2898 -766 -2501
rect -638 -2898 -532 -2501
rect -404 -2898 -298 -2501
rect -170 -2898 -64 -2501
rect 64 -2898 170 -2501
rect 298 -2898 404 -2501
rect 532 -2898 638 -2501
rect 766 -2898 872 -2501
<< metal1 >>
rect -878 2898 -760 2910
rect -878 2501 -872 2898
rect -766 2501 -760 2898
rect -878 2489 -760 2501
rect -644 2898 -526 2910
rect -644 2501 -638 2898
rect -532 2501 -526 2898
rect -644 2489 -526 2501
rect -410 2898 -292 2910
rect -410 2501 -404 2898
rect -298 2501 -292 2898
rect -410 2489 -292 2501
rect -176 2898 -58 2910
rect -176 2501 -170 2898
rect -64 2501 -58 2898
rect -176 2489 -58 2501
rect 58 2898 176 2910
rect 58 2501 64 2898
rect 170 2501 176 2898
rect 58 2489 176 2501
rect 292 2898 410 2910
rect 292 2501 298 2898
rect 404 2501 410 2898
rect 292 2489 410 2501
rect 526 2898 644 2910
rect 526 2501 532 2898
rect 638 2501 644 2898
rect 526 2489 644 2501
rect 760 2898 878 2910
rect 760 2501 766 2898
rect 872 2501 878 2898
rect 760 2489 878 2501
rect -878 -2501 -760 -2489
rect -878 -2898 -872 -2501
rect -766 -2898 -760 -2501
rect -878 -2910 -760 -2898
rect -644 -2501 -526 -2489
rect -644 -2898 -638 -2501
rect -532 -2898 -526 -2501
rect -644 -2910 -526 -2898
rect -410 -2501 -292 -2489
rect -410 -2898 -404 -2501
rect -298 -2898 -292 -2501
rect -410 -2910 -292 -2898
rect -176 -2501 -58 -2489
rect -176 -2898 -170 -2501
rect -64 -2898 -58 -2501
rect -176 -2910 -58 -2898
rect 58 -2501 176 -2489
rect 58 -2898 64 -2501
rect 170 -2898 176 -2501
rect 58 -2910 176 -2898
rect 292 -2501 410 -2489
rect 292 -2898 298 -2501
rect 404 -2898 410 -2501
rect 292 -2910 410 -2898
rect 526 -2501 644 -2489
rect 526 -2898 532 -2501
rect 638 -2898 644 -2501
rect 526 -2910 644 -2898
rect 760 -2501 878 -2489
rect 760 -2898 766 -2501
rect 872 -2898 878 -2501
rect 760 -2910 878 -2898
<< properties >>
string FIXED_BBOX -1001 -3029 1001 3029
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 25.0 m 1 nx 8 wmin 0.690 lmin 0.50 class resistor rho 319.8 val 12.151k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
